magic
tech sky130A
magscale 1 2
timestamp 1636029542
<< metal1 >>
rect 242802 703128 242808 703180
rect 242860 703168 242866 703180
rect 348786 703168 348792 703180
rect 242860 703140 348792 703168
rect 242860 703128 242866 703140
rect 348786 703128 348792 703140
rect 348844 703128 348850 703180
rect 274542 703060 274548 703112
rect 274600 703100 274606 703112
rect 413646 703100 413652 703112
rect 274600 703072 413652 703100
rect 274600 703060 274606 703072
rect 413646 703060 413652 703072
rect 413704 703060 413710 703112
rect 184290 702992 184296 703044
rect 184348 703032 184354 703044
rect 332502 703032 332508 703044
rect 184348 703004 332508 703032
rect 184348 702992 184354 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 201494 702924 201500 702976
rect 201552 702964 201558 702976
rect 202782 702964 202788 702976
rect 201552 702936 202788 702964
rect 201552 702924 201558 702936
rect 202782 702924 202788 702936
rect 202840 702924 202846 702976
rect 280798 702924 280804 702976
rect 280856 702964 280862 702976
rect 429838 702964 429844 702976
rect 280856 702936 429844 702964
rect 280856 702924 280862 702936
rect 429838 702924 429844 702936
rect 429896 702924 429902 702976
rect 188890 702856 188896 702908
rect 188948 702896 188954 702908
rect 364978 702896 364984 702908
rect 188948 702868 364984 702896
rect 188948 702856 188954 702868
rect 364978 702856 364984 702868
rect 365036 702856 365042 702908
rect 218974 702788 218980 702840
rect 219032 702828 219038 702840
rect 269298 702828 269304 702840
rect 219032 702800 269304 702828
rect 219032 702788 219038 702800
rect 269298 702788 269304 702800
rect 269356 702788 269362 702840
rect 285582 702788 285588 702840
rect 285640 702828 285646 702840
rect 462314 702828 462320 702840
rect 285640 702800 462320 702828
rect 285640 702788 285646 702800
rect 462314 702788 462320 702800
rect 462372 702788 462378 702840
rect 169754 702720 169760 702772
rect 169812 702760 169818 702772
rect 170306 702760 170312 702772
rect 169812 702732 170312 702760
rect 169812 702720 169818 702732
rect 170306 702720 170312 702732
rect 170364 702760 170370 702772
rect 224218 702760 224224 702772
rect 170364 702732 224224 702760
rect 170364 702720 170370 702732
rect 224218 702720 224224 702732
rect 224276 702720 224282 702772
rect 248414 702720 248420 702772
rect 248472 702760 248478 702772
rect 494790 702760 494796 702772
rect 248472 702732 494796 702760
rect 248472 702720 248478 702732
rect 494790 702720 494796 702732
rect 494848 702720 494854 702772
rect 206278 702652 206284 702704
rect 206336 702692 206342 702704
rect 397362 702692 397368 702704
rect 206336 702664 397368 702692
rect 206336 702652 206342 702664
rect 397362 702652 397368 702664
rect 397420 702652 397426 702704
rect 24302 702584 24308 702636
rect 24360 702624 24366 702636
rect 85574 702624 85580 702636
rect 24360 702596 85580 702624
rect 24360 702584 24366 702596
rect 85574 702584 85580 702596
rect 85632 702584 85638 702636
rect 137830 702584 137836 702636
rect 137888 702624 137894 702636
rect 215294 702624 215300 702636
rect 137888 702596 215300 702624
rect 137888 702584 137894 702596
rect 215294 702584 215300 702596
rect 215352 702584 215358 702636
rect 222838 702584 222844 702636
rect 222896 702624 222902 702636
rect 478506 702624 478512 702636
rect 222896 702596 478512 702624
rect 222896 702584 222902 702596
rect 478506 702584 478512 702596
rect 478564 702584 478570 702636
rect 8110 702516 8116 702568
rect 8168 702556 8174 702568
rect 96614 702556 96620 702568
rect 8168 702528 96620 702556
rect 8168 702516 8174 702528
rect 96614 702516 96620 702528
rect 96672 702516 96678 702568
rect 154114 702516 154120 702568
rect 154172 702556 154178 702568
rect 233234 702556 233240 702568
rect 154172 702528 233240 702556
rect 154172 702516 154178 702528
rect 233234 702516 233240 702528
rect 233292 702516 233298 702568
rect 271138 702516 271144 702568
rect 271196 702556 271202 702568
rect 527174 702556 527180 702568
rect 271196 702528 527180 702556
rect 271196 702516 271202 702528
rect 527174 702516 527180 702528
rect 527232 702516 527238 702568
rect 67634 702448 67640 702500
rect 67692 702488 67698 702500
rect 169754 702488 169760 702500
rect 67692 702460 169760 702488
rect 67692 702448 67698 702460
rect 169754 702448 169760 702460
rect 169812 702448 169818 702500
rect 180058 702448 180064 702500
rect 180116 702488 180122 702500
rect 235166 702488 235172 702500
rect 180116 702460 235172 702488
rect 180116 702448 180122 702460
rect 235166 702448 235172 702460
rect 235224 702448 235230 702500
rect 255958 702448 255964 702500
rect 256016 702488 256022 702500
rect 543458 702488 543464 702500
rect 256016 702460 543464 702488
rect 256016 702448 256022 702460
rect 543458 702448 543464 702460
rect 543516 702448 543522 702500
rect 62022 700340 62028 700392
rect 62080 700380 62086 700392
rect 72970 700380 72976 700392
rect 62080 700352 72976 700380
rect 62080 700340 62086 700352
rect 72970 700340 72976 700352
rect 73028 700340 73034 700392
rect 84102 700340 84108 700392
rect 84160 700380 84166 700392
rect 89162 700380 89168 700392
rect 84160 700352 89168 700380
rect 84160 700340 84166 700352
rect 89162 700340 89168 700352
rect 89220 700340 89226 700392
rect 71682 700272 71688 700324
rect 71740 700312 71746 700324
rect 105446 700312 105452 700324
rect 71740 700284 105452 700312
rect 71740 700272 71746 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 251818 700272 251824 700324
rect 251876 700312 251882 700324
rect 283834 700312 283840 700324
rect 251876 700284 283840 700312
rect 251876 700272 251882 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 559650 700272 559656 700324
rect 559708 700312 559714 700324
rect 582834 700312 582840 700324
rect 559708 700284 582840 700312
rect 559708 700272 559714 700284
rect 582834 700272 582840 700284
rect 582892 700272 582898 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 33778 683176 33784 683188
rect 3476 683148 33784 683176
rect 3476 683136 3482 683148
rect 33778 683136 33784 683148
rect 33836 683136 33842 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 15838 670732 15844 670744
rect 3568 670704 15844 670732
rect 3568 670692 3574 670704
rect 15838 670692 15844 670704
rect 15896 670692 15902 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 36538 656928 36544 656940
rect 3476 656900 36544 656928
rect 3476 656888 3482 656900
rect 36538 656888 36544 656900
rect 36596 656888 36602 656940
rect 144822 622412 144828 622464
rect 144880 622452 144886 622464
rect 241514 622452 241520 622464
rect 144880 622424 241520 622452
rect 144880 622412 144886 622424
rect 241514 622412 241520 622424
rect 241572 622412 241578 622464
rect 151722 619624 151728 619676
rect 151780 619664 151786 619676
rect 251174 619664 251180 619676
rect 151780 619636 251180 619664
rect 151780 619624 151786 619636
rect 251174 619624 251180 619636
rect 251232 619664 251238 619676
rect 251818 619664 251824 619676
rect 251232 619636 251824 619664
rect 251232 619624 251238 619636
rect 251818 619624 251824 619636
rect 251876 619624 251882 619676
rect 205634 619556 205640 619608
rect 205692 619596 205698 619608
rect 206278 619596 206284 619608
rect 205692 619568 206284 619596
rect 205692 619556 205698 619568
rect 206278 619556 206284 619568
rect 206336 619556 206342 619608
rect 3510 618604 3516 618656
rect 3568 618644 3574 618656
rect 7558 618644 7564 618656
rect 3568 618616 7564 618644
rect 3568 618604 3574 618616
rect 7558 618604 7564 618616
rect 7616 618604 7622 618656
rect 178770 618332 178776 618384
rect 178828 618372 178834 618384
rect 235994 618372 236000 618384
rect 178828 618344 236000 618372
rect 178828 618332 178834 618344
rect 235994 618332 236000 618344
rect 236052 618332 236058 618384
rect 129642 618264 129648 618316
rect 129700 618304 129706 618316
rect 205634 618304 205640 618316
rect 129700 618276 205640 618304
rect 129700 618264 129706 618276
rect 205634 618264 205640 618276
rect 205692 618264 205698 618316
rect 177482 616904 177488 616956
rect 177540 616944 177546 616956
rect 242894 616944 242900 616956
rect 177540 616916 242900 616944
rect 177540 616904 177546 616916
rect 242894 616904 242900 616916
rect 242952 616904 242958 616956
rect 141970 616836 141976 616888
rect 142028 616876 142034 616888
rect 219434 616876 219440 616888
rect 142028 616848 219440 616876
rect 142028 616836 142034 616848
rect 219434 616836 219440 616848
rect 219492 616836 219498 616888
rect 233234 615952 233240 616004
rect 233292 615992 233298 616004
rect 233878 615992 233884 616004
rect 233292 615964 233884 615992
rect 233292 615952 233298 615964
rect 233878 615952 233884 615964
rect 233936 615952 233942 616004
rect 184842 615544 184848 615596
rect 184900 615584 184906 615596
rect 233234 615584 233240 615596
rect 184900 615556 233240 615584
rect 184900 615544 184906 615556
rect 233234 615544 233240 615556
rect 233292 615544 233298 615596
rect 142062 615476 142068 615528
rect 142120 615516 142126 615528
rect 213914 615516 213920 615528
rect 142120 615488 213920 615516
rect 142120 615476 142126 615488
rect 213914 615476 213920 615488
rect 213972 615476 213978 615528
rect 140682 614184 140688 614236
rect 140740 614224 140746 614236
rect 207658 614224 207664 614236
rect 140740 614196 207664 614224
rect 140740 614184 140746 614196
rect 207658 614184 207664 614196
rect 207716 614184 207722 614236
rect 152550 614116 152556 614168
rect 152608 614156 152614 614168
rect 232314 614156 232320 614168
rect 152608 614128 232320 614156
rect 152608 614116 152614 614128
rect 232314 614116 232320 614128
rect 232372 614116 232378 614168
rect 153838 612824 153844 612876
rect 153896 612864 153902 612876
rect 221642 612864 221648 612876
rect 153896 612836 221648 612864
rect 153896 612824 153902 612836
rect 221642 612824 221648 612836
rect 221700 612824 221706 612876
rect 71774 612756 71780 612808
rect 71832 612796 71838 612808
rect 258074 612796 258080 612808
rect 71832 612768 258080 612796
rect 71832 612756 71838 612768
rect 258074 612756 258080 612768
rect 258132 612756 258138 612808
rect 188982 611396 188988 611448
rect 189040 611436 189046 611448
rect 230474 611436 230480 611448
rect 189040 611408 230480 611436
rect 189040 611396 189046 611408
rect 230474 611396 230480 611408
rect 230532 611396 230538 611448
rect 67542 611328 67548 611380
rect 67600 611368 67606 611380
rect 254026 611368 254032 611380
rect 67600 611340 254032 611368
rect 67600 611328 67606 611340
rect 254026 611328 254032 611340
rect 254084 611328 254090 611380
rect 187510 610036 187516 610088
rect 187568 610076 187574 610088
rect 217226 610076 217232 610088
rect 187568 610048 217232 610076
rect 187568 610036 187574 610048
rect 217226 610036 217232 610048
rect 217284 610036 217290 610088
rect 123478 609968 123484 610020
rect 123536 610008 123542 610020
rect 256694 610008 256700 610020
rect 123536 609980 256700 610008
rect 123536 609968 123542 609980
rect 256694 609968 256700 609980
rect 256752 609968 256758 610020
rect 201494 609220 201500 609272
rect 201552 609260 201558 609272
rect 222286 609260 222292 609272
rect 201552 609232 222292 609260
rect 201552 609220 201558 609232
rect 222286 609220 222292 609232
rect 222344 609220 222350 609272
rect 182082 608676 182088 608728
rect 182140 608716 182146 608728
rect 226334 608716 226340 608728
rect 182140 608688 226340 608716
rect 182140 608676 182146 608688
rect 226334 608676 226340 608688
rect 226392 608676 226398 608728
rect 139302 608608 139308 608660
rect 139360 608648 139366 608660
rect 200666 608648 200672 608660
rect 139360 608620 200672 608648
rect 139360 608608 139366 608620
rect 200666 608608 200672 608620
rect 200724 608608 200730 608660
rect 188338 607248 188344 607300
rect 188396 607288 188402 607300
rect 196710 607288 196716 607300
rect 188396 607260 196716 607288
rect 188396 607248 188402 607260
rect 196710 607248 196716 607260
rect 196768 607248 196774 607300
rect 177390 607180 177396 607232
rect 177448 607220 177454 607232
rect 209406 607220 209412 607232
rect 177448 607192 209412 607220
rect 177448 607180 177454 607192
rect 209406 607180 209412 607192
rect 209464 607180 209470 607232
rect 215662 606432 215668 606484
rect 215720 606472 215726 606484
rect 582374 606472 582380 606484
rect 215720 606444 582380 606472
rect 215720 606432 215726 606444
rect 582374 606432 582380 606444
rect 582432 606432 582438 606484
rect 184382 605888 184388 605940
rect 184440 605928 184446 605940
rect 215662 605928 215668 605940
rect 184440 605900 215668 605928
rect 184440 605888 184446 605900
rect 215662 605888 215668 605900
rect 215720 605888 215726 605940
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 94682 605860 94688 605872
rect 3568 605832 94688 605860
rect 3568 605820 3574 605832
rect 94682 605820 94688 605832
rect 94740 605820 94746 605872
rect 98638 605820 98644 605872
rect 98696 605860 98702 605872
rect 144730 605860 144736 605872
rect 98696 605832 144736 605860
rect 98696 605820 98702 605832
rect 144730 605820 144736 605832
rect 144788 605820 144794 605872
rect 180702 605820 180708 605872
rect 180760 605860 180766 605872
rect 214374 605860 214380 605872
rect 180760 605832 214380 605860
rect 180760 605820 180766 605832
rect 214374 605820 214380 605832
rect 214432 605820 214438 605872
rect 183462 604528 183468 604580
rect 183520 604568 183526 604580
rect 206094 604568 206100 604580
rect 183520 604540 206100 604568
rect 183520 604528 183526 604540
rect 206094 604528 206100 604540
rect 206152 604528 206158 604580
rect 169018 604460 169024 604512
rect 169076 604500 169082 604512
rect 216950 604500 216956 604512
rect 169076 604472 216956 604500
rect 169076 604460 169082 604472
rect 216950 604460 216956 604472
rect 217008 604460 217014 604512
rect 241790 604460 241796 604512
rect 241848 604500 241854 604512
rect 242802 604500 242808 604512
rect 241848 604472 242808 604500
rect 241848 604460 241854 604472
rect 242802 604460 242808 604472
rect 242860 604500 242866 604512
rect 274818 604500 274824 604512
rect 242860 604472 274824 604500
rect 242860 604460 242866 604472
rect 274818 604460 274824 604472
rect 274876 604460 274882 604512
rect 289722 604460 289728 604512
rect 289780 604500 289786 604512
rect 582834 604500 582840 604512
rect 289780 604472 582840 604500
rect 289780 604460 289786 604472
rect 582834 604460 582840 604472
rect 582892 604460 582898 604512
rect 246206 603168 246212 603220
rect 246264 603208 246270 603220
rect 254578 603208 254584 603220
rect 246264 603180 254584 603208
rect 246264 603168 246270 603180
rect 254578 603168 254584 603180
rect 254636 603168 254642 603220
rect 177298 603100 177304 603152
rect 177356 603140 177362 603152
rect 203702 603140 203708 603152
rect 177356 603112 203708 603140
rect 177356 603100 177362 603112
rect 203702 603100 203708 603112
rect 203760 603100 203766 603152
rect 241054 603100 241060 603152
rect 241112 603140 241118 603152
rect 281534 603140 281540 603152
rect 241112 603112 281540 603140
rect 241112 603100 241118 603112
rect 281534 603100 281540 603112
rect 281592 603100 281598 603152
rect 222194 602148 222200 602200
rect 222252 602188 222258 602200
rect 223022 602188 223028 602200
rect 222252 602160 223028 602188
rect 222252 602148 222258 602160
rect 223022 602148 223028 602160
rect 223080 602148 223086 602200
rect 191742 601740 191748 601792
rect 191800 601780 191806 601792
rect 263686 601780 263692 601792
rect 191800 601752 263692 601780
rect 191800 601740 191806 601752
rect 263686 601740 263692 601752
rect 263744 601740 263750 601792
rect 104158 601672 104164 601724
rect 104216 601712 104222 601724
rect 211246 601712 211252 601724
rect 104216 601684 211252 601712
rect 104216 601672 104222 601684
rect 211246 601672 211252 601684
rect 211304 601672 211310 601724
rect 252462 601672 252468 601724
rect 252520 601712 252526 601724
rect 259454 601712 259460 601724
rect 252520 601684 259460 601712
rect 252520 601672 252526 601684
rect 259454 601672 259460 601684
rect 259512 601672 259518 601724
rect 224218 601604 224224 601656
rect 224276 601644 224282 601656
rect 225230 601644 225236 601656
rect 224276 601616 225236 601644
rect 224276 601604 224282 601616
rect 225230 601604 225236 601616
rect 225288 601604 225294 601656
rect 233878 601536 233884 601588
rect 233936 601576 233942 601588
rect 235350 601576 235356 601588
rect 233936 601548 235356 601576
rect 233936 601536 233942 601548
rect 235350 601536 235356 601548
rect 235408 601536 235414 601588
rect 192570 600380 192576 600432
rect 192628 600420 192634 600432
rect 204254 600420 204260 600432
rect 192628 600392 204260 600420
rect 192628 600380 192634 600392
rect 204254 600380 204260 600392
rect 204312 600380 204318 600432
rect 239766 600380 239772 600432
rect 239824 600420 239830 600432
rect 271874 600420 271880 600432
rect 239824 600392 271880 600420
rect 239824 600380 239830 600392
rect 271874 600380 271880 600392
rect 271932 600380 271938 600432
rect 148962 600312 148968 600364
rect 149020 600352 149026 600364
rect 200390 600352 200396 600364
rect 149020 600324 200396 600352
rect 149020 600312 149026 600324
rect 200390 600312 200396 600324
rect 200448 600312 200454 600364
rect 216674 600312 216680 600364
rect 216732 600352 216738 600364
rect 227806 600352 227812 600364
rect 216732 600324 227812 600352
rect 216732 600312 216738 600324
rect 227806 600312 227812 600324
rect 227864 600312 227870 600364
rect 251174 600312 251180 600364
rect 251232 600352 251238 600364
rect 299474 600352 299480 600364
rect 251232 600324 299480 600352
rect 251232 600312 251238 600324
rect 299474 600312 299480 600324
rect 299532 600312 299538 600364
rect 180766 599236 200114 599264
rect 180150 599020 180156 599072
rect 180208 599060 180214 599072
rect 180766 599060 180794 599236
rect 192478 599156 192484 599208
rect 192536 599196 192542 599208
rect 197630 599196 197636 599208
rect 192536 599168 197636 599196
rect 192536 599156 192542 599168
rect 197630 599156 197636 599168
rect 197688 599156 197694 599208
rect 193398 599088 193404 599140
rect 193456 599128 193462 599140
rect 193456 599100 195836 599128
rect 193456 599088 193462 599100
rect 180208 599032 180794 599060
rect 180208 599020 180214 599032
rect 66070 598952 66076 599004
rect 66128 598992 66134 599004
rect 187602 598992 187608 599004
rect 66128 598964 187608 598992
rect 66128 598952 66134 598964
rect 187602 598952 187608 598964
rect 187660 598952 187666 599004
rect 192662 598952 192668 599004
rect 192720 598992 192726 599004
rect 195606 598992 195612 599004
rect 192720 598964 195612 598992
rect 192720 598952 192726 598964
rect 195606 598952 195612 598964
rect 195664 598952 195670 599004
rect 195808 598992 195836 599100
rect 200086 599060 200114 599236
rect 229002 599060 229008 599072
rect 200086 599032 229008 599060
rect 229002 599020 229008 599032
rect 229060 599020 229066 599072
rect 247678 599020 247684 599072
rect 247736 599060 247742 599072
rect 257338 599060 257344 599072
rect 247736 599032 257344 599060
rect 247736 599020 247742 599032
rect 257338 599020 257344 599032
rect 257396 599020 257402 599072
rect 205174 598992 205180 599004
rect 195808 598964 205180 598992
rect 205174 598952 205180 598964
rect 205232 598952 205238 599004
rect 222930 598952 222936 599004
rect 222988 598992 222994 599004
rect 280154 598992 280160 599004
rect 222988 598964 280160 598992
rect 222988 598952 222994 598964
rect 280154 598952 280160 598964
rect 280212 598952 280218 599004
rect 192938 598884 192944 598936
rect 192996 598924 193002 598936
rect 195054 598924 195060 598936
rect 192996 598896 195060 598924
rect 192996 598884 193002 598896
rect 195054 598884 195060 598896
rect 195112 598884 195118 598936
rect 197354 598884 197360 598936
rect 197412 598884 197418 598936
rect 245194 598884 245200 598936
rect 245252 598924 245258 598936
rect 256050 598924 256056 598936
rect 245252 598896 256056 598924
rect 245252 598884 245258 598896
rect 256050 598884 256056 598896
rect 256108 598884 256114 598936
rect 193306 598816 193312 598868
rect 193364 598856 193370 598868
rect 197372 598856 197400 598884
rect 193364 598828 197400 598856
rect 193364 598816 193370 598828
rect 246758 598408 246764 598460
rect 246816 598448 246822 598460
rect 246816 598420 248414 598448
rect 246816 598408 246822 598420
rect 112438 597592 112444 597644
rect 112496 597632 112502 597644
rect 189718 597632 189724 597644
rect 112496 597604 189724 597632
rect 112496 597592 112502 597604
rect 189718 597592 189724 597604
rect 189776 597592 189782 597644
rect 161382 597524 161388 597576
rect 161440 597564 161446 597576
rect 192938 597564 192944 597576
rect 161440 597536 192944 597564
rect 161440 597524 161446 597536
rect 192938 597524 192944 597536
rect 192996 597524 193002 597576
rect 248386 597564 248414 598420
rect 255406 597592 255412 597644
rect 255464 597632 255470 597644
rect 287054 597632 287060 597644
rect 255464 597604 287060 597632
rect 255464 597592 255470 597604
rect 287054 597592 287060 597604
rect 287112 597592 287118 597644
rect 273346 597564 273352 597576
rect 248386 597536 273352 597564
rect 273346 597524 273352 597536
rect 273404 597524 273410 597576
rect 150434 596776 150440 596828
rect 150492 596816 150498 596828
rect 184382 596816 184388 596828
rect 150492 596788 184388 596816
rect 150492 596776 150498 596788
rect 184382 596776 184388 596788
rect 184440 596776 184446 596828
rect 253382 596776 253388 596828
rect 253440 596816 253446 596828
rect 293954 596816 293960 596828
rect 253440 596788 293960 596816
rect 253440 596776 253446 596788
rect 293954 596776 293960 596788
rect 294012 596776 294018 596828
rect 86954 596164 86960 596216
rect 87012 596204 87018 596216
rect 150434 596204 150440 596216
rect 87012 596176 150440 596204
rect 87012 596164 87018 596176
rect 150434 596164 150440 596176
rect 150492 596164 150498 596216
rect 255406 596164 255412 596216
rect 255464 596204 255470 596216
rect 267734 596204 267740 596216
rect 255464 596176 267740 596204
rect 255464 596164 255470 596176
rect 267734 596164 267740 596176
rect 267792 596164 267798 596216
rect 92474 595416 92480 595468
rect 92532 595456 92538 595468
rect 165522 595456 165528 595468
rect 92532 595428 165528 595456
rect 92532 595416 92538 595428
rect 165522 595416 165528 595428
rect 165580 595416 165586 595468
rect 165522 594872 165528 594924
rect 165580 594912 165586 594924
rect 166258 594912 166264 594924
rect 165580 594884 166264 594912
rect 165580 594872 165586 594884
rect 166258 594872 166264 594884
rect 166316 594872 166322 594924
rect 170398 594872 170404 594924
rect 170456 594912 170462 594924
rect 190638 594912 190644 594924
rect 170456 594884 190644 594912
rect 170456 594872 170462 594884
rect 190638 594872 190644 594884
rect 190696 594872 190702 594924
rect 159358 594804 159364 594856
rect 159416 594844 159422 594856
rect 191742 594844 191748 594856
rect 159416 594816 191748 594844
rect 159416 594804 159422 594816
rect 191742 594804 191748 594816
rect 191800 594804 191806 594856
rect 175182 594124 175188 594176
rect 175240 594164 175246 594176
rect 192754 594164 192760 594176
rect 175240 594136 192760 594164
rect 175240 594124 175246 594136
rect 192754 594124 192760 594136
rect 192812 594124 192818 594176
rect 143350 594056 143356 594108
rect 143408 594096 143414 594108
rect 192662 594096 192668 594108
rect 143408 594068 192668 594096
rect 143408 594056 143414 594068
rect 192662 594056 192668 594068
rect 192720 594056 192726 594108
rect 255314 594056 255320 594108
rect 255372 594096 255378 594108
rect 285674 594096 285680 594108
rect 255372 594068 285680 594096
rect 255372 594056 255378 594068
rect 285674 594056 285680 594068
rect 285732 594056 285738 594108
rect 69842 593376 69848 593428
rect 69900 593416 69906 593428
rect 143350 593416 143356 593428
rect 69900 593388 143356 593416
rect 69900 593376 69906 593388
rect 143350 593376 143356 593388
rect 143408 593376 143414 593428
rect 285674 593376 285680 593428
rect 285732 593416 285738 593428
rect 582650 593416 582656 593428
rect 285732 593388 582656 593416
rect 285732 593376 285738 593388
rect 582650 593376 582656 593388
rect 582708 593376 582714 593428
rect 175090 592628 175096 592680
rect 175148 592668 175154 592680
rect 192570 592668 192576 592680
rect 175148 592640 192576 592668
rect 175148 592628 175154 592640
rect 192570 592628 192576 592640
rect 192628 592628 192634 592680
rect 256326 592628 256332 592680
rect 256384 592668 256390 592680
rect 256694 592668 256700 592680
rect 256384 592640 256700 592668
rect 256384 592628 256390 592640
rect 256694 592628 256700 592640
rect 256752 592668 256758 592680
rect 284294 592668 284300 592680
rect 256752 592640 284300 592668
rect 256752 592628 256758 592640
rect 284294 592628 284300 592640
rect 284352 592668 284358 592680
rect 299566 592668 299572 592680
rect 284352 592640 299572 592668
rect 284352 592628 284358 592640
rect 299566 592628 299572 592640
rect 299624 592628 299630 592680
rect 164878 592084 164884 592136
rect 164936 592124 164942 592136
rect 191742 592124 191748 592136
rect 164936 592096 191748 592124
rect 164936 592084 164942 592096
rect 191742 592084 191748 592096
rect 191800 592084 191806 592136
rect 89714 592016 89720 592068
rect 89772 592056 89778 592068
rect 175090 592056 175096 592068
rect 89772 592028 175096 592056
rect 89772 592016 89778 592028
rect 175090 592016 175096 592028
rect 175148 592016 175154 592068
rect 95142 591268 95148 591320
rect 95200 591308 95206 591320
rect 192478 591308 192484 591320
rect 95200 591280 192484 591308
rect 95200 591268 95206 591280
rect 192478 591268 192484 591280
rect 192536 591268 192542 591320
rect 253474 591268 253480 591320
rect 253532 591308 253538 591320
rect 298094 591308 298100 591320
rect 253532 591280 298100 591308
rect 253532 591268 253538 591280
rect 298094 591268 298100 591280
rect 298152 591268 298158 591320
rect 163498 590656 163504 590708
rect 163556 590696 163562 590708
rect 191006 590696 191012 590708
rect 163556 590668 191012 590696
rect 163556 590656 163562 590668
rect 191006 590656 191012 590668
rect 191064 590656 191070 590708
rect 255406 590656 255412 590708
rect 255464 590696 255470 590708
rect 265066 590696 265072 590708
rect 255464 590668 265072 590696
rect 255464 590656 255470 590668
rect 265066 590656 265072 590668
rect 265124 590656 265130 590708
rect 77386 589976 77392 590028
rect 77444 590016 77450 590028
rect 84102 590016 84108 590028
rect 77444 589988 84108 590016
rect 77444 589976 77450 589988
rect 84102 589976 84108 589988
rect 84160 590016 84166 590028
rect 122834 590016 122840 590028
rect 84160 589988 122840 590016
rect 84160 589976 84166 589988
rect 122834 589976 122840 589988
rect 122892 589976 122898 590028
rect 36538 589908 36544 589960
rect 36596 589948 36602 589960
rect 74626 589948 74632 589960
rect 36596 589920 74632 589948
rect 36596 589908 36602 589920
rect 74626 589908 74632 589920
rect 74684 589908 74690 589960
rect 116578 589908 116584 589960
rect 116636 589948 116642 589960
rect 190546 589948 190552 589960
rect 116636 589920 190552 589948
rect 116636 589908 116642 589920
rect 190546 589908 190552 589920
rect 190604 589908 190610 589960
rect 254578 589908 254584 589960
rect 254636 589948 254642 589960
rect 292574 589948 292580 589960
rect 254636 589920 292580 589948
rect 254636 589908 254642 589920
rect 292574 589908 292580 589920
rect 292632 589908 292638 589960
rect 255406 589296 255412 589348
rect 255464 589336 255470 589348
rect 261018 589336 261024 589348
rect 255464 589308 261024 589336
rect 255464 589296 255470 589308
rect 261018 589296 261024 589308
rect 261076 589296 261082 589348
rect 40034 589228 40040 589280
rect 40092 589268 40098 589280
rect 95142 589268 95148 589280
rect 40092 589240 95148 589268
rect 40092 589228 40098 589240
rect 95142 589228 95148 589240
rect 95200 589228 95206 589280
rect 133782 588548 133788 588600
rect 133840 588588 133846 588600
rect 177390 588588 177396 588600
rect 133840 588560 177396 588588
rect 133840 588548 133846 588560
rect 177390 588548 177396 588560
rect 177448 588548 177454 588600
rect 85482 587868 85488 587920
rect 85540 587908 85546 587920
rect 133782 587908 133788 587920
rect 85540 587880 133788 587908
rect 85540 587868 85546 587880
rect 133782 587868 133788 587880
rect 133840 587868 133846 587920
rect 255406 587868 255412 587920
rect 255464 587908 255470 587920
rect 287146 587908 287152 587920
rect 255464 587880 287152 587908
rect 255464 587868 255470 587880
rect 287146 587868 287152 587880
rect 287204 587868 287210 587920
rect 81802 587120 81808 587172
rect 81860 587160 81866 587172
rect 186958 587160 186964 587172
rect 81860 587132 186964 587160
rect 81860 587120 81866 587132
rect 186958 587120 186964 587132
rect 187016 587120 187022 587172
rect 256050 587120 256056 587172
rect 256108 587160 256114 587172
rect 270494 587160 270500 587172
rect 256108 587132 270500 587160
rect 256108 587120 256114 587132
rect 270494 587120 270500 587132
rect 270552 587120 270558 587172
rect 191190 586616 191196 586628
rect 180766 586588 191196 586616
rect 150342 586508 150348 586560
rect 150400 586548 150406 586560
rect 180766 586548 180794 586588
rect 191190 586576 191196 586588
rect 191248 586576 191254 586628
rect 150400 586520 180794 586548
rect 150400 586508 150406 586520
rect 187050 586508 187056 586560
rect 187108 586548 187114 586560
rect 190454 586548 190460 586560
rect 187108 586520 190460 586548
rect 187108 586508 187114 586520
rect 190454 586508 190460 586520
rect 190512 586508 190518 586560
rect 71682 585760 71688 585812
rect 71740 585800 71746 585812
rect 106918 585800 106924 585812
rect 71740 585772 106924 585800
rect 71740 585760 71746 585772
rect 106918 585760 106924 585772
rect 106976 585760 106982 585812
rect 67358 585148 67364 585200
rect 67416 585188 67422 585200
rect 71682 585188 71688 585200
rect 67416 585160 71688 585188
rect 67416 585148 67422 585160
rect 71682 585148 71688 585160
rect 71740 585148 71746 585200
rect 92106 585148 92112 585200
rect 92164 585188 92170 585200
rect 118694 585188 118700 585200
rect 92164 585160 118700 585188
rect 92164 585148 92170 585160
rect 118694 585148 118700 585160
rect 118752 585148 118758 585200
rect 168282 585148 168288 585200
rect 168340 585188 168346 585200
rect 191742 585188 191748 585200
rect 168340 585160 191748 585188
rect 168340 585148 168346 585160
rect 191742 585148 191748 585160
rect 191800 585148 191806 585200
rect 255314 584400 255320 584452
rect 255372 584440 255378 584452
rect 258074 584440 258080 584452
rect 255372 584412 258080 584440
rect 255372 584400 255378 584412
rect 258074 584400 258080 584412
rect 258132 584440 258138 584452
rect 277486 584440 277492 584452
rect 258132 584412 277492 584440
rect 258132 584400 258138 584412
rect 277486 584400 277492 584412
rect 277544 584440 277550 584452
rect 582374 584440 582380 584452
rect 277544 584412 582380 584440
rect 277544 584400 277550 584412
rect 582374 584400 582380 584412
rect 582432 584400 582438 584452
rect 73522 583788 73528 583840
rect 73580 583828 73586 583840
rect 111058 583828 111064 583840
rect 73580 583800 111064 583828
rect 73580 583788 73586 583800
rect 111058 583788 111064 583800
rect 111116 583788 111122 583840
rect 157150 583788 157156 583840
rect 157208 583828 157214 583840
rect 191742 583828 191748 583840
rect 157208 583800 191748 583828
rect 157208 583788 157214 583800
rect 191742 583788 191748 583800
rect 191800 583788 191806 583840
rect 79042 583720 79048 583772
rect 79100 583760 79106 583772
rect 158714 583760 158720 583772
rect 79100 583732 158720 583760
rect 79100 583720 79106 583732
rect 158714 583720 158720 583732
rect 158772 583720 158778 583772
rect 255406 583652 255412 583704
rect 255464 583692 255470 583704
rect 274542 583692 274548 583704
rect 255464 583664 274548 583692
rect 255464 583652 255470 583664
rect 274542 583652 274548 583664
rect 274600 583652 274606 583704
rect 88242 583380 88248 583432
rect 88300 583420 88306 583432
rect 88978 583420 88984 583432
rect 88300 583392 88984 583420
rect 88300 583380 88306 583392
rect 88978 583380 88984 583392
rect 89036 583380 89042 583432
rect 94406 583380 94412 583432
rect 94464 583420 94470 583432
rect 98638 583420 98644 583432
rect 94464 583392 98644 583420
rect 94464 583380 94470 583392
rect 98638 583380 98644 583392
rect 98696 583380 98702 583432
rect 148686 582972 148692 583024
rect 148744 583012 148750 583024
rect 191282 583012 191288 583024
rect 148744 582984 191288 583012
rect 148744 582972 148750 582984
rect 191282 582972 191288 582984
rect 191340 582972 191346 583024
rect 274542 582972 274548 583024
rect 274600 583012 274606 583024
rect 284386 583012 284392 583024
rect 274600 582984 284392 583012
rect 274600 582972 274606 582984
rect 284386 582972 284392 582984
rect 284444 582972 284450 583024
rect 77202 582768 77208 582820
rect 77260 582808 77266 582820
rect 79318 582808 79324 582820
rect 77260 582780 79324 582808
rect 77260 582768 77266 582780
rect 79318 582768 79324 582780
rect 79376 582768 79382 582820
rect 76282 582428 76288 582480
rect 76340 582468 76346 582480
rect 95142 582468 95148 582480
rect 76340 582440 95148 582468
rect 76340 582428 76346 582440
rect 95142 582428 95148 582440
rect 95200 582428 95206 582480
rect 93762 582360 93768 582412
rect 93820 582400 93826 582412
rect 177390 582400 177396 582412
rect 93820 582372 177396 582400
rect 93820 582360 93826 582372
rect 177390 582360 177396 582372
rect 177448 582360 177454 582412
rect 182818 582360 182824 582412
rect 182876 582400 182882 582412
rect 191742 582400 191748 582412
rect 182876 582372 191748 582400
rect 182876 582360 182882 582372
rect 191742 582360 191748 582372
rect 191800 582360 191806 582412
rect 158530 581612 158536 581664
rect 158588 581652 158594 581664
rect 177482 581652 177488 581664
rect 158588 581624 177488 581652
rect 158588 581612 158594 581624
rect 177482 581612 177488 581624
rect 177540 581612 177546 581664
rect 67450 581068 67456 581120
rect 67508 581108 67514 581120
rect 124858 581108 124864 581120
rect 67508 581080 124864 581108
rect 67508 581068 67514 581080
rect 124858 581068 124864 581080
rect 124916 581068 124922 581120
rect 80238 581040 80244 581052
rect 4172 581012 80244 581040
rect 3326 580932 3332 580984
rect 3384 580972 3390 580984
rect 4172 580972 4200 581012
rect 80238 581000 80244 581012
rect 80296 581000 80302 581052
rect 176562 581000 176568 581052
rect 176620 581040 176626 581052
rect 191742 581040 191748 581052
rect 176620 581012 191748 581040
rect 176620 581000 176626 581012
rect 191742 581000 191748 581012
rect 191800 581000 191806 581052
rect 3384 580944 4200 580972
rect 3384 580932 3390 580944
rect 69014 580660 69020 580712
rect 69072 580660 69078 580712
rect 86586 580660 86592 580712
rect 86644 580660 86650 580712
rect 91002 580660 91008 580712
rect 91060 580700 91066 580712
rect 98638 580700 98644 580712
rect 91060 580672 98644 580700
rect 91060 580660 91066 580672
rect 98638 580660 98644 580672
rect 98696 580660 98702 580712
rect 63402 579708 63408 579760
rect 63460 579748 63466 579760
rect 66622 579748 66628 579760
rect 63460 579720 66628 579748
rect 63460 579708 63466 579720
rect 66622 579708 66628 579720
rect 66680 579708 66686 579760
rect 53742 579640 53748 579692
rect 53800 579680 53806 579692
rect 69032 579680 69060 580660
rect 86604 580632 86632 580660
rect 86604 580604 93854 580632
rect 93826 579748 93854 580604
rect 255958 580252 255964 580304
rect 256016 580292 256022 580304
rect 278774 580292 278780 580304
rect 256016 580264 278780 580292
rect 256016 580252 256022 580264
rect 278774 580252 278780 580264
rect 278832 580252 278838 580304
rect 161474 579748 161480 579760
rect 93826 579720 161480 579748
rect 161474 579708 161480 579720
rect 161532 579748 161538 579760
rect 188338 579748 188344 579760
rect 161532 579720 188344 579748
rect 161532 579708 161538 579720
rect 188338 579708 188344 579720
rect 188396 579708 188402 579760
rect 53800 579652 69060 579680
rect 53800 579640 53806 579652
rect 98638 579640 98644 579692
rect 98696 579680 98702 579692
rect 169754 579680 169760 579692
rect 98696 579652 169760 579680
rect 98696 579640 98702 579652
rect 169754 579640 169760 579652
rect 169812 579640 169818 579692
rect 95142 578892 95148 578944
rect 95200 578932 95206 578944
rect 108298 578932 108304 578944
rect 95200 578904 108304 578932
rect 95200 578892 95206 578904
rect 108298 578892 108304 578904
rect 108356 578892 108362 578944
rect 158714 578892 158720 578944
rect 158772 578932 158778 578944
rect 159910 578932 159916 578944
rect 158772 578904 159916 578932
rect 158772 578892 158778 578904
rect 159910 578892 159916 578904
rect 159968 578932 159974 578944
rect 184290 578932 184296 578944
rect 159968 578904 184296 578932
rect 159968 578892 159974 578904
rect 184290 578892 184296 578904
rect 184348 578892 184354 578944
rect 55122 578212 55128 578264
rect 55180 578252 55186 578264
rect 66438 578252 66444 578264
rect 55180 578224 66444 578252
rect 55180 578212 55186 578224
rect 66438 578212 66444 578224
rect 66496 578212 66502 578264
rect 96798 578212 96804 578264
rect 96856 578252 96862 578264
rect 134518 578252 134524 578264
rect 96856 578224 134524 578252
rect 96856 578212 96862 578224
rect 134518 578212 134524 578224
rect 134576 578212 134582 578264
rect 186958 578212 186964 578264
rect 187016 578252 187022 578264
rect 191558 578252 191564 578264
rect 187016 578224 191564 578252
rect 187016 578212 187022 578224
rect 191558 578212 191564 578224
rect 191616 578212 191622 578264
rect 98546 578144 98552 578196
rect 98604 578184 98610 578196
rect 191742 578184 191748 578196
rect 98604 578156 191748 578184
rect 98604 578144 98610 578156
rect 191742 578144 191748 578156
rect 191800 578144 191806 578196
rect 137922 577464 137928 577516
rect 137980 577504 137986 577516
rect 187050 577504 187056 577516
rect 137980 577476 187056 577504
rect 137980 577464 137986 577476
rect 187050 577464 187056 577476
rect 187108 577464 187114 577516
rect 255406 577464 255412 577516
rect 255464 577504 255470 577516
rect 298186 577504 298192 577516
rect 255464 577476 298192 577504
rect 255464 577464 255470 577476
rect 298186 577464 298192 577476
rect 298244 577464 298250 577516
rect 255406 576852 255412 576904
rect 255464 576892 255470 576904
rect 264974 576892 264980 576904
rect 255464 576864 264980 576892
rect 255464 576852 255470 576864
rect 264974 576852 264980 576864
rect 265032 576852 265038 576904
rect 3418 576784 3424 576836
rect 3476 576824 3482 576836
rect 67542 576824 67548 576836
rect 3476 576796 67548 576824
rect 3476 576784 3482 576796
rect 67542 576784 67548 576796
rect 67600 576784 67606 576836
rect 97902 576784 97908 576836
rect 97960 576824 97966 576836
rect 123478 576824 123484 576836
rect 97960 576796 123484 576824
rect 97960 576784 97966 576796
rect 123478 576784 123484 576796
rect 123536 576784 123542 576836
rect 94682 576036 94688 576088
rect 94740 576076 94746 576088
rect 96706 576076 96712 576088
rect 94740 576048 96712 576076
rect 94740 576036 94746 576048
rect 96706 576036 96712 576048
rect 96764 576036 96770 576088
rect 181898 575560 181904 575612
rect 181956 575600 181962 575612
rect 191006 575600 191012 575612
rect 181956 575572 191012 575600
rect 181956 575560 181962 575572
rect 191006 575560 191012 575572
rect 191064 575560 191070 575612
rect 67542 575492 67548 575544
rect 67600 575532 67606 575544
rect 67818 575532 67824 575544
rect 67600 575504 67824 575532
rect 67600 575492 67606 575504
rect 67818 575492 67824 575504
rect 67876 575492 67882 575544
rect 119430 575492 119436 575544
rect 119488 575532 119494 575544
rect 191190 575532 191196 575544
rect 119488 575504 191196 575532
rect 119488 575492 119494 575504
rect 191190 575492 191196 575504
rect 191248 575492 191254 575544
rect 255406 575492 255412 575544
rect 255464 575532 255470 575544
rect 270586 575532 270592 575544
rect 255464 575504 270592 575532
rect 255464 575492 255470 575504
rect 270586 575492 270592 575504
rect 270644 575492 270650 575544
rect 172422 574744 172428 574796
rect 172480 574784 172486 574796
rect 185578 574784 185584 574796
rect 172480 574756 185584 574784
rect 172480 574744 172486 574756
rect 185578 574744 185584 574756
rect 185636 574744 185642 574796
rect 96798 574064 96804 574116
rect 96856 574104 96862 574116
rect 151078 574104 151084 574116
rect 96856 574076 151084 574104
rect 96856 574064 96862 574076
rect 151078 574064 151084 574076
rect 151136 574064 151142 574116
rect 166350 574064 166356 574116
rect 166408 574104 166414 574116
rect 191282 574104 191288 574116
rect 166408 574076 191288 574104
rect 166408 574064 166414 574076
rect 191282 574064 191288 574076
rect 191340 574064 191346 574116
rect 255406 574064 255412 574116
rect 255464 574104 255470 574116
rect 273438 574104 273444 574116
rect 255464 574076 273444 574104
rect 255464 574064 255470 574076
rect 273438 574064 273444 574076
rect 273496 574064 273502 574116
rect 97994 573316 98000 573368
rect 98052 573356 98058 573368
rect 137094 573356 137100 573368
rect 98052 573328 137100 573356
rect 98052 573316 98058 573328
rect 137094 573316 137100 573328
rect 137152 573316 137158 573368
rect 163590 572772 163596 572824
rect 163648 572812 163654 572824
rect 191006 572812 191012 572824
rect 163648 572784 191012 572812
rect 163648 572772 163654 572784
rect 191006 572772 191012 572784
rect 191064 572772 191070 572824
rect 64598 572704 64604 572756
rect 64656 572744 64662 572756
rect 66622 572744 66628 572756
rect 64656 572716 66628 572744
rect 64656 572704 64662 572716
rect 66622 572704 66628 572716
rect 66680 572704 66686 572756
rect 96890 572704 96896 572756
rect 96948 572744 96954 572756
rect 111794 572744 111800 572756
rect 96948 572716 111800 572744
rect 96948 572704 96954 572716
rect 111794 572704 111800 572716
rect 111852 572704 111858 572756
rect 136634 572704 136640 572756
rect 136692 572744 136698 572756
rect 137094 572744 137100 572756
rect 136692 572716 137100 572744
rect 136692 572704 136698 572716
rect 137094 572704 137100 572716
rect 137152 572744 137158 572756
rect 191558 572744 191564 572756
rect 137152 572716 191564 572744
rect 137152 572704 137158 572716
rect 191558 572704 191564 572716
rect 191616 572704 191622 572756
rect 255406 572704 255412 572756
rect 255464 572744 255470 572756
rect 283558 572744 283564 572756
rect 255464 572716 283564 572744
rect 255464 572704 255470 572716
rect 283558 572704 283564 572716
rect 283616 572704 283622 572756
rect 97902 572636 97908 572688
rect 97960 572676 97966 572688
rect 112438 572676 112444 572688
rect 97960 572648 112444 572676
rect 97960 572636 97966 572648
rect 112438 572636 112444 572648
rect 112496 572636 112502 572688
rect 184290 572636 184296 572688
rect 184348 572676 184354 572688
rect 191282 572676 191288 572688
rect 184348 572648 191288 572676
rect 184348 572636 184354 572648
rect 191282 572636 191288 572648
rect 191340 572636 191346 572688
rect 111794 571956 111800 572008
rect 111852 571996 111858 572008
rect 183370 571996 183376 572008
rect 111852 571968 183376 571996
rect 111852 571956 111858 571968
rect 183370 571956 183376 571968
rect 183428 571956 183434 572008
rect 60642 571344 60648 571396
rect 60700 571384 60706 571396
rect 66622 571384 66628 571396
rect 60700 571356 66628 571384
rect 60700 571344 60706 571356
rect 66622 571344 66628 571356
rect 66680 571344 66686 571396
rect 97718 571344 97724 571396
rect 97776 571384 97782 571396
rect 101398 571384 101404 571396
rect 97776 571356 101404 571384
rect 97776 571344 97782 571356
rect 101398 571344 101404 571356
rect 101456 571344 101462 571396
rect 255406 571344 255412 571396
rect 255464 571384 255470 571396
rect 278866 571384 278872 571396
rect 255464 571356 278872 571384
rect 255464 571344 255470 571356
rect 278866 571344 278872 571356
rect 278924 571344 278930 571396
rect 188338 571276 188344 571328
rect 188396 571316 188402 571328
rect 190914 571316 190920 571328
rect 188396 571288 190920 571316
rect 188396 571276 188402 571288
rect 190914 571276 190920 571288
rect 190972 571276 190978 571328
rect 182818 570704 182824 570716
rect 161446 570676 182824 570704
rect 157242 570596 157248 570648
rect 157300 570636 157306 570648
rect 161446 570636 161474 570676
rect 182818 570664 182824 570676
rect 182876 570664 182882 570716
rect 157300 570608 161474 570636
rect 157300 570596 157306 570608
rect 182910 570596 182916 570648
rect 182968 570636 182974 570648
rect 183370 570636 183376 570648
rect 182968 570608 183376 570636
rect 182968 570596 182974 570608
rect 183370 570596 183376 570608
rect 183428 570636 183434 570648
rect 191558 570636 191564 570648
rect 183428 570608 191564 570636
rect 183428 570596 183434 570608
rect 191558 570596 191564 570608
rect 191616 570596 191622 570648
rect 255406 570596 255412 570648
rect 255464 570636 255470 570648
rect 255682 570636 255688 570648
rect 255464 570608 255688 570636
rect 255464 570596 255470 570608
rect 255682 570596 255688 570608
rect 255740 570636 255746 570648
rect 582558 570636 582564 570648
rect 255740 570608 582564 570636
rect 255740 570596 255746 570608
rect 582558 570596 582564 570608
rect 582616 570596 582622 570648
rect 57882 569916 57888 569968
rect 57940 569956 57946 569968
rect 66622 569956 66628 569968
rect 57940 569928 66628 569956
rect 57940 569916 57946 569928
rect 66622 569916 66628 569928
rect 66680 569916 66686 569968
rect 97902 569916 97908 569968
rect 97960 569956 97966 569968
rect 146938 569956 146944 569968
rect 97960 569928 146944 569956
rect 97960 569916 97966 569928
rect 146938 569916 146944 569928
rect 146996 569916 147002 569968
rect 97442 569168 97448 569220
rect 97500 569208 97506 569220
rect 178862 569208 178868 569220
rect 97500 569180 178868 569208
rect 97500 569168 97506 569180
rect 178862 569168 178868 569180
rect 178920 569168 178926 569220
rect 255406 568896 255412 568948
rect 255464 568936 255470 568948
rect 258074 568936 258080 568948
rect 255464 568908 258080 568936
rect 255464 568896 255470 568908
rect 258074 568896 258080 568908
rect 258132 568896 258138 568948
rect 255406 568556 255412 568608
rect 255464 568596 255470 568608
rect 289906 568596 289912 568608
rect 255464 568568 289912 568596
rect 255464 568556 255470 568568
rect 289906 568556 289912 568568
rect 289964 568556 289970 568608
rect 96798 568488 96804 568540
rect 96856 568528 96862 568540
rect 129642 568528 129648 568540
rect 96856 568500 129648 568528
rect 96856 568488 96862 568500
rect 129642 568488 129648 568500
rect 129700 568488 129706 568540
rect 128998 567808 129004 567860
rect 129056 567848 129062 567860
rect 186958 567848 186964 567860
rect 129056 567820 186964 567848
rect 129056 567808 129062 567820
rect 186958 567808 186964 567820
rect 187016 567808 187022 567860
rect 255498 567808 255504 567860
rect 255556 567848 255562 567860
rect 281626 567848 281632 567860
rect 255556 567820 281632 567848
rect 255556 567808 255562 567820
rect 281626 567808 281632 567820
rect 281684 567808 281690 567860
rect 255774 567264 255780 567316
rect 255832 567304 255838 567316
rect 258166 567304 258172 567316
rect 255832 567276 258172 567304
rect 255832 567264 255838 567276
rect 258166 567264 258172 567276
rect 258224 567264 258230 567316
rect 188798 567196 188804 567248
rect 188856 567236 188862 567248
rect 191742 567236 191748 567248
rect 188856 567208 191748 567236
rect 188856 567196 188862 567208
rect 191742 567196 191748 567208
rect 191800 567196 191806 567248
rect 289722 566448 289728 566500
rect 289780 566488 289786 566500
rect 582466 566488 582472 566500
rect 289780 566460 582472 566488
rect 289780 566448 289786 566460
rect 582466 566448 582472 566460
rect 582524 566448 582530 566500
rect 255682 565904 255688 565956
rect 255740 565944 255746 565956
rect 274910 565944 274916 565956
rect 255740 565916 274916 565944
rect 255740 565904 255746 565916
rect 274910 565904 274916 565916
rect 274968 565904 274974 565956
rect 52362 565836 52368 565888
rect 52420 565876 52426 565888
rect 67634 565876 67640 565888
rect 52420 565848 67640 565876
rect 52420 565836 52426 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 255590 565836 255596 565888
rect 255648 565876 255654 565888
rect 288618 565876 288624 565888
rect 255648 565848 288624 565876
rect 255648 565836 255654 565848
rect 288618 565836 288624 565848
rect 288676 565876 288682 565888
rect 289722 565876 289728 565888
rect 288676 565848 289728 565876
rect 288676 565836 288682 565848
rect 289722 565836 289728 565848
rect 289780 565836 289786 565888
rect 187694 565768 187700 565820
rect 187752 565808 187758 565820
rect 188890 565808 188896 565820
rect 187752 565780 188896 565808
rect 187752 565768 187758 565780
rect 188890 565768 188896 565780
rect 188948 565808 188954 565820
rect 190822 565808 190828 565820
rect 188948 565780 190828 565808
rect 188948 565768 188954 565780
rect 190822 565768 190828 565780
rect 190880 565768 190886 565820
rect 169202 565088 169208 565140
rect 169260 565128 169266 565140
rect 187694 565128 187700 565140
rect 169260 565100 187700 565128
rect 169260 565088 169266 565100
rect 187694 565088 187700 565100
rect 187752 565088 187758 565140
rect 39942 564408 39948 564460
rect 40000 564448 40006 564460
rect 66806 564448 66812 564460
rect 40000 564420 66812 564448
rect 40000 564408 40006 564420
rect 66806 564408 66812 564420
rect 66864 564408 66870 564460
rect 187694 564408 187700 564460
rect 187752 564448 187758 564460
rect 191098 564448 191104 564460
rect 187752 564420 191104 564448
rect 187752 564408 187758 564420
rect 191098 564408 191104 564420
rect 191156 564408 191162 564460
rect 255590 564408 255596 564460
rect 255648 564448 255654 564460
rect 269114 564448 269120 564460
rect 255648 564420 269120 564448
rect 255648 564408 255654 564420
rect 269114 564408 269120 564420
rect 269172 564408 269178 564460
rect 124858 563660 124864 563712
rect 124916 563700 124922 563712
rect 191006 563700 191012 563712
rect 124916 563672 191012 563700
rect 124916 563660 124922 563672
rect 191006 563660 191012 563672
rect 191064 563660 191070 563712
rect 64690 563048 64696 563100
rect 64748 563088 64754 563100
rect 66714 563088 66720 563100
rect 64748 563060 66720 563088
rect 64748 563048 64754 563060
rect 66714 563048 66720 563060
rect 66772 563048 66778 563100
rect 255590 563048 255596 563100
rect 255648 563088 255654 563100
rect 277394 563088 277400 563100
rect 255648 563060 277400 563088
rect 255648 563048 255654 563060
rect 277394 563048 277400 563060
rect 277452 563048 277458 563100
rect 169570 561688 169576 561740
rect 169628 561728 169634 561740
rect 191742 561728 191748 561740
rect 169628 561700 191748 561728
rect 169628 561688 169634 561700
rect 191742 561688 191748 561700
rect 191800 561688 191806 561740
rect 255590 561688 255596 561740
rect 255648 561728 255654 561740
rect 259638 561728 259644 561740
rect 255648 561700 259644 561728
rect 255648 561688 255654 561700
rect 259638 561688 259644 561700
rect 259696 561688 259702 561740
rect 259362 561008 259368 561060
rect 259420 561048 259426 561060
rect 266354 561048 266360 561060
rect 259420 561020 266360 561048
rect 259420 561008 259426 561020
rect 266354 561008 266360 561020
rect 266412 561008 266418 561060
rect 96890 560940 96896 560992
rect 96948 560980 96954 560992
rect 180150 560980 180156 560992
rect 96948 560952 180156 560980
rect 96948 560940 96954 560952
rect 180150 560940 180156 560952
rect 180208 560940 180214 560992
rect 185670 560396 185676 560448
rect 185728 560436 185734 560448
rect 191098 560436 191104 560448
rect 185728 560408 191104 560436
rect 185728 560396 185734 560408
rect 191098 560396 191104 560408
rect 191156 560396 191162 560448
rect 170950 560260 170956 560312
rect 171008 560300 171014 560312
rect 191190 560300 191196 560312
rect 171008 560272 191196 560300
rect 171008 560260 171014 560272
rect 191190 560260 191196 560272
rect 191248 560260 191254 560312
rect 255590 560260 255596 560312
rect 255648 560300 255654 560312
rect 260926 560300 260932 560312
rect 255648 560272 260932 560300
rect 255648 560260 255654 560272
rect 260926 560260 260932 560272
rect 260984 560260 260990 560312
rect 98086 559512 98092 559564
rect 98144 559552 98150 559564
rect 115198 559552 115204 559564
rect 98144 559524 115204 559552
rect 98144 559512 98150 559524
rect 115198 559512 115204 559524
rect 115256 559512 115262 559564
rect 61930 558900 61936 558952
rect 61988 558940 61994 558952
rect 66806 558940 66812 558952
rect 61988 558912 66812 558940
rect 61988 558900 61994 558912
rect 66806 558900 66812 558912
rect 66864 558900 66870 558952
rect 96982 558900 96988 558952
rect 97040 558940 97046 558952
rect 113818 558940 113824 558952
rect 97040 558912 113824 558940
rect 97040 558900 97046 558912
rect 113818 558900 113824 558912
rect 113876 558900 113882 558952
rect 255590 558900 255596 558952
rect 255648 558940 255654 558952
rect 273254 558940 273260 558952
rect 255648 558912 273260 558940
rect 255648 558900 255654 558912
rect 273254 558900 273260 558912
rect 273312 558900 273318 558952
rect 115198 558832 115204 558884
rect 115256 558872 115262 558884
rect 160738 558872 160744 558884
rect 115256 558844 160744 558872
rect 115256 558832 115262 558844
rect 160738 558832 160744 558844
rect 160796 558832 160802 558884
rect 162762 558152 162768 558204
rect 162820 558192 162826 558204
rect 187694 558192 187700 558204
rect 162820 558164 187700 558192
rect 162820 558152 162826 558164
rect 187694 558152 187700 558164
rect 187752 558152 187758 558204
rect 188338 557608 188344 557660
rect 188396 557648 188402 557660
rect 190914 557648 190920 557660
rect 188396 557620 190920 557648
rect 188396 557608 188402 557620
rect 190914 557608 190920 557620
rect 190972 557608 190978 557660
rect 181990 557540 181996 557592
rect 182048 557580 182054 557592
rect 191742 557580 191748 557592
rect 182048 557552 191748 557580
rect 182048 557540 182054 557552
rect 191742 557540 191748 557552
rect 191800 557540 191806 557592
rect 255590 557540 255596 557592
rect 255648 557580 255654 557592
rect 266354 557580 266360 557592
rect 255648 557552 266360 557580
rect 255648 557540 255654 557552
rect 266354 557540 266360 557552
rect 266412 557540 266418 557592
rect 97902 556792 97908 556844
rect 97960 556832 97966 556844
rect 115290 556832 115296 556844
rect 97960 556804 115296 556832
rect 97960 556792 97966 556804
rect 115290 556792 115296 556804
rect 115348 556792 115354 556844
rect 166442 556180 166448 556232
rect 166500 556220 166506 556232
rect 191742 556220 191748 556232
rect 166500 556192 191748 556220
rect 166500 556180 166506 556192
rect 191742 556180 191748 556192
rect 191800 556180 191806 556232
rect 255590 556180 255596 556232
rect 255648 556220 255654 556232
rect 288434 556220 288440 556232
rect 255648 556192 288440 556220
rect 255648 556180 255654 556192
rect 288434 556180 288440 556192
rect 288492 556180 288498 556232
rect 257338 555432 257344 555484
rect 257396 555472 257402 555484
rect 280246 555472 280252 555484
rect 257396 555444 280252 555472
rect 257396 555432 257402 555444
rect 280246 555432 280252 555444
rect 280304 555432 280310 555484
rect 182818 554820 182824 554872
rect 182876 554860 182882 554872
rect 188338 554860 188344 554872
rect 182876 554832 188344 554860
rect 182876 554820 182882 554832
rect 188338 554820 188344 554832
rect 188396 554820 188402 554872
rect 159450 554752 159456 554804
rect 159508 554792 159514 554804
rect 180150 554792 180156 554804
rect 159508 554764 180156 554792
rect 159508 554752 159514 554764
rect 180150 554752 180156 554764
rect 180208 554752 180214 554804
rect 184658 554752 184664 554804
rect 184716 554792 184722 554804
rect 190822 554792 190828 554804
rect 184716 554764 190828 554792
rect 184716 554752 184722 554764
rect 190822 554752 190828 554764
rect 190880 554752 190886 554804
rect 2774 553800 2780 553852
rect 2832 553840 2838 553852
rect 4798 553840 4804 553852
rect 2832 553812 4804 553840
rect 2832 553800 2838 553812
rect 4798 553800 4804 553812
rect 4856 553800 4862 553852
rect 255590 553460 255596 553512
rect 255648 553500 255654 553512
rect 260834 553500 260840 553512
rect 255648 553472 260840 553500
rect 255648 553460 255654 553472
rect 260834 553460 260840 553472
rect 260892 553460 260898 553512
rect 57790 553392 57796 553444
rect 57848 553432 57854 553444
rect 66714 553432 66720 553444
rect 57848 553404 66720 553432
rect 57848 553392 57854 553404
rect 66714 553392 66720 553404
rect 66772 553392 66778 553444
rect 171778 553392 171784 553444
rect 171836 553432 171842 553444
rect 190914 553432 190920 553444
rect 171836 553404 190920 553432
rect 171836 553392 171842 553404
rect 190914 553392 190920 553404
rect 190972 553392 190978 553444
rect 255682 553392 255688 553444
rect 255740 553432 255746 553444
rect 277578 553432 277584 553444
rect 255740 553404 277584 553432
rect 255740 553392 255746 553404
rect 277578 553392 277584 553404
rect 277636 553392 277642 553444
rect 255590 552644 255596 552696
rect 255648 552684 255654 552696
rect 259362 552684 259368 552696
rect 255648 552656 259368 552684
rect 255648 552644 255654 552656
rect 259362 552644 259368 552656
rect 259420 552684 259426 552696
rect 269206 552684 269212 552696
rect 259420 552656 269212 552684
rect 259420 552644 259426 552656
rect 269206 552644 269212 552656
rect 269264 552644 269270 552696
rect 97902 552304 97908 552356
rect 97960 552344 97966 552356
rect 100754 552344 100760 552356
rect 97960 552316 100760 552344
rect 97960 552304 97966 552316
rect 100754 552304 100760 552316
rect 100812 552304 100818 552356
rect 167638 552032 167644 552084
rect 167696 552072 167702 552084
rect 191742 552072 191748 552084
rect 167696 552044 191748 552072
rect 167696 552032 167702 552044
rect 191742 552032 191748 552044
rect 191800 552032 191806 552084
rect 105538 551284 105544 551336
rect 105596 551324 105602 551336
rect 162210 551324 162216 551336
rect 105596 551296 162216 551324
rect 105596 551284 105602 551296
rect 162210 551284 162216 551296
rect 162268 551284 162274 551336
rect 255590 550672 255596 550724
rect 255648 550712 255654 550724
rect 259546 550712 259552 550724
rect 255648 550684 259552 550712
rect 255648 550672 255654 550684
rect 259546 550672 259552 550684
rect 259604 550672 259610 550724
rect 161566 550604 161572 550656
rect 161624 550644 161630 550656
rect 162210 550644 162216 550656
rect 161624 550616 162216 550644
rect 161624 550604 161630 550616
rect 162210 550604 162216 550616
rect 162268 550644 162274 550656
rect 191374 550644 191380 550656
rect 162268 550616 191380 550644
rect 162268 550604 162274 550616
rect 191374 550604 191380 550616
rect 191432 550604 191438 550656
rect 255590 550536 255596 550588
rect 255648 550576 255654 550588
rect 269298 550576 269304 550588
rect 255648 550548 269304 550576
rect 255648 550536 255654 550548
rect 269298 550536 269304 550548
rect 269356 550576 269362 550588
rect 276106 550576 276112 550588
rect 269356 550548 276112 550576
rect 269356 550536 269362 550548
rect 276106 550536 276112 550548
rect 276164 550536 276170 550588
rect 97902 549856 97908 549908
rect 97960 549896 97966 549908
rect 160094 549896 160100 549908
rect 97960 549868 160100 549896
rect 97960 549856 97966 549868
rect 160094 549856 160100 549868
rect 160152 549856 160158 549908
rect 188338 549352 188344 549364
rect 180766 549324 188344 549352
rect 160094 549244 160100 549296
rect 160152 549284 160158 549296
rect 160738 549284 160744 549296
rect 160152 549256 160744 549284
rect 160152 549244 160158 549256
rect 160738 549244 160744 549256
rect 160796 549284 160802 549296
rect 180766 549284 180794 549324
rect 188338 549312 188344 549324
rect 188396 549312 188402 549364
rect 160796 549256 180794 549284
rect 160796 549244 160802 549256
rect 187694 549244 187700 549296
rect 187752 549284 187758 549296
rect 191742 549284 191748 549296
rect 187752 549256 191748 549284
rect 187752 549244 187758 549256
rect 191742 549244 191748 549256
rect 191800 549244 191806 549296
rect 100754 548496 100760 548548
rect 100812 548536 100818 548548
rect 112438 548536 112444 548548
rect 100812 548508 112444 548536
rect 100812 548496 100818 548508
rect 112438 548496 112444 548508
rect 112496 548496 112502 548548
rect 173618 548496 173624 548548
rect 173676 548536 173682 548548
rect 187694 548536 187700 548548
rect 173676 548508 187700 548536
rect 173676 548496 173682 548508
rect 187694 548496 187700 548508
rect 187752 548496 187758 548548
rect 187418 547884 187424 547936
rect 187476 547924 187482 547936
rect 191558 547924 191564 547936
rect 187476 547896 191564 547924
rect 187476 547884 187482 547896
rect 191558 547884 191564 547896
rect 191616 547884 191622 547936
rect 255590 547884 255596 547936
rect 255648 547924 255654 547936
rect 263594 547924 263600 547936
rect 255648 547896 263600 547924
rect 255648 547884 255654 547896
rect 263594 547884 263600 547896
rect 263652 547884 263658 547936
rect 178678 546524 178684 546576
rect 178736 546564 178742 546576
rect 191558 546564 191564 546576
rect 178736 546536 191564 546564
rect 178736 546524 178742 546536
rect 191558 546524 191564 546536
rect 191616 546524 191622 546576
rect 99374 546456 99380 546508
rect 99432 546496 99438 546508
rect 191282 546496 191288 546508
rect 99432 546468 191288 546496
rect 99432 546456 99438 546468
rect 191282 546456 191288 546468
rect 191340 546456 191346 546508
rect 255590 546456 255596 546508
rect 255648 546496 255654 546508
rect 271966 546496 271972 546508
rect 255648 546468 271972 546496
rect 255648 546456 255654 546468
rect 271966 546456 271972 546468
rect 272024 546456 272030 546508
rect 146938 545708 146944 545760
rect 146996 545748 147002 545760
rect 188430 545748 188436 545760
rect 146996 545720 188436 545748
rect 146996 545708 147002 545720
rect 188430 545708 188436 545720
rect 188488 545708 188494 545760
rect 255590 545232 255596 545284
rect 255648 545272 255654 545284
rect 258258 545272 258264 545284
rect 255648 545244 258264 545272
rect 255648 545232 255654 545244
rect 258258 545232 258264 545244
rect 258316 545232 258322 545284
rect 176470 545096 176476 545148
rect 176528 545136 176534 545148
rect 191190 545136 191196 545148
rect 176528 545108 191196 545136
rect 176528 545096 176534 545108
rect 191190 545096 191196 545108
rect 191248 545096 191254 545148
rect 180150 545028 180156 545080
rect 180208 545068 180214 545080
rect 190638 545068 190644 545080
rect 180208 545040 190644 545068
rect 180208 545028 180214 545040
rect 190638 545028 190644 545040
rect 190696 545028 190702 545080
rect 50982 543736 50988 543788
rect 51040 543776 51046 543788
rect 66806 543776 66812 543788
rect 51040 543748 66812 543776
rect 51040 543736 51046 543748
rect 66806 543736 66812 543748
rect 66864 543736 66870 543788
rect 97534 543736 97540 543788
rect 97592 543776 97598 543788
rect 104250 543776 104256 543788
rect 97592 543748 104256 543776
rect 97592 543736 97598 543748
rect 104250 543736 104256 543748
rect 104308 543736 104314 543788
rect 150250 543736 150256 543788
rect 150308 543776 150314 543788
rect 191098 543776 191104 543788
rect 150308 543748 191104 543776
rect 150308 543736 150314 543748
rect 191098 543736 191104 543748
rect 191156 543736 191162 543788
rect 255590 543736 255596 543788
rect 255648 543776 255654 543788
rect 266446 543776 266452 543788
rect 255648 543748 266452 543776
rect 255648 543736 255654 543748
rect 266446 543736 266452 543748
rect 266504 543736 266510 543788
rect 33778 542988 33784 543040
rect 33836 543028 33842 543040
rect 65978 543028 65984 543040
rect 33836 543000 65984 543028
rect 33836 542988 33842 543000
rect 65978 542988 65984 543000
rect 66036 543028 66042 543040
rect 66530 543028 66536 543040
rect 66036 543000 66536 543028
rect 66036 542988 66042 543000
rect 66530 542988 66536 543000
rect 66588 542988 66594 543040
rect 165062 542444 165068 542496
rect 165120 542484 165126 542496
rect 191558 542484 191564 542496
rect 165120 542456 191564 542484
rect 165120 542444 165126 542456
rect 191558 542444 191564 542456
rect 191616 542444 191622 542496
rect 97534 542376 97540 542428
rect 97592 542416 97598 542428
rect 146110 542416 146116 542428
rect 97592 542388 146116 542416
rect 97592 542376 97598 542388
rect 146110 542376 146116 542388
rect 146168 542416 146174 542428
rect 189074 542416 189080 542428
rect 146168 542388 189080 542416
rect 146168 542376 146174 542388
rect 189074 542376 189080 542388
rect 189132 542376 189138 542428
rect 169754 542308 169760 542360
rect 169812 542348 169818 542360
rect 179414 542348 179420 542360
rect 169812 542320 179420 542348
rect 169812 542308 169818 542320
rect 179414 542308 179420 542320
rect 179472 542348 179478 542360
rect 180058 542348 180064 542360
rect 179472 542320 180064 542348
rect 179472 542308 179478 542320
rect 180058 542308 180064 542320
rect 180116 542308 180122 542360
rect 278038 542308 278044 542360
rect 278096 542348 278102 542360
rect 285858 542348 285864 542360
rect 278096 542320 285864 542348
rect 278096 542308 278102 542320
rect 285858 542308 285864 542320
rect 285916 542308 285922 542360
rect 97902 541628 97908 541680
rect 97960 541668 97966 541680
rect 116578 541668 116584 541680
rect 97960 541640 116584 541668
rect 97960 541628 97966 541640
rect 116578 541628 116584 541640
rect 116636 541628 116642 541680
rect 155770 541628 155776 541680
rect 155828 541668 155834 541680
rect 169754 541668 169760 541680
rect 155828 541640 169760 541668
rect 155828 541628 155834 541640
rect 169754 541628 169760 541640
rect 169812 541628 169818 541680
rect 166534 540948 166540 541000
rect 166592 540988 166598 541000
rect 190822 540988 190828 541000
rect 166592 540960 190828 540988
rect 166592 540948 166598 540960
rect 190822 540948 190828 540960
rect 190880 540948 190886 541000
rect 255590 540948 255596 541000
rect 255648 540988 255654 541000
rect 262306 540988 262312 541000
rect 255648 540960 262312 540988
rect 255648 540948 255654 540960
rect 262306 540948 262312 540960
rect 262364 540948 262370 541000
rect 7558 540200 7564 540252
rect 7616 540240 7622 540252
rect 7616 540212 64874 540240
rect 7616 540200 7622 540212
rect 64846 539900 64874 540212
rect 188338 540200 188344 540252
rect 188396 540240 188402 540252
rect 191558 540240 191564 540252
rect 188396 540212 191564 540240
rect 188396 540200 188402 540212
rect 191558 540200 191564 540212
rect 191616 540200 191622 540252
rect 73154 539900 73160 539912
rect 64846 539872 73160 539900
rect 73154 539860 73160 539872
rect 73212 539860 73218 539912
rect 67266 539792 67272 539844
rect 67324 539832 67330 539844
rect 71774 539832 71780 539844
rect 67324 539804 71780 539832
rect 67324 539792 67330 539804
rect 71774 539792 71780 539804
rect 71832 539792 71838 539844
rect 59078 539588 59084 539640
rect 59136 539628 59142 539640
rect 66622 539628 66628 539640
rect 59136 539600 66628 539628
rect 59136 539588 59142 539600
rect 66622 539588 66628 539600
rect 66680 539588 66686 539640
rect 91738 539588 91744 539640
rect 91796 539628 91802 539640
rect 162854 539628 162860 539640
rect 91796 539600 162860 539628
rect 91796 539588 91802 539600
rect 162854 539588 162860 539600
rect 162912 539588 162918 539640
rect 170490 539588 170496 539640
rect 170548 539628 170554 539640
rect 191466 539628 191472 539640
rect 170548 539600 191472 539628
rect 170548 539588 170554 539600
rect 191466 539588 191472 539600
rect 191524 539588 191530 539640
rect 253106 539316 253112 539368
rect 253164 539356 253170 539368
rect 255682 539356 255688 539368
rect 253164 539328 255688 539356
rect 253164 539316 253170 539328
rect 255682 539316 255688 539328
rect 255740 539316 255746 539368
rect 122098 538840 122104 538892
rect 122156 538880 122162 538892
rect 146938 538880 146944 538892
rect 122156 538852 146944 538880
rect 122156 538840 122162 538852
rect 146938 538840 146944 538852
rect 146996 538840 147002 538892
rect 43438 538296 43444 538348
rect 43496 538336 43502 538348
rect 94590 538336 94596 538348
rect 43496 538308 94596 538336
rect 43496 538296 43502 538308
rect 94590 538296 94596 538308
rect 94648 538336 94654 538348
rect 104158 538336 104164 538348
rect 94648 538308 104164 538336
rect 94648 538296 94654 538308
rect 104158 538296 104164 538308
rect 104216 538296 104222 538348
rect 189074 538296 189080 538348
rect 189132 538336 189138 538348
rect 221366 538336 221372 538348
rect 189132 538308 221372 538336
rect 189132 538296 189138 538308
rect 221366 538296 221372 538308
rect 221424 538296 221430 538348
rect 252094 538296 252100 538348
rect 252152 538336 252158 538348
rect 258166 538336 258172 538348
rect 252152 538308 258172 538336
rect 252152 538296 252158 538308
rect 258166 538296 258172 538308
rect 258224 538296 258230 538348
rect 85850 538228 85856 538280
rect 85908 538268 85914 538280
rect 96430 538268 96436 538280
rect 85908 538240 96436 538268
rect 85908 538228 85914 538240
rect 96430 538228 96436 538240
rect 96488 538268 96494 538280
rect 99374 538268 99380 538280
rect 96488 538240 99380 538268
rect 96488 538228 96494 538240
rect 99374 538228 99380 538240
rect 99432 538228 99438 538280
rect 177390 538228 177396 538280
rect 177448 538268 177454 538280
rect 238662 538268 238668 538280
rect 177448 538240 238668 538268
rect 177448 538228 177454 538240
rect 238662 538228 238668 538240
rect 238720 538228 238726 538280
rect 255590 538228 255596 538280
rect 255648 538268 255654 538280
rect 282914 538268 282920 538280
rect 255648 538240 282920 538268
rect 255648 538228 255654 538240
rect 282914 538228 282920 538240
rect 282972 538228 282978 538280
rect 4798 538160 4804 538212
rect 4856 538200 4862 538212
rect 70946 538200 70952 538212
rect 4856 538172 70952 538200
rect 4856 538160 4862 538172
rect 70946 538160 70952 538172
rect 71004 538160 71010 538212
rect 79226 538160 79232 538212
rect 79284 538200 79290 538212
rect 119430 538200 119436 538212
rect 79284 538172 119436 538200
rect 79284 538160 79290 538172
rect 119430 538160 119436 538172
rect 119488 538160 119494 538212
rect 178862 538160 178868 538212
rect 178920 538200 178926 538212
rect 244366 538200 244372 538212
rect 178920 538172 244372 538200
rect 178920 538160 178926 538172
rect 244366 538160 244372 538172
rect 244424 538160 244430 538212
rect 62022 537480 62028 537532
rect 62080 537520 62086 537532
rect 73154 537520 73160 537532
rect 62080 537492 73160 537520
rect 62080 537480 62086 537492
rect 73154 537480 73160 537492
rect 73212 537480 73218 537532
rect 144638 537480 144644 537532
rect 144696 537520 144702 537532
rect 222102 537520 222108 537532
rect 144696 537492 222108 537520
rect 144696 537480 144702 537492
rect 222102 537480 222108 537492
rect 222160 537480 222166 537532
rect 244274 537480 244280 537532
rect 244332 537520 244338 537532
rect 582374 537520 582380 537532
rect 244332 537492 582380 537520
rect 244332 537480 244338 537492
rect 582374 537480 582380 537492
rect 582432 537480 582438 537532
rect 79226 537004 79232 537056
rect 79284 537044 79290 537056
rect 79962 537044 79968 537056
rect 79284 537016 79968 537044
rect 79284 537004 79290 537016
rect 79962 537004 79968 537016
rect 80020 537004 80026 537056
rect 59170 536800 59176 536852
rect 59228 536840 59234 536852
rect 62022 536840 62028 536852
rect 59228 536812 62028 536840
rect 59228 536800 59234 536812
rect 62022 536800 62028 536812
rect 62080 536800 62086 536852
rect 88242 536800 88248 536852
rect 88300 536840 88306 536852
rect 95418 536840 95424 536852
rect 88300 536812 95424 536840
rect 88300 536800 88306 536812
rect 95418 536800 95424 536812
rect 95476 536800 95482 536852
rect 244366 536800 244372 536852
rect 244424 536840 244430 536852
rect 244826 536840 244832 536852
rect 244424 536812 244832 536840
rect 244424 536800 244430 536812
rect 244826 536800 244832 536812
rect 244884 536800 244890 536852
rect 249702 536800 249708 536852
rect 249760 536840 249766 536852
rect 254118 536840 254124 536852
rect 249760 536812 254124 536840
rect 249760 536800 249766 536812
rect 254118 536800 254124 536812
rect 254176 536800 254182 536852
rect 285582 536840 285588 536852
rect 284588 536812 285588 536840
rect 73154 536732 73160 536784
rect 73212 536772 73218 536784
rect 76742 536772 76748 536784
rect 73212 536744 76748 536772
rect 73212 536732 73218 536744
rect 76742 536732 76748 536744
rect 76800 536732 76806 536784
rect 93394 536732 93400 536784
rect 93452 536772 93458 536784
rect 246758 536772 246764 536784
rect 93452 536744 246764 536772
rect 93452 536732 93458 536744
rect 246758 536732 246764 536744
rect 246816 536772 246822 536784
rect 284588 536772 284616 536812
rect 285582 536800 285588 536812
rect 285640 536840 285646 536852
rect 291194 536840 291200 536852
rect 285640 536812 291200 536840
rect 285640 536800 285646 536812
rect 291194 536800 291200 536812
rect 291252 536800 291258 536852
rect 246816 536744 284616 536772
rect 246816 536732 246822 536744
rect 82170 536664 82176 536716
rect 82228 536704 82234 536716
rect 91738 536704 91744 536716
rect 82228 536676 91744 536704
rect 82228 536664 82234 536676
rect 91738 536664 91744 536676
rect 91796 536664 91802 536716
rect 239214 536664 239220 536716
rect 239272 536704 239278 536716
rect 244274 536704 244280 536716
rect 239272 536676 244280 536704
rect 239272 536664 239278 536676
rect 244274 536664 244280 536676
rect 244332 536664 244338 536716
rect 68922 536528 68928 536580
rect 68980 536568 68986 536580
rect 72418 536568 72424 536580
rect 68980 536540 72424 536568
rect 68980 536528 68986 536540
rect 72418 536528 72424 536540
rect 72476 536528 72482 536580
rect 195974 536188 195980 536240
rect 196032 536228 196038 536240
rect 197630 536228 197636 536240
rect 196032 536200 197636 536228
rect 196032 536188 196038 536200
rect 197630 536188 197636 536200
rect 197688 536188 197694 536240
rect 244918 536120 244924 536172
rect 244976 536160 244982 536172
rect 245930 536160 245936 536172
rect 244976 536132 245936 536160
rect 244976 536120 244982 536132
rect 245930 536120 245936 536132
rect 245988 536120 245994 536172
rect 3418 536052 3424 536104
rect 3476 536092 3482 536104
rect 41322 536092 41328 536104
rect 3476 536064 41328 536092
rect 3476 536052 3482 536064
rect 41322 536052 41328 536064
rect 41380 536092 41386 536104
rect 69382 536092 69388 536104
rect 41380 536064 69388 536092
rect 41380 536052 41386 536064
rect 69382 536052 69388 536064
rect 69440 536052 69446 536104
rect 70946 536052 70952 536104
rect 71004 536092 71010 536104
rect 86218 536092 86224 536104
rect 71004 536064 86224 536092
rect 71004 536052 71010 536064
rect 86218 536052 86224 536064
rect 86276 536052 86282 536104
rect 189810 536052 189816 536104
rect 189868 536092 189874 536104
rect 193582 536092 193588 536104
rect 189868 536064 193588 536092
rect 189868 536052 189874 536064
rect 193582 536052 193588 536064
rect 193640 536052 193646 536104
rect 225230 536052 225236 536104
rect 225288 536092 225294 536104
rect 226978 536092 226984 536104
rect 225288 536064 226984 536092
rect 225288 536052 225294 536064
rect 226978 536052 226984 536064
rect 227036 536052 227042 536104
rect 86678 535916 86684 535968
rect 86736 535956 86742 535968
rect 87598 535956 87604 535968
rect 86736 535928 87604 535956
rect 86736 535916 86742 535928
rect 87598 535916 87604 535928
rect 87656 535916 87662 535968
rect 214650 535508 214656 535560
rect 214708 535548 214714 535560
rect 216398 535548 216404 535560
rect 214708 535520 216404 535548
rect 214708 535508 214714 535520
rect 216398 535508 216404 535520
rect 216456 535508 216462 535560
rect 91002 535440 91008 535492
rect 91060 535480 91066 535492
rect 91830 535480 91836 535492
rect 91060 535452 91836 535480
rect 91060 535440 91066 535452
rect 91830 535440 91836 535452
rect 91888 535440 91894 535492
rect 215938 535440 215944 535492
rect 215996 535480 216002 535492
rect 216950 535480 216956 535492
rect 215996 535452 216956 535480
rect 215996 535440 216002 535452
rect 216950 535440 216956 535452
rect 217008 535440 217014 535492
rect 231670 535440 231676 535492
rect 231728 535480 231734 535492
rect 233878 535480 233884 535492
rect 231728 535452 233884 535480
rect 231728 535440 231734 535452
rect 233878 535440 233884 535452
rect 233936 535440 233942 535492
rect 246298 535440 246304 535492
rect 246356 535480 246362 535492
rect 247494 535480 247500 535492
rect 246356 535452 247500 535480
rect 246356 535440 246362 535452
rect 247494 535440 247500 535452
rect 247552 535440 247558 535492
rect 106918 535372 106924 535424
rect 106976 535412 106982 535424
rect 143534 535412 143540 535424
rect 106976 535384 143540 535412
rect 106976 535372 106982 535384
rect 143534 535372 143540 535384
rect 143592 535412 143598 535424
rect 144638 535412 144644 535424
rect 143592 535384 144644 535412
rect 143592 535372 143598 535384
rect 144638 535372 144644 535384
rect 144696 535372 144702 535424
rect 163866 535372 163872 535424
rect 163924 535412 163930 535424
rect 197354 535412 197360 535424
rect 163924 535384 197360 535412
rect 163924 535372 163930 535384
rect 197354 535372 197360 535384
rect 197412 535372 197418 535424
rect 206370 535236 206376 535288
rect 206428 535276 206434 535288
rect 209958 535276 209964 535288
rect 206428 535248 209964 535276
rect 206428 535236 206434 535248
rect 209958 535236 209964 535248
rect 210016 535236 210022 535288
rect 217318 534828 217324 534880
rect 217376 534868 217382 534880
rect 239766 534868 239772 534880
rect 217376 534840 239772 534868
rect 217376 534828 217382 534840
rect 239766 534828 239772 534840
rect 239824 534828 239830 534880
rect 231210 534760 231216 534812
rect 231268 534800 231274 534812
rect 254026 534800 254032 534812
rect 231268 534772 254032 534800
rect 231268 534760 231274 534772
rect 254026 534760 254032 534772
rect 254084 534760 254090 534812
rect 48130 534692 48136 534744
rect 48188 534732 48194 534744
rect 96890 534732 96896 534744
rect 48188 534704 96896 534732
rect 48188 534692 48194 534704
rect 96890 534692 96896 534704
rect 96948 534692 96954 534744
rect 178770 534692 178776 534744
rect 178828 534732 178834 534744
rect 230382 534732 230388 534744
rect 178828 534704 230388 534732
rect 178828 534692 178834 534704
rect 230382 534692 230388 534704
rect 230440 534692 230446 534744
rect 251910 534692 251916 534744
rect 251968 534732 251974 534744
rect 281718 534732 281724 534744
rect 251968 534704 281724 534732
rect 251968 534692 251974 534704
rect 281718 534692 281724 534704
rect 281776 534692 281782 534744
rect 162854 534420 162860 534472
rect 162912 534460 162918 534472
rect 163866 534460 163872 534472
rect 162912 534432 163872 534460
rect 162912 534420 162918 534432
rect 163866 534420 163872 534432
rect 163924 534420 163930 534472
rect 67358 534012 67364 534064
rect 67416 534052 67422 534064
rect 158714 534052 158720 534064
rect 67416 534024 158720 534052
rect 67416 534012 67422 534024
rect 158714 534012 158720 534024
rect 158772 534012 158778 534064
rect 180610 534012 180616 534064
rect 180668 534052 180674 534064
rect 209406 534052 209412 534064
rect 180668 534024 209412 534052
rect 180668 534012 180674 534024
rect 209406 534012 209412 534024
rect 209464 534012 209470 534064
rect 158714 533536 158720 533588
rect 158772 533576 158778 533588
rect 159450 533576 159456 533588
rect 158772 533548 159456 533576
rect 158772 533536 158778 533548
rect 159450 533536 159456 533548
rect 159508 533536 159514 533588
rect 195974 533400 195980 533452
rect 196032 533440 196038 533452
rect 196894 533440 196900 533452
rect 196032 533412 196900 533440
rect 196032 533400 196038 533412
rect 196894 533400 196900 533412
rect 196952 533400 196958 533452
rect 197354 533400 197360 533452
rect 197412 533440 197418 533452
rect 198182 533440 198188 533452
rect 197412 533412 198188 533440
rect 197412 533400 197418 533412
rect 198182 533400 198188 533412
rect 198240 533400 198246 533452
rect 200390 533440 200396 533452
rect 200086 533412 200396 533440
rect 82722 533332 82728 533384
rect 82780 533372 82786 533384
rect 94682 533372 94688 533384
rect 82780 533344 94688 533372
rect 82780 533332 82786 533344
rect 94682 533332 94688 533344
rect 94740 533332 94746 533384
rect 187694 533332 187700 533384
rect 187752 533372 187758 533384
rect 200086 533372 200114 533412
rect 200390 533400 200396 533412
rect 200448 533400 200454 533452
rect 211798 533400 211804 533452
rect 211856 533440 211862 533452
rect 212534 533440 212540 533452
rect 211856 533412 212540 533440
rect 211856 533400 211862 533412
rect 212534 533400 212540 533412
rect 212592 533400 212598 533452
rect 213178 533400 213184 533452
rect 213236 533440 213242 533452
rect 222654 533440 222660 533452
rect 213236 533412 222660 533440
rect 213236 533400 213242 533412
rect 222654 533400 222660 533412
rect 222712 533400 222718 533452
rect 227806 533400 227812 533452
rect 227864 533440 227870 533452
rect 239398 533440 239404 533452
rect 227864 533412 239404 533440
rect 227864 533400 227870 533412
rect 239398 533400 239404 533412
rect 239456 533400 239462 533452
rect 244550 533400 244556 533452
rect 244608 533440 244614 533452
rect 245010 533440 245016 533452
rect 244608 533412 245016 533440
rect 244608 533400 244614 533412
rect 245010 533400 245016 533412
rect 245068 533400 245074 533452
rect 248414 533400 248420 533452
rect 248472 533440 248478 533452
rect 248966 533440 248972 533452
rect 248472 533412 248972 533440
rect 248472 533400 248478 533412
rect 248966 533400 248972 533412
rect 249024 533400 249030 533452
rect 250438 533400 250444 533452
rect 250496 533440 250502 533452
rect 259638 533440 259644 533452
rect 250496 533412 259644 533440
rect 250496 533400 250502 533412
rect 259638 533400 259644 533412
rect 259696 533400 259702 533452
rect 187752 533344 200114 533372
rect 187752 533332 187758 533344
rect 201494 533332 201500 533384
rect 201552 533372 201558 533384
rect 202046 533372 202052 533384
rect 201552 533344 202052 533372
rect 201552 533332 201558 533344
rect 202046 533332 202052 533344
rect 202104 533332 202110 533384
rect 206278 533332 206284 533384
rect 206336 533372 206342 533384
rect 206336 533344 219434 533372
rect 206336 533332 206342 533344
rect 219406 533304 219434 533344
rect 233234 533332 233240 533384
rect 233292 533372 233298 533384
rect 233694 533372 233700 533384
rect 233292 533344 233700 533372
rect 233292 533332 233298 533344
rect 233694 533332 233700 533344
rect 233752 533332 233758 533384
rect 238662 533332 238668 533384
rect 238720 533372 238726 533384
rect 273530 533372 273536 533384
rect 238720 533344 273536 533372
rect 238720 533332 238726 533344
rect 273530 533332 273536 533344
rect 273588 533332 273594 533384
rect 236638 533304 236644 533316
rect 219406 533276 236644 533304
rect 236638 533264 236644 533276
rect 236696 533264 236702 533316
rect 209038 532924 209044 532976
rect 209096 532964 209102 532976
rect 211246 532964 211252 532976
rect 209096 532936 211252 532964
rect 209096 532924 209102 532936
rect 211246 532924 211252 532936
rect 211304 532924 211310 532976
rect 240134 532856 240140 532908
rect 240192 532896 240198 532908
rect 240686 532896 240692 532908
rect 240192 532868 240692 532896
rect 240192 532856 240198 532868
rect 240686 532856 240692 532868
rect 240744 532856 240750 532908
rect 112438 532652 112444 532704
rect 112496 532692 112502 532704
rect 113082 532692 113088 532704
rect 112496 532664 113088 532692
rect 112496 532652 112502 532664
rect 113082 532652 113088 532664
rect 113140 532692 113146 532704
rect 187694 532692 187700 532704
rect 113140 532664 187700 532692
rect 113140 532652 113146 532664
rect 187694 532652 187700 532664
rect 187752 532652 187758 532704
rect 179322 532584 179328 532636
rect 179380 532624 179386 532636
rect 206830 532624 206836 532636
rect 179380 532596 206836 532624
rect 179380 532584 179386 532596
rect 206830 532584 206836 532596
rect 206888 532584 206894 532636
rect 75822 532040 75828 532092
rect 75880 532080 75886 532092
rect 96798 532080 96804 532092
rect 75880 532052 96804 532080
rect 75880 532040 75886 532052
rect 96798 532040 96804 532052
rect 96856 532040 96862 532092
rect 73430 531972 73436 532024
rect 73488 532012 73494 532024
rect 102778 532012 102784 532024
rect 73488 531984 102784 532012
rect 73488 531972 73494 531984
rect 102778 531972 102784 531984
rect 102836 531972 102842 532024
rect 246206 531972 246212 532024
rect 246264 532012 246270 532024
rect 281810 532012 281816 532024
rect 246264 531984 281816 532012
rect 246264 531972 246270 531984
rect 281810 531972 281816 531984
rect 281868 531972 281874 532024
rect 64690 531224 64696 531276
rect 64748 531264 64754 531276
rect 223574 531264 223580 531276
rect 64748 531236 223580 531264
rect 64748 531224 64754 531236
rect 223574 531224 223580 531236
rect 223632 531224 223638 531276
rect 93118 531156 93124 531208
rect 93176 531196 93182 531208
rect 94038 531196 94044 531208
rect 93176 531168 94044 531196
rect 93176 531156 93182 531168
rect 94038 531156 94044 531168
rect 94096 531156 94102 531208
rect 190362 530544 190368 530596
rect 190420 530584 190426 530596
rect 200206 530584 200212 530596
rect 190420 530556 200212 530584
rect 190420 530544 190426 530556
rect 200206 530544 200212 530556
rect 200264 530544 200270 530596
rect 228358 530544 228364 530596
rect 228416 530584 228422 530596
rect 247586 530584 247592 530596
rect 228416 530556 247592 530584
rect 228416 530544 228422 530556
rect 247586 530544 247592 530556
rect 247644 530544 247650 530596
rect 247678 530544 247684 530596
rect 247736 530584 247742 530596
rect 256694 530584 256700 530596
rect 247736 530556 256700 530584
rect 247736 530544 247742 530556
rect 256694 530544 256700 530556
rect 256752 530544 256758 530596
rect 214558 529932 214564 529984
rect 214616 529972 214622 529984
rect 219618 529972 219624 529984
rect 214616 529944 219624 529972
rect 214616 529932 214622 529944
rect 219618 529932 219624 529944
rect 219676 529932 219682 529984
rect 191650 529864 191656 529916
rect 191708 529904 191714 529916
rect 198826 529904 198832 529916
rect 191708 529876 198832 529904
rect 191708 529864 191714 529876
rect 198826 529864 198832 529876
rect 198884 529864 198890 529916
rect 213914 529728 213920 529780
rect 213972 529768 213978 529780
rect 214742 529768 214748 529780
rect 213972 529740 214748 529768
rect 213972 529728 213978 529740
rect 214742 529728 214748 529740
rect 214800 529728 214806 529780
rect 71866 529252 71872 529304
rect 71924 529292 71930 529304
rect 122098 529292 122104 529304
rect 71924 529264 122104 529292
rect 71924 529252 71930 529264
rect 122098 529252 122104 529264
rect 122156 529252 122162 529304
rect 193122 529252 193128 529304
rect 193180 529292 193186 529304
rect 207198 529292 207204 529304
rect 193180 529264 207204 529292
rect 193180 529252 193186 529264
rect 207198 529252 207204 529264
rect 207256 529252 207262 529304
rect 67450 529184 67456 529236
rect 67508 529224 67514 529236
rect 126882 529224 126888 529236
rect 67508 529196 126888 529224
rect 67508 529184 67514 529196
rect 126882 529184 126888 529196
rect 126940 529224 126946 529236
rect 166534 529224 166540 529236
rect 126940 529196 166540 529224
rect 126940 529184 126946 529196
rect 166534 529184 166540 529196
rect 166592 529184 166598 529236
rect 204530 529184 204536 529236
rect 204588 529224 204594 529236
rect 238018 529224 238024 529236
rect 204588 529196 238024 529224
rect 204588 529184 204594 529196
rect 238018 529184 238024 529196
rect 238076 529184 238082 529236
rect 242894 529184 242900 529236
rect 242952 529224 242958 529236
rect 291286 529224 291292 529236
rect 242952 529196 291292 529224
rect 242952 529184 242958 529196
rect 291286 529184 291292 529196
rect 291344 529184 291350 529236
rect 3142 528504 3148 528556
rect 3200 528544 3206 528556
rect 97994 528544 98000 528556
rect 3200 528516 98000 528544
rect 3200 528504 3206 528516
rect 97994 528504 98000 528516
rect 98052 528504 98058 528556
rect 104250 528504 104256 528556
rect 104308 528544 104314 528556
rect 104802 528544 104808 528556
rect 104308 528516 104808 528544
rect 104308 528504 104314 528516
rect 104802 528504 104808 528516
rect 104860 528544 104866 528556
rect 197630 528544 197636 528556
rect 104860 528516 197636 528544
rect 104860 528504 104866 528516
rect 197630 528504 197636 528516
rect 197688 528504 197694 528556
rect 164970 527892 164976 527944
rect 165028 527932 165034 527944
rect 205634 527932 205640 527944
rect 165028 527904 205640 527932
rect 165028 527892 165034 527904
rect 205634 527892 205640 527904
rect 205692 527892 205698 527944
rect 244918 527892 244924 527944
rect 244976 527932 244982 527944
rect 266538 527932 266544 527944
rect 244976 527904 266544 527932
rect 244976 527892 244982 527904
rect 266538 527892 266544 527904
rect 266596 527892 266602 527944
rect 201586 527824 201592 527876
rect 201644 527864 201650 527876
rect 248598 527864 248604 527876
rect 201644 527836 248604 527864
rect 201644 527824 201650 527836
rect 248598 527824 248604 527836
rect 248656 527824 248662 527876
rect 62022 526396 62028 526448
rect 62080 526436 62086 526448
rect 96706 526436 96712 526448
rect 62080 526408 96712 526436
rect 62080 526396 62086 526408
rect 96706 526396 96712 526408
rect 96764 526396 96770 526448
rect 196066 526396 196072 526448
rect 196124 526436 196130 526448
rect 219434 526436 219440 526448
rect 196124 526408 219440 526436
rect 196124 526396 196130 526408
rect 219434 526396 219440 526408
rect 219492 526396 219498 526448
rect 226242 526260 226248 526312
rect 226300 526300 226306 526312
rect 229278 526300 229284 526312
rect 226300 526272 229284 526300
rect 226300 526260 226306 526272
rect 229278 526260 229284 526272
rect 229336 526260 229342 526312
rect 218698 525036 218704 525088
rect 218756 525076 218762 525088
rect 237466 525076 237472 525088
rect 218756 525048 237472 525076
rect 218756 525036 218762 525048
rect 237466 525036 237472 525048
rect 237524 525036 237530 525088
rect 248506 525036 248512 525088
rect 248564 525076 248570 525088
rect 265158 525076 265164 525088
rect 248564 525048 265164 525076
rect 248564 525036 248570 525048
rect 265158 525036 265164 525048
rect 265216 525036 265222 525088
rect 60642 524356 60648 524408
rect 60700 524396 60706 524408
rect 165614 524396 165620 524408
rect 60700 524368 165620 524396
rect 60700 524356 60706 524368
rect 165614 524356 165620 524368
rect 165672 524396 165678 524408
rect 166442 524396 166448 524408
rect 165672 524368 166448 524396
rect 165672 524356 165678 524368
rect 166442 524356 166448 524368
rect 166500 524356 166506 524408
rect 187326 523744 187332 523796
rect 187384 523784 187390 523796
rect 197446 523784 197452 523796
rect 187384 523756 197452 523784
rect 187384 523744 187390 523756
rect 197446 523744 197452 523756
rect 197504 523744 197510 523796
rect 196618 523676 196624 523728
rect 196676 523716 196682 523728
rect 222194 523716 222200 523728
rect 196676 523688 222200 523716
rect 196676 523676 196682 523688
rect 222194 523676 222200 523688
rect 222252 523676 222258 523728
rect 146938 522928 146944 522980
rect 146996 522968 147002 522980
rect 147398 522968 147404 522980
rect 146996 522940 147404 522968
rect 146996 522928 147002 522940
rect 147398 522928 147404 522940
rect 147456 522968 147462 522980
rect 214650 522968 214656 522980
rect 147456 522940 214656 522968
rect 147456 522928 147462 522940
rect 214650 522928 214656 522940
rect 214708 522928 214714 522980
rect 226978 522928 226984 522980
rect 227036 522968 227042 522980
rect 229094 522968 229100 522980
rect 227036 522940 229100 522968
rect 227036 522928 227042 522940
rect 229094 522928 229100 522940
rect 229152 522928 229158 522980
rect 3418 522248 3424 522300
rect 3476 522288 3482 522300
rect 93118 522288 93124 522300
rect 3476 522260 93124 522288
rect 3476 522248 3482 522260
rect 93118 522248 93124 522260
rect 93176 522288 93182 522300
rect 94498 522288 94504 522300
rect 93176 522260 94504 522288
rect 93176 522248 93182 522260
rect 94498 522248 94504 522260
rect 94556 522248 94562 522300
rect 244550 522248 244556 522300
rect 244608 522288 244614 522300
rect 270678 522288 270684 522300
rect 244608 522260 270684 522288
rect 244608 522248 244614 522260
rect 270678 522248 270684 522260
rect 270736 522248 270742 522300
rect 203518 520956 203524 521008
rect 203576 520996 203582 521008
rect 258166 520996 258172 521008
rect 203576 520968 258172 520996
rect 203576 520956 203582 520968
rect 258166 520956 258172 520968
rect 258224 520956 258230 521008
rect 141878 520888 141884 520940
rect 141936 520928 141942 520940
rect 204254 520928 204260 520940
rect 141936 520900 204260 520928
rect 141936 520888 141942 520900
rect 204254 520888 204260 520900
rect 204312 520888 204318 520940
rect 128262 519596 128268 519648
rect 128320 519636 128326 519648
rect 200114 519636 200120 519648
rect 128320 519608 200120 519636
rect 128320 519596 128326 519608
rect 200114 519596 200120 519608
rect 200172 519596 200178 519648
rect 178862 519528 178868 519580
rect 178920 519568 178926 519580
rect 261018 519568 261024 519580
rect 178920 519540 261024 519568
rect 178920 519528 178926 519540
rect 261018 519528 261024 519540
rect 261076 519528 261082 519580
rect 171042 518236 171048 518288
rect 171100 518276 171106 518288
rect 215938 518276 215944 518288
rect 171100 518248 215944 518276
rect 171100 518236 171106 518248
rect 215938 518236 215944 518248
rect 215996 518236 216002 518288
rect 72418 518168 72424 518220
rect 72476 518208 72482 518220
rect 99466 518208 99472 518220
rect 72476 518180 99472 518208
rect 72476 518168 72482 518180
rect 99466 518168 99472 518180
rect 99524 518168 99530 518220
rect 137830 518168 137836 518220
rect 137888 518208 137894 518220
rect 189810 518208 189816 518220
rect 137888 518180 189816 518208
rect 137888 518168 137894 518180
rect 189810 518168 189816 518180
rect 189868 518168 189874 518220
rect 195238 518168 195244 518220
rect 195296 518208 195302 518220
rect 206370 518208 206376 518220
rect 195296 518180 206376 518208
rect 195296 518168 195302 518180
rect 206370 518168 206376 518180
rect 206428 518168 206434 518220
rect 65794 517148 65800 517200
rect 65852 517188 65858 517200
rect 69658 517188 69664 517200
rect 65852 517160 69664 517188
rect 65852 517148 65858 517160
rect 69658 517148 69664 517160
rect 69716 517148 69722 517200
rect 204898 515448 204904 515500
rect 204956 515488 204962 515500
rect 240226 515488 240232 515500
rect 204956 515460 240232 515488
rect 204956 515448 204962 515460
rect 240226 515448 240232 515460
rect 240284 515448 240290 515500
rect 63402 515380 63408 515432
rect 63460 515420 63466 515432
rect 92566 515420 92572 515432
rect 63460 515392 92572 515420
rect 63460 515380 63466 515392
rect 92566 515380 92572 515392
rect 92624 515380 92630 515432
rect 147582 515380 147588 515432
rect 147640 515420 147646 515432
rect 213178 515420 213184 515432
rect 147640 515392 213184 515420
rect 147640 515380 147646 515392
rect 213178 515380 213184 515392
rect 213236 515380 213242 515432
rect 233326 515380 233332 515432
rect 233384 515420 233390 515432
rect 251450 515420 251456 515432
rect 233384 515392 251456 515420
rect 233384 515380 233390 515392
rect 251450 515380 251456 515392
rect 251508 515380 251514 515432
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 193490 514088 193496 514140
rect 193548 514128 193554 514140
rect 202874 514128 202880 514140
rect 193548 514100 202880 514128
rect 193548 514088 193554 514100
rect 202874 514088 202880 514100
rect 202932 514088 202938 514140
rect 153010 514020 153016 514072
rect 153068 514060 153074 514072
rect 251266 514060 251272 514072
rect 153068 514032 251272 514060
rect 153068 514020 153074 514032
rect 251266 514020 251272 514032
rect 251324 514020 251330 514072
rect 50982 513272 50988 513324
rect 51040 513312 51046 513324
rect 169202 513312 169208 513324
rect 51040 513284 169208 513312
rect 51040 513272 51046 513284
rect 169202 513272 169208 513284
rect 169260 513272 169266 513324
rect 177390 512592 177396 512644
rect 177448 512632 177454 512644
rect 208394 512632 208400 512644
rect 177448 512604 208400 512632
rect 177448 512592 177454 512604
rect 208394 512592 208400 512604
rect 208452 512592 208458 512644
rect 186222 511232 186228 511284
rect 186280 511272 186286 511284
rect 205634 511272 205640 511284
rect 186280 511244 205640 511272
rect 186280 511232 186286 511244
rect 205634 511232 205640 511244
rect 205692 511232 205698 511284
rect 213178 511232 213184 511284
rect 213236 511272 213242 511284
rect 230474 511272 230480 511284
rect 213236 511244 230480 511272
rect 213236 511232 213242 511244
rect 230474 511232 230480 511244
rect 230532 511232 230538 511284
rect 187510 510892 187516 510944
rect 187568 510932 187574 510944
rect 191926 510932 191932 510944
rect 187568 510904 191932 510932
rect 187568 510892 187574 510904
rect 191926 510892 191932 510904
rect 191984 510892 191990 510944
rect 204990 509940 204996 509992
rect 205048 509980 205054 509992
rect 253198 509980 253204 509992
rect 205048 509952 253204 509980
rect 205048 509940 205054 509952
rect 253198 509940 253204 509952
rect 253256 509940 253262 509992
rect 146202 509872 146208 509924
rect 146260 509912 146266 509924
rect 205082 509912 205088 509924
rect 146260 509884 205088 509912
rect 146260 509872 146266 509884
rect 205082 509872 205088 509884
rect 205140 509872 205146 509924
rect 76006 509192 76012 509244
rect 76064 509232 76070 509244
rect 212442 509232 212448 509244
rect 76064 509204 212448 509232
rect 76064 509192 76070 509204
rect 212442 509192 212448 509204
rect 212500 509192 212506 509244
rect 212442 508512 212448 508564
rect 212500 508552 212506 508564
rect 222194 508552 222200 508564
rect 212500 508524 222200 508552
rect 212500 508512 212506 508524
rect 222194 508512 222200 508524
rect 222252 508512 222258 508564
rect 76006 508308 76012 508360
rect 76064 508348 76070 508360
rect 76558 508348 76564 508360
rect 76064 508320 76564 508348
rect 76064 508308 76070 508320
rect 76558 508308 76564 508320
rect 76616 508308 76622 508360
rect 206370 507152 206376 507204
rect 206428 507192 206434 507204
rect 258074 507192 258080 507204
rect 206428 507164 258080 507192
rect 206428 507152 206434 507164
rect 258074 507152 258080 507164
rect 258132 507152 258138 507204
rect 143258 507084 143264 507136
rect 143316 507124 143322 507136
rect 247678 507124 247684 507136
rect 143316 507096 247684 507124
rect 143316 507084 143322 507096
rect 247678 507084 247684 507096
rect 247736 507084 247742 507136
rect 169478 505724 169484 505776
rect 169536 505764 169542 505776
rect 254210 505764 254216 505776
rect 169536 505736 254216 505764
rect 169536 505724 169542 505736
rect 254210 505724 254216 505736
rect 254268 505724 254274 505776
rect 136542 504432 136548 504484
rect 136600 504472 136606 504484
rect 195974 504472 195980 504484
rect 136600 504444 195980 504472
rect 136600 504432 136606 504444
rect 195974 504432 195980 504444
rect 196032 504432 196038 504484
rect 168098 504364 168104 504416
rect 168156 504404 168162 504416
rect 232498 504404 232504 504416
rect 168156 504376 232504 504404
rect 168156 504364 168162 504376
rect 232498 504364 232504 504376
rect 232556 504364 232562 504416
rect 237374 504364 237380 504416
rect 237432 504404 237438 504416
rect 253198 504404 253204 504416
rect 237432 504376 253204 504404
rect 237432 504364 237438 504376
rect 253198 504364 253204 504376
rect 253256 504364 253262 504416
rect 173526 502936 173532 502988
rect 173584 502976 173590 502988
rect 244458 502976 244464 502988
rect 173584 502948 244464 502976
rect 173584 502936 173590 502948
rect 244458 502936 244464 502948
rect 244516 502936 244522 502988
rect 170766 501576 170772 501628
rect 170824 501616 170830 501628
rect 253934 501616 253940 501628
rect 170824 501588 253940 501616
rect 170824 501576 170830 501588
rect 253934 501576 253940 501588
rect 253992 501576 253998 501628
rect 210418 500284 210424 500336
rect 210476 500324 210482 500336
rect 253290 500324 253296 500336
rect 210476 500296 253296 500324
rect 210476 500284 210482 500296
rect 253290 500284 253296 500296
rect 253348 500284 253354 500336
rect 161198 500216 161204 500268
rect 161256 500256 161262 500268
rect 217318 500256 217324 500268
rect 161256 500228 217324 500256
rect 161256 500216 161262 500228
rect 217318 500216 217324 500228
rect 217376 500216 217382 500268
rect 186958 498856 186964 498908
rect 187016 498896 187022 498908
rect 216766 498896 216772 498908
rect 187016 498868 216772 498896
rect 187016 498856 187022 498868
rect 216766 498856 216772 498868
rect 216824 498856 216830 498908
rect 162670 498788 162676 498840
rect 162728 498828 162734 498840
rect 195238 498828 195244 498840
rect 162728 498800 195244 498828
rect 162728 498788 162734 498800
rect 195238 498788 195244 498800
rect 195296 498788 195302 498840
rect 233878 497496 233884 497548
rect 233936 497536 233942 497548
rect 277854 497536 277860 497548
rect 233936 497508 277860 497536
rect 233936 497496 233942 497508
rect 277854 497496 277860 497508
rect 277912 497496 277918 497548
rect 172238 497428 172244 497480
rect 172296 497468 172302 497480
rect 250438 497468 250444 497480
rect 172296 497440 250444 497468
rect 172296 497428 172302 497440
rect 250438 497428 250444 497440
rect 250496 497428 250502 497480
rect 187418 496136 187424 496188
rect 187476 496176 187482 496188
rect 214650 496176 214656 496188
rect 187476 496148 214656 496176
rect 187476 496136 187482 496148
rect 214650 496136 214656 496148
rect 214708 496136 214714 496188
rect 217318 496136 217324 496188
rect 217376 496176 217382 496188
rect 231210 496176 231216 496188
rect 217376 496148 231216 496176
rect 217376 496136 217382 496148
rect 231210 496136 231216 496148
rect 231268 496136 231274 496188
rect 108942 496068 108948 496120
rect 109000 496108 109006 496120
rect 277670 496108 277676 496120
rect 109000 496080 277676 496108
rect 109000 496068 109006 496080
rect 277670 496068 277676 496080
rect 277728 496068 277734 496120
rect 108298 495456 108304 495508
rect 108356 495496 108362 495508
rect 108942 495496 108948 495508
rect 108356 495468 108948 495496
rect 108356 495456 108362 495468
rect 108942 495456 108948 495468
rect 109000 495456 109006 495508
rect 185578 494776 185584 494828
rect 185636 494816 185642 494828
rect 214006 494816 214012 494828
rect 185636 494788 214012 494816
rect 185636 494776 185642 494788
rect 214006 494776 214012 494788
rect 214064 494776 214070 494828
rect 220906 494776 220912 494828
rect 220964 494816 220970 494828
rect 256786 494816 256792 494828
rect 220964 494788 256792 494816
rect 220964 494776 220970 494788
rect 256786 494776 256792 494788
rect 256844 494776 256850 494828
rect 154482 494708 154488 494760
rect 154540 494748 154546 494760
rect 222930 494748 222936 494760
rect 154540 494720 222936 494748
rect 154540 494708 154546 494720
rect 222930 494708 222936 494720
rect 222988 494708 222994 494760
rect 97994 492668 98000 492720
rect 98052 492708 98058 492720
rect 210234 492708 210240 492720
rect 98052 492680 210240 492708
rect 98052 492668 98058 492680
rect 210234 492668 210240 492680
rect 210292 492708 210298 492720
rect 210510 492708 210516 492720
rect 210292 492680 210516 492708
rect 210292 492668 210298 492680
rect 210510 492668 210516 492680
rect 210568 492668 210574 492720
rect 157058 491988 157064 492040
rect 157116 492028 157122 492040
rect 171778 492028 171784 492040
rect 157116 492000 171784 492028
rect 157116 491988 157122 492000
rect 171778 491988 171784 492000
rect 171836 491988 171842 492040
rect 165522 491920 165528 491972
rect 165580 491960 165586 491972
rect 197354 491960 197360 491972
rect 165580 491932 197360 491960
rect 165580 491920 165586 491932
rect 197354 491920 197360 491932
rect 197412 491920 197418 491972
rect 227622 491920 227628 491972
rect 227680 491960 227686 491972
rect 248414 491960 248420 491972
rect 227680 491932 248420 491960
rect 227680 491920 227686 491932
rect 248414 491920 248420 491932
rect 248472 491920 248478 491972
rect 184750 489132 184756 489184
rect 184808 489172 184814 489184
rect 203518 489172 203524 489184
rect 184808 489144 203524 489172
rect 184808 489132 184814 489144
rect 203518 489132 203524 489144
rect 203576 489132 203582 489184
rect 222102 489132 222108 489184
rect 222160 489172 222166 489184
rect 246298 489172 246304 489184
rect 222160 489144 246304 489172
rect 222160 489132 222166 489144
rect 246298 489132 246304 489144
rect 246356 489132 246362 489184
rect 166534 487840 166540 487892
rect 166592 487880 166598 487892
rect 220078 487880 220084 487892
rect 166592 487852 220084 487880
rect 166592 487840 166598 487852
rect 220078 487840 220084 487852
rect 220136 487840 220142 487892
rect 187510 487772 187516 487824
rect 187568 487812 187574 487824
rect 251818 487812 251824 487824
rect 187568 487784 251824 487812
rect 187568 487772 187574 487784
rect 251818 487772 251824 487784
rect 251876 487772 251882 487824
rect 235994 486684 236000 486736
rect 236052 486724 236058 486736
rect 238110 486724 238116 486736
rect 236052 486696 238116 486724
rect 236052 486684 236058 486696
rect 238110 486684 238116 486696
rect 238168 486684 238174 486736
rect 210510 486480 210516 486532
rect 210568 486520 210574 486532
rect 232498 486520 232504 486532
rect 210568 486492 232504 486520
rect 210568 486480 210574 486492
rect 232498 486480 232504 486492
rect 232556 486480 232562 486532
rect 160002 486412 160008 486464
rect 160060 486452 160066 486464
rect 184658 486452 184664 486464
rect 160060 486424 184664 486452
rect 160060 486412 160066 486424
rect 184658 486412 184664 486424
rect 184716 486452 184722 486464
rect 218146 486452 218152 486464
rect 184716 486424 218152 486452
rect 184716 486412 184722 486424
rect 218146 486412 218152 486424
rect 218204 486412 218210 486464
rect 199470 485052 199476 485104
rect 199528 485092 199534 485104
rect 241606 485092 241612 485104
rect 199528 485064 241612 485092
rect 199528 485052 199534 485064
rect 241606 485052 241612 485064
rect 241664 485052 241670 485104
rect 155678 484440 155684 484492
rect 155736 484480 155742 484492
rect 182910 484480 182916 484492
rect 155736 484452 182916 484480
rect 155736 484440 155742 484452
rect 182910 484440 182916 484452
rect 182968 484480 182974 484492
rect 183370 484480 183376 484492
rect 182968 484452 183376 484480
rect 182968 484440 182974 484452
rect 183370 484440 183376 484452
rect 183428 484440 183434 484492
rect 122742 484372 122748 484424
rect 122800 484412 122806 484424
rect 223574 484412 223580 484424
rect 122800 484384 223580 484412
rect 122800 484372 122806 484384
rect 223574 484372 223580 484384
rect 223632 484372 223638 484424
rect 183370 484304 183376 484356
rect 183428 484344 183434 484356
rect 579798 484344 579804 484356
rect 183428 484316 579804 484344
rect 183428 484304 183434 484316
rect 579798 484304 579804 484316
rect 579856 484304 579862 484356
rect 178954 483624 178960 483676
rect 179012 483664 179018 483676
rect 195422 483664 195428 483676
rect 179012 483636 195428 483664
rect 179012 483624 179018 483636
rect 195422 483624 195428 483636
rect 195480 483624 195486 483676
rect 233234 483624 233240 483676
rect 233292 483664 233298 483676
rect 249794 483664 249800 483676
rect 233292 483636 249800 483664
rect 233292 483624 233298 483636
rect 249794 483624 249800 483636
rect 249852 483624 249858 483676
rect 242894 482944 242900 482996
rect 242952 482984 242958 482996
rect 243538 482984 243544 482996
rect 242952 482956 243544 482984
rect 242952 482944 242958 482956
rect 243538 482944 243544 482956
rect 243596 482944 243602 482996
rect 177482 482264 177488 482316
rect 177540 482304 177546 482316
rect 217318 482304 217324 482316
rect 177540 482276 217324 482304
rect 177540 482264 177546 482276
rect 217318 482264 217324 482276
rect 217376 482264 217382 482316
rect 239398 482264 239404 482316
rect 239456 482304 239462 482316
rect 276198 482304 276204 482316
rect 239456 482276 276204 482304
rect 239456 482264 239462 482276
rect 276198 482264 276204 482276
rect 276256 482264 276262 482316
rect 133782 481652 133788 481704
rect 133840 481692 133846 481704
rect 242894 481692 242900 481704
rect 133840 481664 242900 481692
rect 133840 481652 133846 481664
rect 242894 481652 242900 481664
rect 242952 481652 242958 481704
rect 181898 480292 181904 480344
rect 181956 480332 181962 480344
rect 267918 480332 267924 480344
rect 181956 480304 267924 480332
rect 181956 480292 181962 480304
rect 267918 480292 267924 480304
rect 267976 480292 267982 480344
rect 126238 480224 126244 480276
rect 126296 480264 126302 480276
rect 240778 480264 240784 480276
rect 126296 480236 240784 480264
rect 126296 480224 126302 480236
rect 240778 480224 240784 480236
rect 240836 480224 240842 480276
rect 176378 479476 176384 479528
rect 176436 479516 176442 479528
rect 213914 479516 213920 479528
rect 176436 479488 213920 479516
rect 176436 479476 176442 479488
rect 213914 479476 213920 479488
rect 213972 479476 213978 479528
rect 218054 479476 218060 479528
rect 218112 479516 218118 479528
rect 254118 479516 254124 479528
rect 218112 479488 254124 479516
rect 218112 479476 218118 479488
rect 254118 479476 254124 479488
rect 254176 479476 254182 479528
rect 132402 478932 132408 478984
rect 132460 478972 132466 478984
rect 199470 478972 199476 478984
rect 132460 478944 199476 478972
rect 132460 478932 132466 478944
rect 199470 478932 199476 478944
rect 199528 478932 199534 478984
rect 198734 478864 198740 478916
rect 198792 478904 198798 478916
rect 199378 478904 199384 478916
rect 198792 478876 199384 478904
rect 198792 478864 198798 478876
rect 199378 478864 199384 478876
rect 199436 478904 199442 478916
rect 215294 478904 215300 478916
rect 199436 478876 215300 478904
rect 199436 478864 199442 478876
rect 215294 478864 215300 478876
rect 215352 478864 215358 478916
rect 148778 478184 148784 478236
rect 148836 478224 148842 478236
rect 198734 478224 198740 478236
rect 148836 478196 198740 478224
rect 148836 478184 148842 478196
rect 198734 478184 198740 478196
rect 198792 478184 198798 478236
rect 111058 478116 111064 478168
rect 111116 478156 111122 478168
rect 251450 478156 251456 478168
rect 111116 478128 251456 478156
rect 111116 478116 111122 478128
rect 251450 478116 251456 478128
rect 251508 478116 251514 478168
rect 110414 477504 110420 477556
rect 110472 477544 110478 477556
rect 111058 477544 111064 477556
rect 110472 477516 111064 477544
rect 110472 477504 110478 477516
rect 111058 477504 111064 477516
rect 111116 477504 111122 477556
rect 251450 477504 251456 477556
rect 251508 477544 251514 477556
rect 251910 477544 251916 477556
rect 251508 477516 251916 477544
rect 251508 477504 251514 477516
rect 251910 477504 251916 477516
rect 251968 477504 251974 477556
rect 85482 476756 85488 476808
rect 85540 476796 85546 476808
rect 94130 476796 94136 476808
rect 85540 476768 94136 476796
rect 85540 476756 85546 476768
rect 94130 476756 94136 476768
rect 94188 476756 94194 476808
rect 224954 476756 224960 476808
rect 225012 476796 225018 476808
rect 269758 476796 269764 476808
rect 225012 476768 269764 476796
rect 225012 476756 225018 476768
rect 269758 476756 269764 476768
rect 269816 476756 269822 476808
rect 198734 476552 198740 476604
rect 198792 476592 198798 476604
rect 199470 476592 199476 476604
rect 198792 476564 199476 476592
rect 198792 476552 198798 476564
rect 199470 476552 199476 476564
rect 199528 476552 199534 476604
rect 141418 476076 141424 476128
rect 141476 476116 141482 476128
rect 258258 476116 258264 476128
rect 141476 476088 258264 476116
rect 141476 476076 141482 476088
rect 258258 476076 258264 476088
rect 258316 476076 258322 476128
rect 3326 475328 3332 475380
rect 3384 475368 3390 475380
rect 43438 475368 43444 475380
rect 3384 475340 43444 475368
rect 3384 475328 3390 475340
rect 43438 475328 43444 475340
rect 43496 475328 43502 475380
rect 206462 475328 206468 475380
rect 206520 475368 206526 475380
rect 222838 475368 222844 475380
rect 206520 475340 222844 475368
rect 206520 475328 206526 475340
rect 222838 475328 222844 475340
rect 222896 475328 222902 475380
rect 226334 474784 226340 474836
rect 226392 474824 226398 474836
rect 226978 474824 226984 474836
rect 226392 474796 226984 474824
rect 226392 474784 226398 474796
rect 226978 474784 226984 474796
rect 227036 474824 227042 474836
rect 302234 474824 302240 474836
rect 227036 474796 302240 474824
rect 227036 474784 227042 474796
rect 302234 474784 302240 474796
rect 302292 474784 302298 474836
rect 164050 474716 164056 474768
rect 164108 474756 164114 474768
rect 251358 474756 251364 474768
rect 164108 474728 251364 474756
rect 164108 474716 164114 474728
rect 251358 474716 251364 474728
rect 251416 474716 251422 474768
rect 146938 474648 146944 474700
rect 146996 474688 147002 474700
rect 147398 474688 147404 474700
rect 146996 474660 147404 474688
rect 146996 474648 147002 474660
rect 147398 474648 147404 474660
rect 147456 474648 147462 474700
rect 146938 473424 146944 473476
rect 146996 473464 147002 473476
rect 253474 473464 253480 473476
rect 146996 473436 253480 473464
rect 146996 473424 147002 473436
rect 253474 473424 253480 473436
rect 253532 473424 253538 473476
rect 108850 473356 108856 473408
rect 108908 473396 108914 473408
rect 249058 473396 249064 473408
rect 108908 473368 249064 473396
rect 108908 473356 108914 473368
rect 249058 473356 249064 473368
rect 249116 473356 249122 473408
rect 93946 472608 93952 472660
rect 94004 472648 94010 472660
rect 94590 472648 94596 472660
rect 94004 472620 94596 472648
rect 94004 472608 94010 472620
rect 94590 472608 94596 472620
rect 94648 472648 94654 472660
rect 209774 472648 209780 472660
rect 94648 472620 209780 472648
rect 94648 472608 94654 472620
rect 209774 472608 209780 472620
rect 209832 472608 209838 472660
rect 217318 472608 217324 472660
rect 217376 472648 217382 472660
rect 269206 472648 269212 472660
rect 217376 472620 269212 472648
rect 217376 472608 217382 472620
rect 269206 472608 269212 472620
rect 269264 472608 269270 472660
rect 287054 472608 287060 472660
rect 287112 472648 287118 472660
rect 287606 472648 287612 472660
rect 287112 472620 287612 472648
rect 287112 472608 287118 472620
rect 287606 472608 287612 472620
rect 287664 472648 287670 472660
rect 582466 472648 582472 472660
rect 287664 472620 582472 472648
rect 287664 472608 287670 472620
rect 582466 472608 582472 472620
rect 582524 472608 582530 472660
rect 151078 471996 151084 472048
rect 151136 472036 151142 472048
rect 186038 472036 186044 472048
rect 151136 472008 186044 472036
rect 151136 471996 151142 472008
rect 186038 471996 186044 472008
rect 186096 472036 186102 472048
rect 229094 472036 229100 472048
rect 186096 472008 229100 472036
rect 186096 471996 186102 472008
rect 229094 471996 229100 472008
rect 229152 471996 229158 472048
rect 102134 471928 102140 471980
rect 102192 471968 102198 471980
rect 102778 471968 102784 471980
rect 102192 471940 102784 471968
rect 102192 471928 102198 471940
rect 102778 471928 102784 471940
rect 102836 471928 102842 471980
rect 79962 471248 79968 471300
rect 80020 471288 80026 471300
rect 101398 471288 101404 471300
rect 80020 471260 101404 471288
rect 80020 471248 80026 471260
rect 101398 471248 101404 471260
rect 101456 471248 101462 471300
rect 246942 471248 246948 471300
rect 247000 471288 247006 471300
rect 249702 471288 249708 471300
rect 247000 471260 249708 471288
rect 247000 471248 247006 471260
rect 249702 471248 249708 471260
rect 249760 471288 249766 471300
rect 287054 471288 287060 471300
rect 249760 471260 287060 471288
rect 249760 471248 249766 471260
rect 287054 471248 287060 471260
rect 287112 471248 287118 471300
rect 251174 471112 251180 471164
rect 251232 471152 251238 471164
rect 251818 471152 251824 471164
rect 251232 471124 251824 471152
rect 251232 471112 251238 471124
rect 251818 471112 251824 471124
rect 251876 471112 251882 471164
rect 135898 470636 135904 470688
rect 135956 470676 135962 470688
rect 251174 470676 251180 470688
rect 135956 470648 251180 470676
rect 135956 470636 135962 470648
rect 251174 470636 251180 470648
rect 251232 470636 251238 470688
rect 102134 470568 102140 470620
rect 102192 470608 102198 470620
rect 240226 470608 240232 470620
rect 102192 470580 240232 470608
rect 102192 470568 102198 470580
rect 240226 470568 240232 470580
rect 240284 470568 240290 470620
rect 180610 469820 180616 469872
rect 180668 469860 180674 469872
rect 206278 469860 206284 469872
rect 180668 469832 206284 469860
rect 180668 469820 180674 469832
rect 206278 469820 206284 469832
rect 206336 469820 206342 469872
rect 228450 469820 228456 469872
rect 228508 469860 228514 469872
rect 239398 469860 239404 469872
rect 228508 469832 239404 469860
rect 228508 469820 228514 469832
rect 239398 469820 239404 469832
rect 239456 469820 239462 469872
rect 174538 469208 174544 469260
rect 174596 469248 174602 469260
rect 174998 469248 175004 469260
rect 174596 469220 175004 469248
rect 174596 469208 174602 469220
rect 174998 469208 175004 469220
rect 175056 469248 175062 469260
rect 242158 469248 242164 469260
rect 175056 469220 242164 469248
rect 175056 469208 175062 469220
rect 242158 469208 242164 469220
rect 242216 469208 242222 469260
rect 241422 469140 241428 469192
rect 241480 469180 241486 469192
rect 259546 469180 259552 469192
rect 241480 469152 259552 469180
rect 241480 469140 241486 469152
rect 259546 469140 259552 469152
rect 259604 469140 259610 469192
rect 195330 468528 195336 468580
rect 195388 468568 195394 468580
rect 213178 468568 213184 468580
rect 195388 468540 213184 468568
rect 195388 468528 195394 468540
rect 213178 468528 213184 468540
rect 213236 468528 213242 468580
rect 223574 468528 223580 468580
rect 223632 468568 223638 468580
rect 246942 468568 246948 468580
rect 223632 468540 246948 468568
rect 223632 468528 223638 468540
rect 246942 468528 246948 468540
rect 247000 468528 247006 468580
rect 79318 468460 79324 468512
rect 79376 468500 79382 468512
rect 91186 468500 91192 468512
rect 79376 468472 91192 468500
rect 79376 468460 79382 468472
rect 91186 468460 91192 468472
rect 91244 468460 91250 468512
rect 93854 468460 93860 468512
rect 93912 468500 93918 468512
rect 160738 468500 160744 468512
rect 93912 468472 160744 468500
rect 93912 468460 93918 468472
rect 160738 468460 160744 468472
rect 160796 468500 160802 468512
rect 227714 468500 227720 468512
rect 160796 468472 227720 468500
rect 160796 468460 160802 468472
rect 227714 468460 227720 468472
rect 227772 468460 227778 468512
rect 240226 468460 240232 468512
rect 240284 468500 240290 468512
rect 241422 468500 241428 468512
rect 240284 468472 241428 468500
rect 240284 468460 240290 468472
rect 241422 468460 241428 468472
rect 241480 468460 241486 468512
rect 197354 467100 197360 467152
rect 197412 467140 197418 467152
rect 255498 467140 255504 467152
rect 197412 467112 255504 467140
rect 197412 467100 197418 467112
rect 255498 467100 255504 467112
rect 255556 467100 255562 467152
rect 140590 466488 140596 466540
rect 140648 466528 140654 466540
rect 204254 466528 204260 466540
rect 140648 466500 204260 466528
rect 140648 466488 140654 466500
rect 204254 466488 204260 466500
rect 204312 466488 204318 466540
rect 68922 466420 68928 466472
rect 68980 466460 68986 466472
rect 188338 466460 188344 466472
rect 68980 466432 188344 466460
rect 68980 466420 68986 466432
rect 188338 466420 188344 466432
rect 188396 466420 188402 466472
rect 224954 466420 224960 466472
rect 225012 466460 225018 466472
rect 226242 466460 226248 466472
rect 225012 466432 226248 466460
rect 225012 466420 225018 466432
rect 226242 466420 226248 466432
rect 226300 466460 226306 466472
rect 299566 466460 299572 466472
rect 226300 466432 299572 466460
rect 226300 466420 226306 466432
rect 299566 466420 299572 466432
rect 299624 466420 299630 466472
rect 158438 465672 158444 465724
rect 158496 465712 158502 465724
rect 165062 465712 165068 465724
rect 158496 465684 165068 465712
rect 158496 465672 158502 465684
rect 165062 465672 165068 465684
rect 165120 465672 165126 465724
rect 183278 465672 183284 465724
rect 183336 465712 183342 465724
rect 191926 465712 191932 465724
rect 183336 465684 191932 465712
rect 183336 465672 183342 465684
rect 191926 465672 191932 465684
rect 191984 465672 191990 465724
rect 193030 465672 193036 465724
rect 193088 465712 193094 465724
rect 212718 465712 212724 465724
rect 193088 465684 212724 465712
rect 193088 465672 193094 465684
rect 212718 465672 212724 465684
rect 212776 465672 212782 465724
rect 94498 465536 94504 465588
rect 94556 465576 94562 465588
rect 95142 465576 95148 465588
rect 94556 465548 95148 465576
rect 94556 465536 94562 465548
rect 95142 465536 95148 465548
rect 95200 465536 95206 465588
rect 95142 465060 95148 465112
rect 95200 465100 95206 465112
rect 216674 465100 216680 465112
rect 95200 465072 216680 465100
rect 95200 465060 95206 465072
rect 216674 465060 216680 465072
rect 216732 465060 216738 465112
rect 237374 465060 237380 465112
rect 237432 465100 237438 465112
rect 238018 465100 238024 465112
rect 237432 465072 238024 465100
rect 237432 465060 237438 465072
rect 238018 465060 238024 465072
rect 238076 465100 238082 465112
rect 289998 465100 290004 465112
rect 238076 465072 290004 465100
rect 238076 465060 238082 465072
rect 289998 465060 290004 465072
rect 290056 465060 290062 465112
rect 201494 464992 201500 465044
rect 201552 465032 201558 465044
rect 207106 465032 207112 465044
rect 201552 465004 207112 465032
rect 201552 464992 201558 465004
rect 207106 464992 207112 465004
rect 207164 464992 207170 465044
rect 77294 464312 77300 464364
rect 77352 464352 77358 464364
rect 110506 464352 110512 464364
rect 77352 464324 110512 464352
rect 77352 464312 77358 464324
rect 110506 464312 110512 464324
rect 110564 464312 110570 464364
rect 130378 464312 130384 464364
rect 130436 464352 130442 464364
rect 197354 464352 197360 464364
rect 130436 464324 197360 464352
rect 130436 464312 130442 464324
rect 197354 464312 197360 464324
rect 197412 464312 197418 464364
rect 273898 464312 273904 464364
rect 273956 464352 273962 464364
rect 280246 464352 280252 464364
rect 273956 464324 280252 464352
rect 273956 464312 273962 464324
rect 280246 464312 280252 464324
rect 280304 464312 280310 464364
rect 165614 464176 165620 464228
rect 165672 464216 165678 464228
rect 166442 464216 166448 464228
rect 165672 464188 166448 464216
rect 165672 464176 165678 464188
rect 166442 464176 166448 464188
rect 166500 464176 166506 464228
rect 226334 463768 226340 463820
rect 226392 463808 226398 463820
rect 227622 463808 227628 463820
rect 226392 463780 227628 463808
rect 226392 463768 226398 463780
rect 227622 463768 227628 463780
rect 227680 463808 227686 463820
rect 274726 463808 274732 463820
rect 227680 463780 274732 463808
rect 227680 463768 227686 463780
rect 274726 463768 274732 463780
rect 274784 463768 274790 463820
rect 106274 463700 106280 463752
rect 106332 463740 106338 463752
rect 165614 463740 165620 463752
rect 106332 463712 165620 463740
rect 106332 463700 106338 463712
rect 165614 463700 165620 463712
rect 165672 463700 165678 463752
rect 167638 463700 167644 463752
rect 167696 463740 167702 463752
rect 248414 463740 248420 463752
rect 167696 463712 248420 463740
rect 167696 463700 167702 463712
rect 248414 463700 248420 463712
rect 248472 463740 248478 463752
rect 248598 463740 248604 463752
rect 248472 463712 248604 463740
rect 248472 463700 248478 463712
rect 248598 463700 248604 463712
rect 248656 463700 248662 463752
rect 204254 463632 204260 463684
rect 204312 463672 204318 463684
rect 273438 463672 273444 463684
rect 204312 463644 273444 463672
rect 204312 463632 204318 463644
rect 273438 463632 273444 463644
rect 273496 463632 273502 463684
rect 87598 462952 87604 463004
rect 87656 462992 87662 463004
rect 104894 462992 104900 463004
rect 87656 462964 104900 462992
rect 87656 462952 87662 462964
rect 104894 462952 104900 462964
rect 104952 462952 104958 463004
rect 190270 462952 190276 463004
rect 190328 462992 190334 463004
rect 204990 462992 204996 463004
rect 190328 462964 204996 462992
rect 190328 462952 190334 462964
rect 204990 462952 204996 462964
rect 205048 462952 205054 463004
rect 3418 462408 3424 462460
rect 3476 462448 3482 462460
rect 7558 462448 7564 462460
rect 3476 462420 7564 462448
rect 3476 462408 3482 462420
rect 7558 462408 7564 462420
rect 7616 462408 7622 462460
rect 104894 462340 104900 462392
rect 104952 462380 104958 462392
rect 242986 462380 242992 462392
rect 104952 462352 242992 462380
rect 104952 462340 104958 462352
rect 242986 462340 242992 462352
rect 243044 462340 243050 462392
rect 82814 462272 82820 462324
rect 82872 462312 82878 462324
rect 108850 462312 108856 462324
rect 82872 462284 108856 462312
rect 82872 462272 82878 462284
rect 108850 462272 108856 462284
rect 108908 462312 108914 462324
rect 109034 462312 109040 462324
rect 108908 462284 109040 462312
rect 108908 462272 108914 462284
rect 109034 462272 109040 462284
rect 109092 462272 109098 462324
rect 251174 462272 251180 462324
rect 251232 462312 251238 462324
rect 251910 462312 251916 462324
rect 251232 462284 251916 462312
rect 251232 462272 251238 462284
rect 251910 462272 251916 462284
rect 251968 462272 251974 462324
rect 216674 461660 216680 461712
rect 216732 461700 216738 461712
rect 231854 461700 231860 461712
rect 216732 461672 231860 461700
rect 216732 461660 216738 461672
rect 231854 461660 231860 461672
rect 231912 461660 231918 461712
rect 67634 461592 67640 461644
rect 67692 461632 67698 461644
rect 83458 461632 83464 461644
rect 67692 461604 83464 461632
rect 67692 461592 67698 461604
rect 83458 461592 83464 461604
rect 83516 461592 83522 461644
rect 110506 461592 110512 461644
rect 110564 461632 110570 461644
rect 117314 461632 117320 461644
rect 110564 461604 117320 461632
rect 110564 461592 110570 461604
rect 117314 461592 117320 461604
rect 117372 461592 117378 461644
rect 213822 461592 213828 461644
rect 213880 461632 213886 461644
rect 270586 461632 270592 461644
rect 213880 461604 270592 461632
rect 213880 461592 213886 461604
rect 270586 461592 270592 461604
rect 270644 461592 270650 461644
rect 216674 461524 216680 461576
rect 216732 461564 216738 461576
rect 217318 461564 217324 461576
rect 216732 461536 217324 461564
rect 216732 461524 216738 461536
rect 217318 461524 217324 461536
rect 217376 461524 217382 461576
rect 184658 460980 184664 461032
rect 184716 461020 184722 461032
rect 216674 461020 216680 461032
rect 184716 460992 216680 461020
rect 184716 460980 184722 460992
rect 216674 460980 216680 460992
rect 216732 460980 216738 461032
rect 104802 460912 104808 460964
rect 104860 460952 104866 460964
rect 188154 460952 188160 460964
rect 104860 460924 188160 460952
rect 104860 460912 104866 460924
rect 188154 460912 188160 460924
rect 188212 460912 188218 460964
rect 251174 460912 251180 460964
rect 251232 460952 251238 460964
rect 292666 460952 292672 460964
rect 251232 460924 292672 460952
rect 251232 460912 251238 460924
rect 292666 460912 292672 460924
rect 292724 460912 292730 460964
rect 66162 460164 66168 460216
rect 66220 460204 66226 460216
rect 85666 460204 85672 460216
rect 66220 460176 85672 460204
rect 66220 460164 66226 460176
rect 85666 460164 85672 460176
rect 85724 460164 85730 460216
rect 86218 460164 86224 460216
rect 86276 460204 86282 460216
rect 114554 460204 114560 460216
rect 86276 460176 114560 460204
rect 86276 460164 86282 460176
rect 114554 460164 114560 460176
rect 114612 460164 114618 460216
rect 142798 460164 142804 460216
rect 142856 460204 142862 460216
rect 249794 460204 249800 460216
rect 142856 460176 249800 460204
rect 142856 460164 142862 460176
rect 249794 460164 249800 460176
rect 249852 460204 249858 460216
rect 259546 460204 259552 460216
rect 249852 460176 259552 460204
rect 249852 460164 249858 460176
rect 259546 460164 259552 460176
rect 259604 460164 259610 460216
rect 112438 459552 112444 459604
rect 112496 459592 112502 459604
rect 113082 459592 113088 459604
rect 112496 459564 113088 459592
rect 112496 459552 112502 459564
rect 113082 459552 113088 459564
rect 113140 459592 113146 459604
rect 129642 459592 129648 459604
rect 113140 459564 129648 459592
rect 113140 459552 113146 459564
rect 129642 459552 129648 459564
rect 129700 459592 129706 459604
rect 249610 459592 249616 459604
rect 129700 459564 249616 459592
rect 129700 459552 129706 459564
rect 249610 459552 249616 459564
rect 249668 459552 249674 459604
rect 187786 459484 187792 459536
rect 187844 459524 187850 459536
rect 211798 459524 211804 459536
rect 187844 459496 211804 459524
rect 187844 459484 187850 459496
rect 211798 459484 211804 459496
rect 211856 459484 211862 459536
rect 253198 458872 253204 458924
rect 253256 458912 253262 458924
rect 262398 458912 262404 458924
rect 253256 458884 262404 458912
rect 253256 458872 253262 458884
rect 262398 458872 262404 458884
rect 262456 458872 262462 458924
rect 241514 458804 241520 458856
rect 241572 458844 241578 458856
rect 254026 458844 254032 458856
rect 241572 458816 254032 458844
rect 241572 458804 241578 458816
rect 254026 458804 254032 458816
rect 254084 458804 254090 458856
rect 276290 458668 276296 458720
rect 276348 458708 276354 458720
rect 277302 458708 277308 458720
rect 276348 458680 277308 458708
rect 276348 458668 276354 458680
rect 277302 458668 277308 458680
rect 277360 458708 277366 458720
rect 278866 458708 278872 458720
rect 277360 458680 278872 458708
rect 277360 458668 277366 458680
rect 278866 458668 278872 458680
rect 278924 458668 278930 458720
rect 160738 458260 160744 458312
rect 160796 458300 160802 458312
rect 197354 458300 197360 458312
rect 160796 458272 197360 458300
rect 160796 458260 160802 458272
rect 197354 458260 197360 458272
rect 197412 458300 197418 458312
rect 197998 458300 198004 458312
rect 197412 458272 198004 458300
rect 197412 458260 197418 458272
rect 197998 458260 198004 458272
rect 198056 458260 198062 458312
rect 75178 458192 75184 458244
rect 75236 458232 75242 458244
rect 75822 458232 75828 458244
rect 75236 458204 75828 458232
rect 75236 458192 75242 458204
rect 75822 458192 75828 458204
rect 75880 458232 75886 458244
rect 187694 458232 187700 458244
rect 75880 458204 187700 458232
rect 75880 458192 75886 458204
rect 187694 458192 187700 458204
rect 187752 458192 187758 458244
rect 100018 457444 100024 457496
rect 100076 457484 100082 457496
rect 142890 457484 142896 457496
rect 100076 457456 142896 457484
rect 100076 457444 100082 457456
rect 142890 457444 142896 457456
rect 142948 457444 142954 457496
rect 154022 457444 154028 457496
rect 154080 457484 154086 457496
rect 187602 457484 187608 457496
rect 154080 457456 187608 457484
rect 154080 457444 154086 457456
rect 187602 457444 187608 457456
rect 187660 457444 187666 457496
rect 188154 457444 188160 457496
rect 188212 457484 188218 457496
rect 246390 457484 246396 457496
rect 188212 457456 246396 457484
rect 188212 457444 188218 457456
rect 246390 457444 246396 457456
rect 246448 457444 246454 457496
rect 247494 457444 247500 457496
rect 247552 457484 247558 457496
rect 277670 457484 277676 457496
rect 247552 457456 277676 457484
rect 247552 457444 247558 457456
rect 277670 457444 277676 457456
rect 277728 457444 277734 457496
rect 156598 457376 156604 457428
rect 156656 457416 156662 457428
rect 163498 457416 163504 457428
rect 156656 457388 163504 457416
rect 156656 457376 156662 457388
rect 163498 457376 163504 457388
rect 163556 457376 163562 457428
rect 184198 456764 184204 456816
rect 184256 456804 184262 456816
rect 213270 456804 213276 456816
rect 184256 456776 213276 456804
rect 184256 456764 184262 456776
rect 213270 456764 213276 456776
rect 213328 456804 213334 456816
rect 213822 456804 213828 456816
rect 213328 456776 213828 456804
rect 213328 456764 213334 456776
rect 213822 456764 213828 456776
rect 213880 456764 213886 456816
rect 237466 456764 237472 456816
rect 237524 456804 237530 456816
rect 238110 456804 238116 456816
rect 237524 456776 238116 456804
rect 237524 456764 237530 456776
rect 238110 456764 238116 456776
rect 238168 456804 238174 456816
rect 253566 456804 253572 456816
rect 238168 456776 253572 456804
rect 238168 456764 238174 456776
rect 253566 456764 253572 456776
rect 253624 456764 253630 456816
rect 187510 456084 187516 456136
rect 187568 456124 187574 456136
rect 188338 456124 188344 456136
rect 187568 456096 188344 456124
rect 187568 456084 187574 456096
rect 188338 456084 188344 456096
rect 188396 456084 188402 456136
rect 218146 456084 218152 456136
rect 218204 456124 218210 456136
rect 218974 456124 218980 456136
rect 218204 456096 218980 456124
rect 218204 456084 218210 456096
rect 218974 456084 218980 456096
rect 219032 456084 219038 456136
rect 251266 456084 251272 456136
rect 251324 456124 251330 456136
rect 252094 456124 252100 456136
rect 251324 456096 252100 456124
rect 251324 456084 251330 456096
rect 252094 456084 252100 456096
rect 252152 456084 252158 456136
rect 187694 456016 187700 456068
rect 187752 456056 187758 456068
rect 196066 456056 196072 456068
rect 187752 456028 196072 456056
rect 187752 456016 187758 456028
rect 196066 456016 196072 456028
rect 196124 456016 196130 456068
rect 240134 456016 240140 456068
rect 240192 456056 240198 456068
rect 254210 456056 254216 456068
rect 240192 456028 254216 456056
rect 240192 456016 240198 456028
rect 254210 456016 254216 456028
rect 254268 456016 254274 456068
rect 288342 456016 288348 456068
rect 288400 456056 288406 456068
rect 580166 456056 580172 456068
rect 288400 456028 580172 456056
rect 288400 456016 288406 456028
rect 580166 456016 580172 456028
rect 580224 456016 580230 456068
rect 225046 455744 225052 455796
rect 225104 455784 225110 455796
rect 226978 455784 226984 455796
rect 225104 455756 226984 455784
rect 225104 455744 225110 455756
rect 226978 455744 226984 455756
rect 227036 455744 227042 455796
rect 82078 455404 82084 455456
rect 82136 455444 82142 455456
rect 82722 455444 82728 455456
rect 82136 455416 82728 455444
rect 82136 455404 82142 455416
rect 82722 455404 82728 455416
rect 82780 455444 82786 455456
rect 211154 455444 211160 455456
rect 82780 455416 211160 455444
rect 82780 455404 82786 455416
rect 211154 455404 211160 455416
rect 211212 455404 211218 455456
rect 233970 455404 233976 455456
rect 234028 455444 234034 455456
rect 258074 455444 258080 455456
rect 234028 455416 258080 455444
rect 234028 455404 234034 455416
rect 258074 455404 258080 455416
rect 258132 455404 258138 455456
rect 73154 455336 73160 455388
rect 73212 455376 73218 455388
rect 112990 455376 112996 455388
rect 73212 455348 112996 455376
rect 73212 455336 73218 455348
rect 112990 455336 112996 455348
rect 113048 455376 113054 455388
rect 128998 455376 129004 455388
rect 113048 455348 129004 455376
rect 113048 455336 113054 455348
rect 128998 455336 129004 455348
rect 129056 455336 129062 455388
rect 214650 455336 214656 455388
rect 214708 455376 214714 455388
rect 233988 455376 234016 455404
rect 214708 455348 234016 455376
rect 214708 455336 214714 455348
rect 242986 455336 242992 455388
rect 243044 455376 243050 455388
rect 243538 455376 243544 455388
rect 243044 455348 243544 455376
rect 243044 455336 243050 455348
rect 243538 455336 243544 455348
rect 243596 455376 243602 455388
rect 276106 455376 276112 455388
rect 243596 455348 276112 455376
rect 243596 455336 243602 455348
rect 276106 455336 276112 455348
rect 276164 455376 276170 455388
rect 276382 455376 276388 455388
rect 276164 455348 276388 455376
rect 276164 455336 276170 455348
rect 276382 455336 276388 455348
rect 276440 455336 276446 455388
rect 221642 455268 221648 455320
rect 221700 455308 221706 455320
rect 222102 455308 222108 455320
rect 221700 455280 222108 455308
rect 221700 455268 221706 455280
rect 222102 455268 222108 455280
rect 222160 455268 222166 455320
rect 63402 454656 63408 454708
rect 63460 454696 63466 454708
rect 74534 454696 74540 454708
rect 63460 454668 74540 454696
rect 63460 454656 63466 454668
rect 74534 454656 74540 454668
rect 74592 454696 74598 454708
rect 154390 454696 154396 454708
rect 74592 454668 154396 454696
rect 74592 454656 74598 454668
rect 154390 454656 154396 454668
rect 154448 454696 154454 454708
rect 178862 454696 178868 454708
rect 154448 454668 178868 454696
rect 154448 454656 154454 454668
rect 178862 454656 178868 454668
rect 178920 454656 178926 454708
rect 276382 454656 276388 454708
rect 276440 454696 276446 454708
rect 280246 454696 280252 454708
rect 276440 454668 280252 454696
rect 276440 454656 276446 454668
rect 280246 454656 280252 454668
rect 280304 454656 280310 454708
rect 188430 454112 188436 454164
rect 188488 454152 188494 454164
rect 207106 454152 207112 454164
rect 188488 454124 207112 454152
rect 188488 454112 188494 454124
rect 207106 454112 207112 454124
rect 207164 454112 207170 454164
rect 187050 454044 187056 454096
rect 187108 454084 187114 454096
rect 209866 454084 209872 454096
rect 187108 454056 209872 454084
rect 187108 454044 187114 454056
rect 209866 454044 209872 454056
rect 209924 454084 209930 454096
rect 210418 454084 210424 454096
rect 209924 454056 210424 454084
rect 209924 454044 209930 454056
rect 210418 454044 210424 454056
rect 210476 454044 210482 454096
rect 221642 454044 221648 454096
rect 221700 454084 221706 454096
rect 261110 454084 261116 454096
rect 221700 454056 261116 454084
rect 221700 454044 221706 454056
rect 261110 454044 261116 454056
rect 261168 454044 261174 454096
rect 221182 453976 221188 454028
rect 221240 454016 221246 454028
rect 223482 454016 223488 454028
rect 221240 453988 223488 454016
rect 221240 453976 221246 453988
rect 223482 453976 223488 453988
rect 223540 453976 223546 454028
rect 227806 453976 227812 454028
rect 227864 454016 227870 454028
rect 228726 454016 228732 454028
rect 227864 453988 228732 454016
rect 227864 453976 227870 453988
rect 228726 453976 228732 453988
rect 228784 453976 228790 454028
rect 249610 453976 249616 454028
rect 249668 454016 249674 454028
rect 253382 454016 253388 454028
rect 249668 453988 253388 454016
rect 249668 453976 249674 453988
rect 253382 453976 253388 453988
rect 253440 453976 253446 454028
rect 260098 453976 260104 454028
rect 260156 454016 260162 454028
rect 262306 454016 262312 454028
rect 260156 453988 262312 454016
rect 260156 453976 260162 453988
rect 262306 453976 262312 453988
rect 262364 453976 262370 454028
rect 198826 453908 198832 453960
rect 198884 453948 198890 453960
rect 200390 453948 200396 453960
rect 198884 453920 200396 453948
rect 198884 453908 198890 453920
rect 200390 453908 200396 453920
rect 200448 453908 200454 453960
rect 194502 453296 194508 453348
rect 194560 453336 194566 453348
rect 241422 453336 241428 453348
rect 194560 453308 241428 453336
rect 194560 453296 194566 453308
rect 241422 453296 241428 453308
rect 241480 453296 241486 453348
rect 122190 452684 122196 452736
rect 122248 452724 122254 452736
rect 195238 452724 195244 452736
rect 122248 452696 195244 452724
rect 122248 452684 122254 452696
rect 195238 452684 195244 452696
rect 195296 452684 195302 452736
rect 77938 452616 77944 452668
rect 77996 452656 78002 452668
rect 166442 452656 166448 452668
rect 77996 452628 166448 452656
rect 77996 452616 78002 452628
rect 166442 452616 166448 452628
rect 166500 452616 166506 452668
rect 204162 452616 204168 452668
rect 204220 452656 204226 452668
rect 218698 452656 218704 452668
rect 204220 452628 218704 452656
rect 204220 452616 204226 452628
rect 218698 452616 218704 452628
rect 218756 452616 218762 452668
rect 223022 452616 223028 452668
rect 223080 452656 223086 452668
rect 260098 452656 260104 452668
rect 223080 452628 260104 452656
rect 223080 452616 223086 452628
rect 260098 452616 260104 452628
rect 260156 452616 260162 452668
rect 75822 451868 75828 451920
rect 75880 451908 75886 451920
rect 98730 451908 98736 451920
rect 75880 451880 98736 451908
rect 75880 451868 75886 451880
rect 98730 451868 98736 451880
rect 98788 451868 98794 451920
rect 105538 451868 105544 451920
rect 105596 451908 105602 451920
rect 158806 451908 158812 451920
rect 105596 451880 158812 451908
rect 105596 451868 105602 451880
rect 158806 451868 158812 451880
rect 158864 451868 158870 451920
rect 279418 451868 279424 451920
rect 279476 451908 279482 451920
rect 287146 451908 287152 451920
rect 279476 451880 287152 451908
rect 279476 451868 279482 451880
rect 287146 451868 287152 451880
rect 287204 451868 287210 451920
rect 182174 451324 182180 451376
rect 182232 451364 182238 451376
rect 195606 451364 195612 451376
rect 182232 451336 195612 451364
rect 182232 451324 182238 451336
rect 195606 451324 195612 451336
rect 195664 451324 195670 451376
rect 227714 451324 227720 451376
rect 227772 451364 227778 451376
rect 272058 451364 272064 451376
rect 227772 451336 272064 451364
rect 227772 451324 227778 451336
rect 272058 451324 272064 451336
rect 272116 451324 272122 451376
rect 116578 451256 116584 451308
rect 116636 451296 116642 451308
rect 116636 451268 240088 451296
rect 116636 451256 116642 451268
rect 240060 451228 240088 451268
rect 240134 451256 240140 451308
rect 240192 451296 240198 451308
rect 241330 451296 241336 451308
rect 240192 451268 241336 451296
rect 240192 451256 240198 451268
rect 241330 451256 241336 451268
rect 241388 451296 241394 451308
rect 261018 451296 261024 451308
rect 241388 451268 261024 451296
rect 241388 451256 241394 451268
rect 261018 451256 261024 451268
rect 261076 451256 261082 451308
rect 240686 451228 240692 451240
rect 240060 451200 240692 451228
rect 240686 451188 240692 451200
rect 240744 451188 240750 451240
rect 251818 450984 251824 451036
rect 251876 451024 251882 451036
rect 256970 451024 256976 451036
rect 251876 450996 256976 451024
rect 251876 450984 251882 450996
rect 256970 450984 256976 450996
rect 257028 450984 257034 451036
rect 113818 450644 113824 450696
rect 113876 450684 113882 450696
rect 114462 450684 114468 450696
rect 113876 450656 114468 450684
rect 113876 450644 113882 450656
rect 114462 450644 114468 450656
rect 114520 450644 114526 450696
rect 180058 450576 180064 450628
rect 180116 450616 180122 450628
rect 188798 450616 188804 450628
rect 180116 450588 188804 450616
rect 180116 450576 180122 450588
rect 188798 450576 188804 450588
rect 188856 450576 188862 450628
rect 4798 450508 4804 450560
rect 4856 450548 4862 450560
rect 104158 450548 104164 450560
rect 4856 450520 104164 450548
rect 4856 450508 4862 450520
rect 104158 450508 104164 450520
rect 104216 450508 104222 450560
rect 184290 450508 184296 450560
rect 184348 450548 184354 450560
rect 204162 450548 204168 450560
rect 184348 450520 204168 450548
rect 184348 450508 184354 450520
rect 204162 450508 204168 450520
rect 204220 450508 204226 450560
rect 193214 450236 193220 450288
rect 193272 450276 193278 450288
rect 193490 450276 193496 450288
rect 193272 450248 193496 450276
rect 193272 450236 193278 450248
rect 193490 450236 193496 450248
rect 193548 450236 193554 450288
rect 114462 449964 114468 450016
rect 114520 450004 114526 450016
rect 172330 450004 172336 450016
rect 114520 449976 172336 450004
rect 114520 449964 114526 449976
rect 172330 449964 172336 449976
rect 172388 449964 172394 450016
rect 78674 449896 78680 449948
rect 78732 449936 78738 449948
rect 174998 449936 175004 449948
rect 78732 449908 175004 449936
rect 78732 449896 78738 449908
rect 174998 449896 175004 449908
rect 175056 449896 175062 449948
rect 188798 449896 188804 449948
rect 188856 449936 188862 449948
rect 250898 449936 250904 449948
rect 188856 449908 250904 449936
rect 188856 449896 188862 449908
rect 250898 449896 250904 449908
rect 250956 449936 250962 449948
rect 258166 449936 258172 449948
rect 250956 449908 258172 449936
rect 250956 449896 250962 449908
rect 258166 449896 258172 449908
rect 258224 449896 258230 449948
rect 192754 449760 192760 449812
rect 192812 449800 192818 449812
rect 195330 449800 195336 449812
rect 192812 449772 195336 449800
rect 192812 449760 192818 449772
rect 195330 449760 195336 449772
rect 195388 449760 195394 449812
rect 172330 449692 172336 449744
rect 172388 449732 172394 449744
rect 194502 449732 194508 449744
rect 172388 449704 194508 449732
rect 172388 449692 172394 449704
rect 194502 449692 194508 449704
rect 194560 449692 194566 449744
rect 251910 449692 251916 449744
rect 251968 449732 251974 449744
rect 251968 449704 258074 449732
rect 251968 449692 251974 449704
rect 95234 449216 95240 449268
rect 95292 449256 95298 449268
rect 151078 449256 151084 449268
rect 95292 449228 151084 449256
rect 95292 449216 95298 449228
rect 151078 449216 151084 449228
rect 151136 449216 151142 449268
rect 57882 449148 57888 449200
rect 57940 449188 57946 449200
rect 169018 449188 169024 449200
rect 57940 449160 169024 449188
rect 57940 449148 57946 449160
rect 169018 449148 169024 449160
rect 169076 449148 169082 449200
rect 258046 449188 258074 449704
rect 268010 449188 268016 449200
rect 258046 449160 268016 449188
rect 268010 449148 268016 449160
rect 268068 449148 268074 449200
rect 184842 449080 184848 449132
rect 184900 449120 184906 449132
rect 191558 449120 191564 449132
rect 184900 449092 191564 449120
rect 184900 449080 184906 449092
rect 191558 449080 191564 449092
rect 191616 449080 191622 449132
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 36538 448576 36544 448588
rect 3200 448548 36544 448576
rect 3200 448536 3206 448548
rect 36538 448536 36544 448548
rect 36596 448536 36602 448588
rect 66070 448536 66076 448588
rect 66128 448576 66134 448588
rect 70486 448576 70492 448588
rect 66128 448548 70492 448576
rect 66128 448536 66134 448548
rect 70486 448536 70492 448548
rect 70544 448536 70550 448588
rect 95142 448536 95148 448588
rect 95200 448576 95206 448588
rect 95878 448576 95884 448588
rect 95200 448548 95884 448576
rect 95200 448536 95206 448548
rect 95878 448536 95884 448548
rect 95936 448536 95942 448588
rect 177574 447856 177580 447908
rect 177632 447896 177638 447908
rect 188430 447896 188436 447908
rect 177632 447868 188436 447896
rect 177632 447856 177638 447868
rect 188430 447856 188436 447868
rect 188488 447856 188494 447908
rect 66162 447788 66168 447840
rect 66220 447828 66226 447840
rect 191558 447828 191564 447840
rect 66220 447800 191564 447828
rect 66220 447788 66226 447800
rect 191558 447788 191564 447800
rect 191616 447788 191622 447840
rect 176102 447040 176108 447092
rect 176160 447080 176166 447092
rect 176470 447080 176476 447092
rect 176160 447052 176476 447080
rect 176160 447040 176166 447052
rect 176470 447040 176476 447052
rect 176528 447080 176534 447092
rect 191006 447080 191012 447092
rect 176528 447052 191012 447080
rect 176528 447040 176534 447052
rect 191006 447040 191012 447052
rect 191064 447040 191070 447092
rect 67174 446428 67180 446480
rect 67232 446468 67238 446480
rect 165062 446468 165068 446480
rect 67232 446440 165068 446468
rect 67232 446428 67238 446440
rect 165062 446428 165068 446440
rect 165120 446428 165126 446480
rect 76650 446360 76656 446412
rect 76708 446400 76714 446412
rect 176102 446400 176108 446412
rect 76708 446372 176108 446400
rect 76708 446360 76714 446372
rect 176102 446360 176108 446372
rect 176160 446360 176166 446412
rect 255590 446360 255596 446412
rect 255648 446400 255654 446412
rect 269206 446400 269212 446412
rect 255648 446372 269212 446400
rect 255648 446360 255654 446372
rect 269206 446360 269212 446372
rect 269264 446360 269270 446412
rect 173710 445748 173716 445800
rect 173768 445788 173774 445800
rect 177298 445788 177304 445800
rect 173768 445760 177304 445788
rect 173768 445748 173774 445760
rect 177298 445748 177304 445760
rect 177356 445748 177362 445800
rect 160094 445680 160100 445732
rect 160152 445720 160158 445732
rect 160738 445720 160744 445732
rect 160152 445692 160744 445720
rect 160152 445680 160158 445692
rect 160738 445680 160744 445692
rect 160796 445680 160802 445732
rect 177316 445720 177344 445748
rect 191006 445720 191012 445732
rect 177316 445692 191012 445720
rect 191006 445680 191012 445692
rect 191064 445680 191070 445732
rect 143350 445000 143356 445052
rect 143408 445040 143414 445052
rect 184198 445040 184204 445052
rect 143408 445012 184204 445040
rect 143408 445000 143414 445012
rect 184198 445000 184204 445012
rect 184256 445000 184262 445052
rect 269758 445000 269764 445052
rect 269816 445040 269822 445052
rect 278866 445040 278872 445052
rect 269816 445012 278872 445040
rect 269816 445000 269822 445012
rect 278866 445000 278872 445012
rect 278924 445000 278930 445052
rect 83458 444456 83464 444508
rect 83516 444496 83522 444508
rect 142890 444496 142896 444508
rect 83516 444468 142896 444496
rect 83516 444456 83522 444468
rect 142890 444456 142896 444468
rect 142948 444496 142954 444508
rect 143350 444496 143356 444508
rect 142948 444468 143356 444496
rect 142948 444456 142954 444468
rect 143350 444456 143356 444468
rect 143408 444456 143414 444508
rect 72418 444388 72424 444440
rect 72476 444428 72482 444440
rect 160094 444428 160100 444440
rect 72476 444400 160100 444428
rect 72476 444388 72482 444400
rect 160094 444388 160100 444400
rect 160152 444388 160158 444440
rect 86954 444320 86960 444372
rect 87012 444360 87018 444372
rect 88242 444360 88248 444372
rect 87012 444332 88248 444360
rect 87012 444320 87018 444332
rect 88242 444320 88248 444332
rect 88300 444320 88306 444372
rect 255498 443844 255504 443896
rect 255556 443884 255562 443896
rect 255556 443856 258074 443884
rect 255556 443844 255562 443856
rect 88242 443708 88248 443760
rect 88300 443748 88306 443760
rect 184290 443748 184296 443760
rect 88300 443720 184296 443748
rect 88300 443708 88306 443720
rect 184290 443708 184296 443720
rect 184348 443708 184354 443760
rect 68922 443640 68928 443692
rect 68980 443680 68986 443692
rect 80054 443680 80060 443692
rect 68980 443652 80060 443680
rect 68980 443640 68986 443652
rect 80054 443640 80060 443652
rect 80112 443640 80118 443692
rect 184566 443640 184572 443692
rect 184624 443680 184630 443692
rect 187142 443680 187148 443692
rect 184624 443652 187148 443680
rect 184624 443640 184630 443652
rect 187142 443640 187148 443652
rect 187200 443640 187206 443692
rect 258046 443680 258074 443856
rect 258258 443680 258264 443692
rect 258046 443652 258264 443680
rect 258258 443640 258264 443652
rect 258316 443680 258322 443692
rect 269298 443680 269304 443692
rect 258316 443652 269304 443680
rect 258316 443640 258322 443652
rect 269298 443640 269304 443652
rect 269356 443640 269362 443692
rect 193030 443068 193036 443080
rect 180766 443040 193036 443068
rect 71130 442960 71136 443012
rect 71188 443000 71194 443012
rect 180766 443000 180794 443040
rect 193030 443028 193036 443040
rect 193088 443028 193094 443080
rect 71188 442972 180794 443000
rect 71188 442960 71194 442972
rect 257338 442280 257344 442332
rect 257396 442320 257402 442332
rect 263686 442320 263692 442332
rect 257396 442292 263692 442320
rect 257396 442280 257402 442292
rect 263686 442280 263692 442292
rect 263744 442280 263750 442332
rect 163958 442212 163964 442264
rect 164016 442252 164022 442264
rect 190270 442252 190276 442264
rect 164016 442224 190276 442252
rect 164016 442212 164022 442224
rect 190270 442212 190276 442224
rect 190328 442252 190334 442264
rect 191558 442252 191564 442264
rect 190328 442224 191564 442252
rect 190328 442212 190334 442224
rect 191558 442212 191564 442224
rect 191616 442212 191622 442264
rect 255498 442212 255504 442264
rect 255556 442252 255562 442264
rect 259638 442252 259644 442264
rect 255556 442224 259644 442252
rect 255556 442212 255562 442224
rect 259638 442212 259644 442224
rect 259696 442252 259702 442264
rect 285766 442252 285772 442264
rect 259696 442224 285772 442252
rect 259696 442212 259702 442224
rect 285766 442212 285772 442224
rect 285824 442212 285830 442264
rect 61838 441668 61844 441720
rect 61896 441708 61902 441720
rect 138658 441708 138664 441720
rect 61896 441680 138664 441708
rect 61896 441668 61902 441680
rect 138658 441668 138664 441680
rect 138716 441668 138722 441720
rect 68278 441600 68284 441652
rect 68336 441640 68342 441652
rect 163958 441640 163964 441652
rect 68336 441612 163964 441640
rect 68336 441600 68342 441612
rect 163958 441600 163964 441612
rect 164016 441600 164022 441652
rect 173618 441532 173624 441584
rect 173676 441572 173682 441584
rect 191558 441572 191564 441584
rect 173676 441544 191564 441572
rect 173676 441532 173682 441544
rect 191558 441532 191564 441544
rect 191616 441532 191622 441584
rect 104158 441464 104164 441516
rect 104216 441504 104222 441516
rect 174538 441504 174544 441516
rect 104216 441476 174544 441504
rect 104216 441464 104222 441476
rect 174538 441464 174544 441476
rect 174596 441464 174602 441516
rect 69750 440852 69756 440904
rect 69808 440892 69814 440904
rect 122190 440892 122196 440904
rect 69808 440864 122196 440892
rect 69808 440852 69814 440864
rect 122190 440852 122196 440864
rect 122248 440852 122254 440904
rect 190270 440852 190276 440904
rect 190328 440892 190334 440904
rect 193306 440892 193312 440904
rect 190328 440864 193312 440892
rect 190328 440852 190334 440864
rect 193306 440852 193312 440864
rect 193364 440852 193370 440904
rect 183370 440240 183376 440292
rect 183428 440280 183434 440292
rect 186958 440280 186964 440292
rect 183428 440252 186964 440280
rect 183428 440240 183434 440252
rect 186958 440240 186964 440252
rect 187016 440240 187022 440292
rect 76834 439560 76840 439612
rect 76892 439600 76898 439612
rect 89714 439600 89720 439612
rect 76892 439572 89720 439600
rect 76892 439560 76898 439572
rect 89714 439560 89720 439572
rect 89772 439560 89778 439612
rect 50982 439492 50988 439544
rect 51040 439532 51046 439544
rect 83734 439532 83740 439544
rect 51040 439504 83740 439532
rect 51040 439492 51046 439504
rect 83734 439492 83740 439504
rect 83792 439492 83798 439544
rect 255498 439492 255504 439544
rect 255556 439532 255562 439544
rect 288710 439532 288716 439544
rect 255556 439504 288716 439532
rect 255556 439492 255562 439504
rect 288710 439492 288716 439504
rect 288768 439492 288774 439544
rect 183462 438948 183468 439000
rect 183520 438988 183526 439000
rect 186958 438988 186964 439000
rect 183520 438960 186964 438988
rect 183520 438948 183526 438960
rect 186958 438948 186964 438960
rect 187016 438948 187022 439000
rect 104802 438880 104808 438932
rect 104860 438920 104866 438932
rect 107654 438920 107660 438932
rect 104860 438892 107660 438920
rect 104860 438880 104866 438892
rect 107654 438880 107660 438892
rect 107712 438880 107718 438932
rect 186038 438880 186044 438932
rect 186096 438920 186102 438932
rect 187694 438920 187700 438932
rect 186096 438892 187700 438920
rect 186096 438880 186102 438892
rect 187694 438880 187700 438892
rect 187752 438880 187758 438932
rect 147674 438812 147680 438864
rect 147732 438852 147738 438864
rect 148686 438852 148692 438864
rect 147732 438824 148692 438852
rect 147732 438812 147738 438824
rect 148686 438812 148692 438824
rect 148744 438852 148750 438864
rect 191650 438852 191656 438864
rect 148744 438824 191656 438852
rect 148744 438812 148750 438824
rect 191650 438812 191656 438824
rect 191708 438812 191714 438864
rect 255498 438812 255504 438864
rect 255556 438852 255562 438864
rect 263778 438852 263784 438864
rect 255556 438824 263784 438852
rect 255556 438812 255562 438824
rect 263778 438812 263784 438824
rect 263836 438812 263842 438864
rect 255958 438744 255964 438796
rect 256016 438784 256022 438796
rect 260190 438784 260196 438796
rect 256016 438756 260196 438784
rect 256016 438744 256022 438756
rect 260190 438744 260196 438756
rect 260248 438744 260254 438796
rect 73890 438200 73896 438252
rect 73948 438240 73954 438252
rect 77938 438240 77944 438252
rect 73948 438212 77944 438240
rect 73948 438200 73954 438212
rect 77938 438200 77944 438212
rect 77996 438200 78002 438252
rect 67358 438132 67364 438184
rect 67416 438172 67422 438184
rect 76650 438172 76656 438184
rect 67416 438144 76656 438172
rect 67416 438132 67422 438144
rect 76650 438132 76656 438144
rect 76708 438132 76714 438184
rect 81434 438132 81440 438184
rect 81492 438172 81498 438184
rect 88978 438172 88984 438184
rect 81492 438144 88984 438172
rect 81492 438132 81498 438144
rect 88978 438132 88984 438144
rect 89036 438132 89042 438184
rect 90634 438132 90640 438184
rect 90692 438172 90698 438184
rect 147674 438172 147680 438184
rect 90692 438144 147680 438172
rect 90692 438132 90698 438144
rect 147674 438132 147680 438144
rect 147732 438132 147738 438184
rect 78582 437452 78588 437504
rect 78640 437492 78646 437504
rect 176470 437492 176476 437504
rect 78640 437464 176476 437492
rect 78640 437452 78646 437464
rect 176470 437452 176476 437464
rect 176528 437492 176534 437504
rect 177574 437492 177580 437504
rect 176528 437464 177580 437492
rect 176528 437452 176534 437464
rect 177574 437452 177580 437464
rect 177632 437452 177638 437504
rect 183462 437452 183468 437504
rect 183520 437492 183526 437504
rect 184566 437492 184572 437504
rect 183520 437464 184572 437492
rect 183520 437452 183526 437464
rect 184566 437452 184572 437464
rect 184624 437452 184630 437504
rect 263778 437452 263784 437504
rect 263836 437492 263842 437504
rect 266630 437492 266636 437504
rect 263836 437464 266636 437492
rect 263836 437452 263842 437464
rect 266630 437452 266636 437464
rect 266688 437452 266694 437504
rect 76558 437384 76564 437436
rect 76616 437424 76622 437436
rect 82906 437424 82912 437436
rect 76616 437396 82912 437424
rect 76616 437384 76622 437396
rect 82906 437384 82912 437396
rect 82964 437384 82970 437436
rect 101398 437384 101404 437436
rect 101456 437424 101462 437436
rect 104158 437424 104164 437436
rect 101456 437396 104164 437424
rect 101456 437384 101462 437396
rect 104158 437384 104164 437396
rect 104216 437384 104222 437436
rect 102502 437316 102508 437368
rect 102560 437356 102566 437368
rect 105538 437356 105544 437368
rect 102560 437328 105544 437356
rect 102560 437316 102566 437328
rect 105538 437316 105544 437328
rect 105596 437316 105602 437368
rect 110782 436704 110788 436756
rect 110840 436744 110846 436756
rect 180058 436744 180064 436756
rect 110840 436716 180064 436744
rect 110840 436704 110846 436716
rect 180058 436704 180064 436716
rect 180116 436704 180122 436756
rect 95878 436296 95884 436348
rect 95936 436336 95942 436348
rect 96982 436336 96988 436348
rect 95936 436308 96988 436336
rect 95936 436296 95942 436308
rect 96982 436296 96988 436308
rect 97040 436296 97046 436348
rect 68922 436268 68928 436280
rect 64846 436240 68928 436268
rect 52270 436160 52276 436212
rect 52328 436200 52334 436212
rect 64846 436200 64874 436240
rect 68922 436228 68928 436240
rect 68980 436228 68986 436280
rect 70486 436200 70492 436212
rect 52328 436172 64874 436200
rect 68572 436172 70492 436200
rect 52328 436160 52334 436172
rect 41230 436092 41236 436144
rect 41288 436132 41294 436144
rect 68572 436132 68600 436172
rect 70486 436160 70492 436172
rect 70544 436160 70550 436212
rect 71774 436200 71780 436212
rect 71148 436172 71780 436200
rect 41288 436104 68600 436132
rect 41288 436092 41294 436104
rect 68646 436092 68652 436144
rect 68704 436132 68710 436144
rect 71148 436132 71176 436172
rect 71774 436160 71780 436172
rect 71832 436200 71838 436212
rect 72694 436200 72700 436212
rect 71832 436172 72700 436200
rect 71832 436160 71838 436172
rect 72694 436160 72700 436172
rect 72752 436160 72758 436212
rect 68704 436104 71176 436132
rect 68704 436092 68710 436104
rect 71682 436092 71688 436144
rect 71740 436132 71746 436144
rect 72418 436132 72424 436144
rect 71740 436104 72424 436132
rect 71740 436092 71746 436104
rect 72418 436092 72424 436104
rect 72476 436092 72482 436144
rect 96338 436092 96344 436144
rect 96396 436132 96402 436144
rect 100018 436132 100024 436144
rect 96396 436104 100024 436132
rect 96396 436092 96402 436104
rect 100018 436092 100024 436104
rect 100076 436092 100082 436144
rect 103882 436092 103888 436144
rect 103940 436132 103946 436144
rect 104158 436132 104164 436144
rect 103940 436104 104164 436132
rect 103940 436092 103946 436104
rect 104158 436092 104164 436104
rect 104216 436132 104222 436144
rect 116026 436132 116032 436144
rect 104216 436104 116032 436132
rect 104216 436092 104222 436104
rect 116026 436092 116032 436104
rect 116084 436132 116090 436144
rect 116578 436132 116584 436144
rect 116084 436104 116584 436132
rect 116084 436092 116090 436104
rect 116578 436092 116584 436104
rect 116636 436092 116642 436144
rect 188338 436092 188344 436144
rect 188396 436132 188402 436144
rect 191650 436132 191656 436144
rect 188396 436104 191656 436132
rect 188396 436092 188402 436104
rect 191650 436092 191656 436104
rect 191708 436092 191714 436144
rect 255498 436024 255504 436076
rect 255556 436064 255562 436076
rect 267918 436064 267924 436076
rect 255556 436036 267924 436064
rect 255556 436024 255562 436036
rect 267918 436024 267924 436036
rect 267976 436064 267982 436076
rect 276290 436064 276296 436076
rect 267976 436036 276296 436064
rect 267976 436024 267982 436036
rect 276290 436024 276296 436036
rect 276348 436024 276354 436076
rect 170398 435344 170404 435396
rect 170456 435384 170462 435396
rect 181530 435384 181536 435396
rect 170456 435356 181536 435384
rect 170456 435344 170462 435356
rect 181530 435344 181536 435356
rect 181588 435344 181594 435396
rect 264238 435344 264244 435396
rect 264296 435384 264302 435396
rect 274818 435384 274824 435396
rect 264296 435356 274824 435384
rect 264296 435344 264302 435356
rect 274818 435344 274824 435356
rect 274876 435344 274882 435396
rect 3418 434800 3424 434852
rect 3476 434840 3482 434852
rect 112254 434840 112260 434852
rect 3476 434812 112260 434840
rect 3476 434800 3482 434812
rect 112254 434800 112260 434812
rect 112312 434800 112318 434852
rect 62022 434732 62028 434784
rect 62080 434772 62086 434784
rect 191650 434772 191656 434784
rect 62080 434744 191656 434772
rect 62080 434732 62086 434744
rect 191650 434732 191656 434744
rect 191708 434732 191714 434784
rect 115750 434664 115756 434716
rect 115808 434704 115814 434716
rect 126238 434704 126244 434716
rect 115808 434676 126244 434704
rect 115808 434664 115814 434676
rect 126238 434664 126244 434676
rect 126296 434664 126302 434716
rect 68186 433984 68192 434036
rect 68244 434024 68250 434036
rect 191650 434024 191656 434036
rect 68244 433996 191656 434024
rect 68244 433984 68250 433996
rect 191650 433984 191656 433996
rect 191708 433984 191714 434036
rect 255498 433984 255504 434036
rect 255556 434024 255562 434036
rect 262858 434024 262864 434036
rect 255556 433996 262864 434024
rect 255556 433984 255562 433996
rect 262858 433984 262864 433996
rect 262916 433984 262922 434036
rect 67266 433780 67272 433832
rect 67324 433820 67330 433832
rect 71130 433820 71136 433832
rect 67324 433792 71136 433820
rect 67324 433780 67330 433792
rect 71130 433780 71136 433792
rect 71188 433780 71194 433832
rect 70670 433644 70676 433696
rect 70728 433644 70734 433696
rect 53742 433304 53748 433356
rect 53800 433344 53806 433356
rect 57698 433344 57704 433356
rect 53800 433316 57704 433344
rect 53800 433304 53806 433316
rect 57698 433304 57704 433316
rect 57756 433344 57762 433356
rect 66806 433344 66812 433356
rect 57756 433316 66812 433344
rect 57756 433304 57762 433316
rect 66806 433304 66812 433316
rect 66864 433304 66870 433356
rect 67726 433236 67732 433288
rect 67784 433276 67790 433288
rect 70688 433276 70716 433644
rect 276014 433344 276020 433356
rect 269040 433316 276020 433344
rect 269040 433288 269068 433316
rect 276014 433304 276020 433316
rect 276072 433304 276078 433356
rect 67784 433248 70716 433276
rect 67784 433236 67790 433248
rect 115842 433236 115848 433288
rect 115900 433276 115906 433288
rect 146938 433276 146944 433288
rect 115900 433248 146944 433276
rect 115900 433236 115906 433248
rect 146938 433236 146944 433248
rect 146996 433236 147002 433288
rect 155586 433236 155592 433288
rect 155644 433276 155650 433288
rect 155770 433276 155776 433288
rect 155644 433248 155776 433276
rect 155644 433236 155650 433248
rect 155770 433236 155776 433248
rect 155828 433236 155834 433288
rect 269022 433236 269028 433288
rect 269080 433236 269086 433288
rect 67542 433168 67548 433220
rect 67600 433208 67606 433220
rect 68278 433208 68284 433220
rect 67600 433180 68284 433208
rect 67600 433168 67606 433180
rect 68278 433168 68284 433180
rect 68336 433168 68342 433220
rect 155586 432556 155592 432608
rect 155644 432596 155650 432608
rect 191650 432596 191656 432608
rect 155644 432568 191656 432596
rect 155644 432556 155650 432568
rect 191650 432556 191656 432568
rect 191708 432556 191714 432608
rect 262858 432556 262864 432608
rect 262916 432596 262922 432608
rect 267918 432596 267924 432608
rect 262916 432568 267924 432596
rect 262916 432556 262922 432568
rect 267918 432556 267924 432568
rect 267976 432596 267982 432608
rect 269022 432596 269028 432608
rect 267976 432568 269028 432596
rect 267976 432556 267982 432568
rect 269022 432556 269028 432568
rect 269080 432556 269086 432608
rect 65702 432488 65708 432540
rect 65760 432528 65766 432540
rect 66162 432528 66168 432540
rect 65760 432500 66168 432528
rect 65760 432488 65766 432500
rect 66162 432488 66168 432500
rect 66220 432488 66226 432540
rect 63310 431944 63316 431996
rect 63368 431984 63374 431996
rect 178954 431984 178960 431996
rect 63368 431956 178960 431984
rect 63368 431944 63374 431956
rect 178954 431944 178960 431956
rect 179012 431944 179018 431996
rect 254210 431944 254216 431996
rect 254268 431984 254274 431996
rect 263778 431984 263784 431996
rect 254268 431956 263784 431984
rect 254268 431944 254274 431956
rect 263778 431944 263784 431956
rect 263836 431944 263842 431996
rect 56502 431196 56508 431248
rect 56560 431236 56566 431248
rect 67358 431236 67364 431248
rect 56560 431208 67364 431236
rect 56560 431196 56566 431208
rect 67358 431196 67364 431208
rect 67416 431196 67422 431248
rect 165430 431196 165436 431248
rect 165488 431236 165494 431248
rect 191742 431236 191748 431248
rect 165488 431208 191748 431236
rect 165488 431196 165494 431208
rect 191742 431196 191748 431208
rect 191800 431196 191806 431248
rect 255406 431196 255412 431248
rect 255464 431236 255470 431248
rect 262490 431236 262496 431248
rect 255464 431208 262496 431236
rect 255464 431196 255470 431208
rect 262490 431196 262496 431208
rect 262548 431196 262554 431248
rect 138658 430516 138664 430568
rect 138716 430556 138722 430568
rect 164970 430556 164976 430568
rect 138716 430528 164976 430556
rect 138716 430516 138722 430528
rect 164970 430516 164976 430528
rect 165028 430556 165034 430568
rect 165430 430556 165436 430568
rect 165028 430528 165436 430556
rect 165028 430516 165034 430528
rect 165430 430516 165436 430528
rect 165488 430516 165494 430568
rect 178954 430516 178960 430568
rect 179012 430556 179018 430568
rect 191006 430556 191012 430568
rect 179012 430528 191012 430556
rect 179012 430516 179018 430528
rect 191006 430516 191012 430528
rect 191064 430516 191070 430568
rect 114922 430448 114928 430500
rect 114980 430488 114986 430500
rect 141418 430488 141424 430500
rect 114980 430460 141424 430488
rect 114980 430448 114986 430460
rect 141418 430448 141424 430460
rect 141476 430448 141482 430500
rect 155770 429836 155776 429888
rect 155828 429876 155834 429888
rect 188338 429876 188344 429888
rect 155828 429848 188344 429876
rect 155828 429836 155834 429848
rect 188338 429836 188344 429848
rect 188396 429836 188402 429888
rect 255406 429496 255412 429548
rect 255464 429536 255470 429548
rect 259546 429536 259552 429548
rect 255464 429508 259552 429536
rect 255464 429496 255470 429508
rect 259546 429496 259552 429508
rect 259604 429496 259610 429548
rect 64690 429360 64696 429412
rect 64748 429400 64754 429412
rect 67266 429400 67272 429412
rect 64748 429372 67272 429400
rect 64748 429360 64754 429372
rect 67266 429360 67272 429372
rect 67324 429360 67330 429412
rect 48222 429156 48228 429208
rect 48280 429196 48286 429208
rect 66806 429196 66812 429208
rect 48280 429168 66812 429196
rect 48280 429156 48286 429168
rect 66806 429156 66812 429168
rect 66864 429156 66870 429208
rect 115842 429088 115848 429140
rect 115900 429128 115906 429140
rect 154022 429128 154028 429140
rect 115900 429100 154028 429128
rect 115900 429088 115906 429100
rect 154022 429088 154028 429100
rect 154080 429088 154086 429140
rect 154390 429088 154396 429140
rect 154448 429128 154454 429140
rect 190822 429128 190828 429140
rect 154448 429100 190828 429128
rect 154448 429088 154454 429100
rect 190822 429088 190828 429100
rect 190880 429088 190886 429140
rect 65794 427320 65800 427372
rect 65852 427360 65858 427372
rect 67542 427360 67548 427372
rect 65852 427332 67548 427360
rect 65852 427320 65858 427332
rect 67542 427320 67548 427332
rect 67600 427320 67606 427372
rect 122190 427048 122196 427100
rect 122248 427088 122254 427100
rect 133138 427088 133144 427100
rect 122248 427060 133144 427088
rect 122248 427048 122254 427060
rect 133138 427048 133144 427060
rect 133196 427048 133202 427100
rect 169018 427048 169024 427100
rect 169076 427088 169082 427100
rect 178034 427088 178040 427100
rect 169076 427060 178040 427088
rect 169076 427048 169082 427060
rect 178034 427048 178040 427060
rect 178092 427048 178098 427100
rect 284386 427048 284392 427100
rect 284444 427088 284450 427100
rect 291378 427088 291384 427100
rect 284444 427060 291384 427088
rect 284444 427048 284450 427060
rect 291378 427048 291384 427060
rect 291436 427088 291442 427100
rect 582558 427088 582564 427100
rect 291436 427060 582564 427088
rect 291436 427048 291442 427060
rect 582558 427048 582564 427060
rect 582616 427048 582622 427100
rect 115842 426436 115848 426488
rect 115900 426476 115906 426488
rect 125594 426476 125600 426488
rect 115900 426448 125600 426476
rect 115900 426436 115906 426448
rect 125594 426436 125600 426448
rect 125652 426436 125658 426488
rect 178034 426436 178040 426488
rect 178092 426476 178098 426488
rect 179322 426476 179328 426488
rect 178092 426448 179328 426476
rect 178092 426436 178098 426448
rect 179322 426436 179328 426448
rect 179380 426476 179386 426488
rect 191742 426476 191748 426488
rect 179380 426448 191748 426476
rect 179380 426436 179386 426448
rect 191742 426436 191748 426448
rect 191800 426436 191806 426488
rect 255406 426436 255412 426488
rect 255464 426476 255470 426488
rect 284386 426476 284392 426488
rect 255464 426448 284392 426476
rect 255464 426436 255470 426448
rect 284386 426436 284392 426448
rect 284444 426436 284450 426488
rect 67542 426368 67548 426420
rect 67600 426408 67606 426420
rect 68186 426408 68192 426420
rect 67600 426380 68192 426408
rect 67600 426368 67606 426380
rect 68186 426368 68192 426380
rect 68244 426368 68250 426420
rect 115750 426368 115756 426420
rect 115808 426408 115814 426420
rect 117498 426408 117504 426420
rect 115808 426380 117504 426408
rect 115808 426368 115814 426380
rect 117498 426368 117504 426380
rect 117556 426408 117562 426420
rect 119338 426408 119344 426420
rect 117556 426380 119344 426408
rect 117556 426368 117562 426380
rect 119338 426368 119344 426380
rect 119396 426368 119402 426420
rect 49602 425688 49608 425740
rect 49660 425728 49666 425740
rect 66990 425728 66996 425740
rect 49660 425700 66996 425728
rect 49660 425688 49666 425700
rect 66990 425688 66996 425700
rect 67048 425688 67054 425740
rect 256602 425688 256608 425740
rect 256660 425728 256666 425740
rect 273530 425728 273536 425740
rect 256660 425700 273536 425728
rect 256660 425688 256666 425700
rect 273530 425688 273536 425700
rect 273588 425688 273594 425740
rect 165614 425076 165620 425128
rect 165672 425116 165678 425128
rect 191742 425116 191748 425128
rect 165672 425088 191748 425116
rect 165672 425076 165678 425088
rect 191742 425076 191748 425088
rect 191800 425076 191806 425128
rect 115842 425008 115848 425060
rect 115900 425048 115906 425060
rect 130378 425048 130384 425060
rect 115900 425020 130384 425048
rect 115900 425008 115906 425020
rect 130378 425008 130384 425020
rect 130436 425008 130442 425060
rect 151722 425008 151728 425060
rect 151780 425048 151786 425060
rect 165632 425048 165660 425076
rect 151780 425020 165660 425048
rect 151780 425008 151786 425020
rect 182082 425008 182088 425060
rect 182140 425048 182146 425060
rect 191006 425048 191012 425060
rect 182140 425020 191012 425048
rect 182140 425008 182146 425020
rect 191006 425008 191012 425020
rect 191064 425008 191070 425060
rect 115106 424940 115112 424992
rect 115164 424980 115170 424992
rect 117314 424980 117320 424992
rect 115164 424952 117320 424980
rect 115164 424940 115170 424952
rect 117314 424940 117320 424952
rect 117372 424940 117378 424992
rect 169386 424464 169392 424516
rect 169444 424504 169450 424516
rect 182082 424504 182088 424516
rect 169444 424476 182088 424504
rect 169444 424464 169450 424476
rect 182082 424464 182088 424476
rect 182140 424464 182146 424516
rect 169570 424328 169576 424380
rect 169628 424368 169634 424380
rect 182818 424368 182824 424380
rect 169628 424340 182824 424368
rect 169628 424328 169634 424340
rect 182818 424328 182824 424340
rect 182876 424328 182882 424380
rect 256602 424328 256608 424380
rect 256660 424368 256666 424380
rect 274818 424368 274824 424380
rect 256660 424340 274824 424368
rect 256660 424328 256666 424340
rect 274818 424328 274824 424340
rect 274876 424328 274882 424380
rect 59262 423648 59268 423700
rect 59320 423688 59326 423700
rect 66714 423688 66720 423700
rect 59320 423660 66720 423688
rect 59320 423648 59326 423660
rect 66714 423648 66720 423660
rect 66772 423648 66778 423700
rect 60734 423580 60740 423632
rect 60792 423620 60798 423632
rect 62022 423620 62028 423632
rect 60792 423592 62028 423620
rect 60792 423580 60798 423592
rect 62022 423580 62028 423592
rect 62080 423620 62086 423632
rect 66806 423620 66812 423632
rect 62080 423592 66812 423620
rect 62080 423580 62086 423592
rect 66806 423580 66812 423592
rect 66864 423580 66870 423632
rect 115842 423580 115848 423632
rect 115900 423620 115906 423632
rect 170398 423620 170404 423632
rect 115900 423592 170404 423620
rect 115900 423580 115906 423592
rect 170398 423580 170404 423592
rect 170456 423580 170462 423632
rect 146110 423512 146116 423564
rect 146168 423552 146174 423564
rect 151078 423552 151084 423564
rect 146168 423524 151084 423552
rect 146168 423512 146174 423524
rect 151078 423512 151084 423524
rect 151136 423512 151142 423564
rect 253566 423376 253572 423428
rect 253624 423416 253630 423428
rect 256970 423416 256976 423428
rect 253624 423388 256976 423416
rect 253624 423376 253630 423388
rect 256970 423376 256976 423388
rect 257028 423376 257034 423428
rect 44082 422900 44088 422952
rect 44140 422940 44146 422952
rect 60734 422940 60740 422952
rect 44140 422912 60740 422940
rect 44140 422900 44146 422912
rect 60734 422900 60740 422912
rect 60792 422900 60798 422952
rect 151078 422288 151084 422340
rect 151136 422328 151142 422340
rect 191742 422328 191748 422340
rect 151136 422300 191748 422328
rect 151136 422288 151142 422300
rect 191742 422288 191748 422300
rect 191800 422288 191806 422340
rect 255498 422288 255504 422340
rect 255556 422328 255562 422340
rect 277762 422328 277768 422340
rect 255556 422300 277768 422328
rect 255556 422288 255562 422300
rect 277762 422288 277768 422300
rect 277820 422288 277826 422340
rect 152918 421540 152924 421592
rect 152976 421580 152982 421592
rect 177390 421580 177396 421592
rect 152976 421552 177396 421580
rect 152976 421540 152982 421552
rect 177390 421540 177396 421552
rect 177448 421540 177454 421592
rect 65978 420996 65984 421048
rect 66036 421036 66042 421048
rect 67542 421036 67548 421048
rect 66036 421008 67548 421036
rect 66036 420996 66042 421008
rect 67542 420996 67548 421008
rect 67600 420996 67606 421048
rect 50982 420928 50988 420980
rect 51040 420968 51046 420980
rect 66806 420968 66812 420980
rect 51040 420940 66812 420968
rect 51040 420928 51046 420940
rect 66806 420928 66812 420940
rect 66864 420928 66870 420980
rect 146110 420928 146116 420980
rect 146168 420968 146174 420980
rect 152550 420968 152556 420980
rect 146168 420940 152556 420968
rect 146168 420928 146174 420940
rect 152550 420928 152556 420940
rect 152608 420968 152614 420980
rect 153102 420968 153108 420980
rect 152608 420940 153108 420968
rect 152608 420928 152614 420940
rect 153102 420928 153108 420940
rect 153160 420928 153166 420980
rect 255498 420928 255504 420980
rect 255556 420968 255562 420980
rect 298278 420968 298284 420980
rect 255556 420940 298284 420968
rect 255556 420928 255562 420940
rect 298278 420928 298284 420940
rect 298336 420928 298342 420980
rect 61838 420860 61844 420912
rect 61896 420900 61902 420912
rect 66898 420900 66904 420912
rect 61896 420872 66904 420900
rect 61896 420860 61902 420872
rect 66898 420860 66904 420872
rect 66956 420860 66962 420912
rect 57882 420180 57888 420232
rect 57940 420220 57946 420232
rect 66806 420220 66812 420232
rect 57940 420192 66812 420220
rect 57940 420180 57946 420192
rect 66806 420180 66812 420192
rect 66864 420180 66870 420232
rect 186958 420180 186964 420232
rect 187016 420220 187022 420232
rect 192478 420220 192484 420232
rect 187016 420192 192484 420220
rect 187016 420180 187022 420192
rect 192478 420180 192484 420192
rect 192536 420180 192542 420232
rect 174630 419500 174636 419552
rect 174688 419540 174694 419552
rect 192386 419540 192392 419552
rect 174688 419512 192392 419540
rect 174688 419500 174694 419512
rect 192386 419500 192392 419512
rect 192444 419500 192450 419552
rect 255498 419500 255504 419552
rect 255556 419540 255562 419552
rect 280430 419540 280436 419552
rect 255556 419512 280436 419540
rect 255556 419500 255562 419512
rect 280430 419500 280436 419512
rect 280488 419540 280494 419552
rect 285858 419540 285864 419552
rect 280488 419512 285864 419540
rect 280488 419500 280494 419512
rect 285858 419500 285864 419512
rect 285916 419500 285922 419552
rect 115842 419432 115848 419484
rect 115900 419472 115906 419484
rect 142798 419472 142804 419484
rect 115900 419444 142804 419472
rect 115900 419432 115906 419444
rect 142798 419432 142804 419444
rect 142856 419432 142862 419484
rect 255406 419432 255412 419484
rect 255464 419472 255470 419484
rect 281534 419472 281540 419484
rect 255464 419444 281540 419472
rect 255464 419432 255470 419444
rect 281534 419432 281540 419444
rect 281592 419432 281598 419484
rect 122098 419364 122104 419416
rect 122156 419404 122162 419416
rect 123018 419404 123024 419416
rect 122156 419376 123024 419404
rect 122156 419364 122162 419376
rect 123018 419364 123024 419376
rect 123076 419364 123082 419416
rect 281534 418752 281540 418804
rect 281592 418792 281598 418804
rect 285858 418792 285864 418804
rect 281592 418764 285864 418792
rect 281592 418752 281598 418764
rect 285858 418752 285864 418764
rect 285916 418792 285922 418804
rect 582374 418792 582380 418804
rect 285916 418764 582380 418792
rect 285916 418752 285922 418764
rect 582374 418752 582380 418764
rect 582432 418752 582438 418804
rect 63218 418276 63224 418328
rect 63276 418316 63282 418328
rect 66438 418316 66444 418328
rect 63276 418288 66444 418316
rect 63276 418276 63282 418288
rect 66438 418276 66444 418288
rect 66496 418276 66502 418328
rect 63402 418072 63408 418124
rect 63460 418112 63466 418124
rect 66438 418112 66444 418124
rect 63460 418084 66444 418112
rect 63460 418072 63466 418084
rect 66438 418072 66444 418084
rect 66496 418072 66502 418124
rect 153102 417392 153108 417444
rect 153160 417432 153166 417444
rect 155678 417432 155684 417444
rect 153160 417404 155684 417432
rect 153160 417392 153166 417404
rect 155678 417392 155684 417404
rect 155736 417432 155742 417444
rect 179414 417432 179420 417444
rect 155736 417404 179420 417432
rect 155736 417392 155742 417404
rect 179414 417392 179420 417404
rect 179472 417392 179478 417444
rect 283650 417392 283656 417444
rect 283708 417432 283714 417444
rect 582650 417432 582656 417444
rect 283708 417404 582656 417432
rect 283708 417392 283714 417404
rect 582650 417392 582656 417404
rect 582708 417392 582714 417444
rect 117406 417188 117412 417240
rect 117464 417228 117470 417240
rect 122190 417228 122196 417240
rect 117464 417200 122196 417228
rect 117464 417188 117470 417200
rect 122190 417188 122196 417200
rect 122248 417188 122254 417240
rect 126238 417188 126244 417240
rect 126296 417228 126302 417240
rect 126882 417228 126888 417240
rect 126296 417200 126888 417228
rect 126296 417188 126302 417200
rect 126882 417188 126888 417200
rect 126940 417188 126946 417240
rect 57790 416780 57796 416832
rect 57848 416820 57854 416832
rect 57848 416792 61884 416820
rect 57848 416780 57854 416792
rect 61856 416764 61884 416792
rect 115842 416780 115848 416832
rect 115900 416820 115906 416832
rect 117406 416820 117412 416832
rect 115900 416792 117412 416820
rect 115900 416780 115906 416792
rect 117406 416780 117412 416792
rect 117464 416780 117470 416832
rect 126882 416780 126888 416832
rect 126940 416820 126946 416832
rect 148318 416820 148324 416832
rect 126940 416792 148324 416820
rect 126940 416780 126946 416792
rect 148318 416780 148324 416792
rect 148376 416780 148382 416832
rect 177298 416780 177304 416832
rect 177356 416820 177362 416832
rect 191742 416820 191748 416832
rect 177356 416792 191748 416820
rect 177356 416780 177362 416792
rect 191742 416780 191748 416792
rect 191800 416780 191806 416832
rect 255498 416780 255504 416832
rect 255556 416820 255562 416832
rect 283190 416820 283196 416832
rect 255556 416792 283196 416820
rect 255556 416780 255562 416792
rect 283190 416780 283196 416792
rect 283248 416820 283254 416832
rect 283650 416820 283656 416832
rect 283248 416792 283656 416820
rect 283248 416780 283254 416792
rect 283650 416780 283656 416792
rect 283708 416780 283714 416832
rect 61838 416712 61844 416764
rect 61896 416712 61902 416764
rect 179414 416712 179420 416764
rect 179472 416752 179478 416764
rect 191650 416752 191656 416764
rect 179472 416724 191656 416752
rect 179472 416712 179478 416724
rect 191650 416712 191656 416724
rect 191708 416712 191714 416764
rect 255406 416712 255412 416764
rect 255464 416752 255470 416764
rect 278958 416752 278964 416764
rect 255464 416724 278964 416752
rect 255464 416712 255470 416724
rect 278958 416712 278964 416724
rect 279016 416752 279022 416764
rect 279326 416752 279332 416764
rect 279016 416724 279332 416752
rect 279016 416712 279022 416724
rect 279326 416712 279332 416724
rect 279384 416712 279390 416764
rect 122098 416032 122104 416084
rect 122156 416072 122162 416084
rect 189718 416072 189724 416084
rect 122156 416044 189724 416072
rect 122156 416032 122162 416044
rect 189718 416032 189724 416044
rect 189776 416032 189782 416084
rect 115842 415624 115848 415676
rect 115900 415664 115906 415676
rect 120074 415664 120080 415676
rect 115900 415636 120080 415664
rect 115900 415624 115906 415636
rect 120074 415624 120080 415636
rect 120132 415624 120138 415676
rect 61838 415420 61844 415472
rect 61896 415460 61902 415472
rect 66898 415460 66904 415472
rect 61896 415432 66904 415460
rect 61896 415420 61902 415432
rect 66898 415420 66904 415432
rect 66956 415420 66962 415472
rect 114922 414672 114928 414724
rect 114980 414712 114986 414724
rect 124858 414712 124864 414724
rect 114980 414684 124864 414712
rect 114980 414672 114986 414684
rect 124858 414672 124864 414684
rect 124916 414672 124922 414724
rect 176562 414672 176568 414724
rect 176620 414712 176626 414724
rect 189718 414712 189724 414724
rect 176620 414684 189724 414712
rect 176620 414672 176626 414684
rect 189718 414672 189724 414684
rect 189776 414672 189782 414724
rect 54846 413992 54852 414044
rect 54904 414032 54910 414044
rect 66806 414032 66812 414044
rect 54904 414004 66812 414032
rect 54904 413992 54910 414004
rect 66806 413992 66812 414004
rect 66864 413992 66870 414044
rect 154022 413992 154028 414044
rect 154080 414032 154086 414044
rect 191190 414032 191196 414044
rect 154080 414004 191196 414032
rect 154080 413992 154086 414004
rect 191190 413992 191196 414004
rect 191248 413992 191254 414044
rect 57974 413244 57980 413296
rect 58032 413284 58038 413296
rect 66622 413284 66628 413296
rect 58032 413256 66628 413284
rect 58032 413244 58038 413256
rect 66622 413244 66628 413256
rect 66680 413244 66686 413296
rect 123018 412700 123024 412752
rect 123076 412740 123082 412752
rect 142798 412740 142804 412752
rect 123076 412712 142804 412740
rect 123076 412700 123082 412712
rect 142798 412700 142804 412712
rect 142856 412700 142862 412752
rect 115842 412632 115848 412684
rect 115900 412672 115906 412684
rect 147030 412672 147036 412684
rect 115900 412644 147036 412672
rect 115900 412632 115906 412644
rect 147030 412632 147036 412644
rect 147088 412632 147094 412684
rect 115750 412564 115756 412616
rect 115808 412604 115814 412616
rect 123018 412604 123024 412616
rect 115808 412576 123024 412604
rect 115808 412564 115814 412576
rect 123018 412564 123024 412576
rect 123076 412564 123082 412616
rect 255498 412564 255504 412616
rect 255556 412604 255562 412616
rect 281810 412604 281816 412616
rect 255556 412576 281816 412604
rect 255556 412564 255562 412576
rect 281810 412564 281816 412576
rect 281868 412564 281874 412616
rect 52178 411884 52184 411936
rect 52236 411924 52242 411936
rect 55030 411924 55036 411936
rect 52236 411896 55036 411924
rect 52236 411884 52242 411896
rect 55030 411884 55036 411896
rect 55088 411924 55094 411936
rect 57974 411924 57980 411936
rect 55088 411896 57980 411924
rect 55088 411884 55094 411896
rect 57974 411884 57980 411896
rect 58032 411884 58038 411936
rect 165430 411884 165436 411936
rect 165488 411924 165494 411936
rect 191742 411924 191748 411936
rect 165488 411896 191748 411924
rect 165488 411884 165494 411896
rect 191742 411884 191748 411896
rect 191800 411884 191806 411936
rect 64782 411272 64788 411324
rect 64840 411312 64846 411324
rect 66898 411312 66904 411324
rect 64840 411284 66904 411312
rect 64840 411272 64846 411284
rect 66898 411272 66904 411284
rect 66956 411272 66962 411324
rect 115842 411204 115848 411256
rect 115900 411244 115906 411256
rect 126238 411244 126244 411256
rect 115900 411216 126244 411244
rect 115900 411204 115906 411216
rect 126238 411204 126244 411216
rect 126296 411204 126302 411256
rect 59998 410524 60004 410576
rect 60056 410564 60062 410576
rect 66806 410564 66812 410576
rect 60056 410536 66812 410564
rect 60056 410524 60062 410536
rect 66806 410524 66812 410536
rect 66864 410524 66870 410576
rect 154390 410524 154396 410576
rect 154448 410564 154454 410576
rect 161474 410564 161480 410576
rect 154448 410536 161480 410564
rect 154448 410524 154454 410536
rect 161474 410524 161480 410536
rect 161532 410524 161538 410576
rect 183186 410524 183192 410576
rect 183244 410564 183250 410576
rect 191742 410564 191748 410576
rect 183244 410536 191748 410564
rect 183244 410524 183250 410536
rect 191742 410524 191748 410536
rect 191800 410524 191806 410576
rect 115934 409844 115940 409896
rect 115992 409884 115998 409896
rect 154390 409884 154396 409896
rect 115992 409856 154396 409884
rect 115992 409844 115998 409856
rect 154390 409844 154396 409856
rect 154448 409844 154454 409896
rect 135990 409776 135996 409828
rect 136048 409816 136054 409828
rect 141878 409816 141884 409828
rect 136048 409788 141884 409816
rect 136048 409776 136054 409788
rect 141878 409776 141884 409788
rect 141936 409816 141942 409828
rect 177298 409816 177304 409828
rect 141936 409788 177304 409816
rect 141936 409776 141942 409788
rect 177298 409776 177304 409788
rect 177356 409776 177362 409828
rect 115842 409708 115848 409760
rect 115900 409748 115906 409760
rect 122098 409748 122104 409760
rect 115900 409720 122104 409748
rect 115900 409708 115906 409720
rect 122098 409708 122104 409720
rect 122156 409708 122162 409760
rect 39850 409096 39856 409148
rect 39908 409136 39914 409148
rect 52362 409136 52368 409148
rect 39908 409108 52368 409136
rect 39908 409096 39914 409108
rect 52362 409096 52368 409108
rect 52420 409136 52426 409148
rect 59998 409136 60004 409148
rect 52420 409108 60004 409136
rect 52420 409096 52426 409108
rect 59998 409096 60004 409108
rect 60056 409096 60062 409148
rect 128998 409096 129004 409148
rect 129056 409136 129062 409148
rect 135990 409136 135996 409148
rect 129056 409108 135996 409136
rect 129056 409096 129062 409108
rect 135990 409096 135996 409108
rect 136048 409096 136054 409148
rect 153838 409096 153844 409148
rect 153896 409136 153902 409148
rect 184290 409136 184296 409148
rect 153896 409108 184296 409136
rect 153896 409096 153902 409108
rect 184290 409096 184296 409108
rect 184348 409096 184354 409148
rect 271782 409096 271788 409148
rect 271840 409136 271846 409148
rect 280154 409136 280160 409148
rect 271840 409108 280160 409136
rect 271840 409096 271846 409108
rect 280154 409096 280160 409108
rect 280212 409096 280218 409148
rect 63310 408484 63316 408536
rect 63368 408524 63374 408536
rect 66438 408524 66444 408536
rect 63368 408496 66444 408524
rect 63368 408484 63374 408496
rect 66438 408484 66444 408496
rect 66496 408484 66502 408536
rect 115842 408484 115848 408536
rect 115900 408524 115906 408536
rect 141418 408524 141424 408536
rect 115900 408496 141424 408524
rect 115900 408484 115906 408496
rect 141418 408484 141424 408496
rect 141476 408484 141482 408536
rect 255406 408484 255412 408536
rect 255464 408524 255470 408536
rect 270770 408524 270776 408536
rect 255464 408496 270776 408524
rect 255464 408484 255470 408496
rect 270770 408484 270776 408496
rect 270828 408524 270834 408536
rect 271782 408524 271788 408536
rect 270828 408496 271788 408524
rect 270828 408484 270834 408496
rect 271782 408484 271788 408496
rect 271840 408484 271846 408536
rect 255406 407804 255412 407856
rect 255464 407844 255470 407856
rect 262398 407844 262404 407856
rect 255464 407816 262404 407844
rect 255464 407804 255470 407816
rect 262398 407804 262404 407816
rect 262456 407804 262462 407856
rect 48130 407736 48136 407788
rect 48188 407776 48194 407788
rect 66806 407776 66812 407788
rect 48188 407748 66812 407776
rect 48188 407736 48194 407748
rect 66806 407736 66812 407748
rect 66864 407736 66870 407788
rect 186130 407736 186136 407788
rect 186188 407776 186194 407788
rect 193306 407776 193312 407788
rect 186188 407748 193312 407776
rect 186188 407736 186194 407748
rect 193306 407736 193312 407748
rect 193364 407736 193370 407788
rect 255498 407736 255504 407788
rect 255556 407776 255562 407788
rect 267826 407776 267832 407788
rect 255556 407748 267832 407776
rect 255556 407736 255562 407748
rect 267826 407736 267832 407748
rect 267884 407736 267890 407788
rect 124858 407124 124864 407176
rect 124916 407164 124922 407176
rect 185578 407164 185584 407176
rect 124916 407136 185584 407164
rect 124916 407124 124922 407136
rect 185578 407124 185584 407136
rect 185636 407124 185642 407176
rect 113082 407056 113088 407108
rect 113140 407096 113146 407108
rect 135898 407096 135904 407108
rect 113140 407068 135904 407096
rect 113140 407056 113146 407068
rect 135898 407056 135904 407068
rect 135956 407056 135962 407108
rect 50890 406376 50896 406428
rect 50948 406416 50954 406428
rect 64598 406416 64604 406428
rect 50948 406388 64604 406416
rect 50948 406376 50954 406388
rect 64598 406376 64604 406388
rect 64656 406416 64662 406428
rect 66438 406416 66444 406428
rect 64656 406388 66444 406416
rect 64656 406376 64662 406388
rect 66438 406376 66444 406388
rect 66496 406376 66502 406428
rect 119338 406376 119344 406428
rect 119396 406416 119402 406428
rect 143258 406416 143264 406428
rect 119396 406388 143264 406416
rect 119396 406376 119402 406388
rect 143258 406376 143264 406388
rect 143316 406416 143322 406428
rect 177390 406416 177396 406428
rect 143316 406388 177396 406416
rect 143316 406376 143322 406388
rect 177390 406376 177396 406388
rect 177448 406376 177454 406428
rect 186130 405968 186136 406020
rect 186188 406008 186194 406020
rect 187050 406008 187056 406020
rect 186188 405980 187056 406008
rect 186188 405968 186194 405980
rect 187050 405968 187056 405980
rect 187108 405968 187114 406020
rect 191006 405736 191012 405748
rect 161446 405708 191012 405736
rect 161446 405680 161474 405708
rect 191006 405696 191012 405708
rect 191064 405696 191070 405748
rect 255498 405696 255504 405748
rect 255556 405736 255562 405748
rect 281810 405736 281816 405748
rect 255556 405708 281816 405736
rect 255556 405696 255562 405708
rect 281810 405696 281816 405708
rect 281868 405696 281874 405748
rect 153010 405628 153016 405680
rect 153068 405668 153074 405680
rect 161446 405668 161480 405680
rect 153068 405640 161480 405668
rect 153068 405628 153074 405640
rect 161474 405628 161480 405640
rect 161532 405628 161538 405680
rect 181622 405628 181628 405680
rect 181680 405668 181686 405680
rect 181990 405668 181996 405680
rect 181680 405640 181996 405668
rect 181680 405628 181686 405640
rect 181990 405628 181996 405640
rect 182048 405668 182054 405680
rect 191742 405668 191748 405680
rect 182048 405640 191748 405668
rect 182048 405628 182054 405640
rect 191742 405628 191748 405640
rect 191800 405628 191806 405680
rect 62022 404336 62028 404388
rect 62080 404376 62086 404388
rect 66898 404376 66904 404388
rect 62080 404348 66904 404376
rect 62080 404336 62086 404348
rect 66898 404336 66904 404348
rect 66956 404336 66962 404388
rect 115842 404336 115848 404388
rect 115900 404376 115906 404388
rect 146938 404376 146944 404388
rect 115900 404348 146944 404376
rect 115900 404336 115906 404348
rect 146938 404336 146944 404348
rect 146996 404336 147002 404388
rect 178862 404336 178868 404388
rect 178920 404376 178926 404388
rect 181622 404376 181628 404388
rect 178920 404348 181628 404376
rect 178920 404336 178926 404348
rect 181622 404336 181628 404348
rect 181680 404336 181686 404388
rect 154298 404268 154304 404320
rect 154356 404308 154362 404320
rect 158714 404308 158720 404320
rect 154356 404280 158720 404308
rect 154356 404268 154362 404280
rect 158714 404268 158720 404280
rect 158772 404268 158778 404320
rect 162762 404268 162768 404320
rect 162820 404308 162826 404320
rect 191742 404308 191748 404320
rect 162820 404280 191748 404308
rect 162820 404268 162826 404280
rect 191742 404268 191748 404280
rect 191800 404268 191806 404320
rect 262858 403588 262864 403640
rect 262916 403628 262922 403640
rect 270494 403628 270500 403640
rect 262916 403600 270500 403628
rect 262916 403588 262922 403600
rect 270494 403588 270500 403600
rect 270552 403588 270558 403640
rect 119982 403044 119988 403096
rect 120040 403084 120046 403096
rect 154298 403084 154304 403096
rect 120040 403056 154304 403084
rect 120040 403044 120046 403056
rect 154298 403044 154304 403056
rect 154356 403044 154362 403096
rect 54754 402976 54760 403028
rect 54812 403016 54818 403028
rect 66438 403016 66444 403028
rect 54812 402988 66444 403016
rect 54812 402976 54818 402988
rect 66438 402976 66444 402988
rect 66496 402976 66502 403028
rect 115842 402976 115848 403028
rect 115900 403016 115906 403028
rect 151170 403016 151176 403028
rect 115900 402988 151176 403016
rect 115900 402976 115906 402988
rect 151170 402976 151176 402988
rect 151228 402976 151234 403028
rect 157978 402976 157984 403028
rect 158036 403016 158042 403028
rect 162762 403016 162768 403028
rect 158036 402988 162768 403016
rect 158036 402976 158042 402988
rect 162762 402976 162768 402988
rect 162820 402976 162826 403028
rect 255406 402976 255412 403028
rect 255464 403016 255470 403028
rect 291378 403016 291384 403028
rect 255464 402988 291384 403016
rect 255464 402976 255470 402988
rect 291378 402976 291384 402988
rect 291436 402976 291442 403028
rect 55122 402908 55128 402960
rect 55180 402948 55186 402960
rect 67634 402948 67640 402960
rect 55180 402920 67640 402948
rect 55180 402908 55186 402920
rect 67634 402908 67640 402920
rect 67692 402908 67698 402960
rect 161382 402296 161388 402348
rect 161440 402336 161446 402348
rect 176654 402336 176660 402348
rect 161440 402308 176660 402336
rect 161440 402296 161446 402308
rect 176654 402296 176660 402308
rect 176712 402296 176718 402348
rect 115934 402228 115940 402280
rect 115992 402268 115998 402280
rect 184750 402268 184756 402280
rect 115992 402240 184756 402268
rect 115992 402228 115998 402240
rect 184750 402228 184756 402240
rect 184808 402228 184814 402280
rect 184750 401684 184756 401736
rect 184808 401724 184814 401736
rect 186958 401724 186964 401736
rect 184808 401696 186964 401724
rect 184808 401684 184814 401696
rect 186958 401684 186964 401696
rect 187016 401684 187022 401736
rect 176654 401616 176660 401668
rect 176712 401656 176718 401668
rect 177942 401656 177948 401668
rect 176712 401628 177948 401656
rect 176712 401616 176718 401628
rect 177942 401616 177948 401628
rect 178000 401656 178006 401668
rect 191006 401656 191012 401668
rect 178000 401628 191012 401656
rect 178000 401616 178006 401628
rect 191006 401616 191012 401628
rect 191064 401616 191070 401668
rect 255406 401616 255412 401668
rect 255464 401656 255470 401668
rect 259546 401656 259552 401668
rect 255464 401628 259552 401656
rect 255464 401616 255470 401628
rect 259546 401616 259552 401628
rect 259604 401616 259610 401668
rect 169018 401548 169024 401600
rect 169076 401588 169082 401600
rect 173526 401588 173532 401600
rect 169076 401560 173532 401588
rect 169076 401548 169082 401560
rect 173526 401548 173532 401560
rect 173584 401588 173590 401600
rect 191742 401588 191748 401600
rect 173584 401560 191748 401588
rect 173584 401548 173590 401560
rect 191742 401548 191748 401560
rect 191800 401548 191806 401600
rect 114830 400936 114836 400988
rect 114888 400976 114894 400988
rect 119982 400976 119988 400988
rect 114888 400948 119988 400976
rect 114888 400936 114894 400948
rect 119982 400936 119988 400948
rect 120040 400936 120046 400988
rect 118786 400868 118792 400920
rect 118844 400908 118850 400920
rect 143534 400908 143540 400920
rect 118844 400880 143540 400908
rect 118844 400868 118850 400880
rect 143534 400868 143540 400880
rect 143592 400868 143598 400920
rect 177850 400596 177856 400648
rect 177908 400636 177914 400648
rect 178770 400636 178776 400648
rect 177908 400608 178776 400636
rect 177908 400596 177914 400608
rect 178770 400596 178776 400608
rect 178828 400596 178834 400648
rect 58986 400188 58992 400240
rect 59044 400228 59050 400240
rect 66438 400228 66444 400240
rect 59044 400200 66444 400228
rect 59044 400188 59050 400200
rect 66438 400188 66444 400200
rect 66496 400188 66502 400240
rect 115382 400188 115388 400240
rect 115440 400228 115446 400240
rect 122098 400228 122104 400240
rect 115440 400200 122104 400228
rect 115440 400188 115446 400200
rect 122098 400188 122104 400200
rect 122156 400188 122162 400240
rect 128998 400188 129004 400240
rect 129056 400228 129062 400240
rect 177850 400228 177856 400240
rect 129056 400200 177856 400228
rect 129056 400188 129062 400200
rect 177850 400188 177856 400200
rect 177908 400188 177914 400240
rect 255406 400188 255412 400240
rect 255464 400228 255470 400240
rect 280338 400228 280344 400240
rect 255464 400200 280344 400228
rect 255464 400188 255470 400200
rect 280338 400188 280344 400200
rect 280396 400188 280402 400240
rect 147030 399440 147036 399492
rect 147088 399480 147094 399492
rect 180242 399480 180248 399492
rect 147088 399452 180248 399480
rect 147088 399440 147094 399452
rect 180242 399440 180248 399452
rect 180300 399440 180306 399492
rect 53650 398828 53656 398880
rect 53708 398868 53714 398880
rect 66806 398868 66812 398880
rect 53708 398840 66812 398868
rect 53708 398828 53714 398840
rect 66806 398828 66812 398840
rect 66864 398828 66870 398880
rect 188338 398828 188344 398880
rect 188396 398868 188402 398880
rect 191006 398868 191012 398880
rect 188396 398840 191012 398868
rect 188396 398828 188402 398840
rect 191006 398828 191012 398840
rect 191064 398828 191070 398880
rect 61930 398760 61936 398812
rect 61988 398800 61994 398812
rect 67082 398800 67088 398812
rect 61988 398772 67088 398800
rect 61988 398760 61994 398772
rect 67082 398760 67088 398772
rect 67140 398760 67146 398812
rect 276474 398760 276480 398812
rect 276532 398800 276538 398812
rect 277486 398800 277492 398812
rect 276532 398772 277492 398800
rect 276532 398760 276538 398772
rect 277486 398760 277492 398772
rect 277544 398760 277550 398812
rect 115842 398284 115848 398336
rect 115900 398324 115906 398336
rect 116118 398324 116124 398336
rect 115900 398296 116124 398324
rect 115900 398284 115906 398296
rect 116118 398284 116124 398296
rect 116176 398324 116182 398336
rect 118786 398324 118792 398336
rect 116176 398296 118792 398324
rect 116176 398284 116182 398296
rect 118786 398284 118792 398296
rect 118844 398284 118850 398336
rect 253566 398148 253572 398200
rect 253624 398188 253630 398200
rect 262490 398188 262496 398200
rect 253624 398160 262496 398188
rect 253624 398148 253630 398160
rect 262490 398148 262496 398160
rect 262548 398148 262554 398200
rect 118786 398080 118792 398132
rect 118844 398120 118850 398132
rect 149054 398120 149060 398132
rect 118844 398092 149060 398120
rect 118844 398080 118850 398092
rect 149054 398080 149060 398092
rect 149112 398080 149118 398132
rect 255406 398080 255412 398132
rect 255464 398120 255470 398132
rect 276014 398120 276020 398132
rect 255464 398092 276020 398120
rect 255464 398080 255470 398092
rect 276014 398080 276020 398092
rect 276072 398120 276078 398132
rect 276474 398120 276480 398132
rect 276072 398092 276480 398120
rect 276072 398080 276078 398092
rect 276474 398080 276480 398092
rect 276532 398080 276538 398132
rect 168098 397536 168104 397588
rect 168156 397576 168162 397588
rect 169754 397576 169760 397588
rect 168156 397548 169760 397576
rect 168156 397536 168162 397548
rect 169754 397536 169760 397548
rect 169812 397576 169818 397588
rect 190822 397576 190828 397588
rect 169812 397548 190828 397576
rect 169812 397536 169818 397548
rect 190822 397536 190828 397548
rect 190880 397536 190886 397588
rect 4798 397468 4804 397520
rect 4856 397508 4862 397520
rect 64598 397508 64604 397520
rect 4856 397480 64604 397508
rect 4856 397468 4862 397480
rect 64598 397468 64604 397480
rect 64656 397508 64662 397520
rect 66806 397508 66812 397520
rect 64656 397480 66812 397508
rect 64656 397468 64662 397480
rect 66806 397468 66812 397480
rect 66864 397468 66870 397520
rect 126238 397468 126244 397520
rect 126296 397508 126302 397520
rect 178678 397508 178684 397520
rect 126296 397480 178684 397508
rect 126296 397468 126302 397480
rect 178678 397468 178684 397480
rect 178736 397468 178742 397520
rect 162118 397264 162124 397316
rect 162176 397304 162182 397316
rect 162670 397304 162676 397316
rect 162176 397276 162676 397304
rect 162176 397264 162182 397276
rect 162670 397264 162676 397276
rect 162728 397264 162734 397316
rect 115750 397060 115756 397112
rect 115808 397100 115814 397112
rect 118786 397100 118792 397112
rect 115808 397072 118792 397100
rect 115808 397060 115814 397072
rect 118786 397060 118792 397072
rect 118844 397060 118850 397112
rect 41322 396720 41328 396772
rect 41380 396760 41386 396772
rect 60734 396760 60740 396772
rect 41380 396732 60740 396760
rect 41380 396720 41386 396732
rect 60734 396720 60740 396732
rect 60792 396720 60798 396772
rect 130378 396720 130384 396772
rect 130436 396760 130442 396772
rect 137922 396760 137928 396772
rect 130436 396732 137928 396760
rect 130436 396720 130442 396732
rect 137922 396720 137928 396732
rect 137980 396760 137986 396772
rect 180886 396760 180892 396772
rect 137980 396732 180892 396760
rect 137980 396720 137986 396732
rect 180886 396720 180892 396732
rect 180944 396720 180950 396772
rect 258718 396720 258724 396772
rect 258776 396760 258782 396772
rect 276198 396760 276204 396772
rect 258776 396732 276204 396760
rect 258776 396720 258782 396732
rect 276198 396720 276204 396732
rect 276256 396720 276262 396772
rect 60734 396040 60740 396092
rect 60792 396080 60798 396092
rect 61930 396080 61936 396092
rect 60792 396052 61936 396080
rect 60792 396040 60798 396052
rect 61930 396040 61936 396052
rect 61988 396080 61994 396092
rect 66254 396080 66260 396092
rect 61988 396052 66260 396080
rect 61988 396040 61994 396052
rect 66254 396040 66260 396052
rect 66312 396040 66318 396092
rect 115842 396040 115848 396092
rect 115900 396080 115906 396092
rect 124950 396080 124956 396092
rect 115900 396052 124956 396080
rect 115900 396040 115906 396052
rect 124950 396040 124956 396052
rect 125008 396040 125014 396092
rect 162118 396040 162124 396092
rect 162176 396080 162182 396092
rect 192662 396080 192668 396092
rect 162176 396052 192668 396080
rect 162176 396040 162182 396052
rect 192662 396040 192668 396052
rect 192720 396040 192726 396092
rect 153010 395972 153016 396024
rect 153068 396012 153074 396024
rect 156598 396012 156604 396024
rect 153068 395984 156604 396012
rect 153068 395972 153074 395984
rect 156598 395972 156604 395984
rect 156656 395972 156662 396024
rect 162210 395972 162216 396024
rect 162268 396012 162274 396024
rect 170858 396012 170864 396024
rect 162268 395984 170864 396012
rect 162268 395972 162274 395984
rect 170858 395972 170864 395984
rect 170916 396012 170922 396024
rect 191742 396012 191748 396024
rect 170916 395984 191748 396012
rect 170916 395972 170922 395984
rect 191742 395972 191748 395984
rect 191800 395972 191806 396024
rect 258994 395292 259000 395344
rect 259052 395332 259058 395344
rect 273438 395332 273444 395344
rect 259052 395304 273444 395332
rect 259052 395292 259058 395304
rect 273438 395292 273444 395304
rect 273496 395292 273502 395344
rect 115842 394748 115848 394800
rect 115900 394788 115906 394800
rect 144178 394788 144184 394800
rect 115900 394760 144184 394788
rect 115900 394748 115906 394760
rect 144178 394748 144184 394760
rect 144236 394748 144242 394800
rect 153010 394720 153016 394732
rect 115952 394692 153016 394720
rect 115842 394612 115848 394664
rect 115900 394652 115906 394664
rect 115952 394652 115980 394692
rect 153010 394680 153016 394692
rect 153068 394680 153074 394732
rect 255406 394680 255412 394732
rect 255464 394720 255470 394732
rect 272150 394720 272156 394732
rect 255464 394692 272156 394720
rect 255464 394680 255470 394692
rect 272150 394680 272156 394692
rect 272208 394680 272214 394732
rect 115900 394624 115980 394652
rect 115900 394612 115906 394624
rect 117222 394000 117228 394052
rect 117280 394040 117286 394052
rect 136634 394040 136640 394052
rect 117280 394012 136640 394040
rect 117280 394000 117286 394012
rect 136634 394000 136640 394012
rect 136692 394000 136698 394052
rect 137278 394000 137284 394052
rect 137336 394040 137342 394052
rect 159358 394040 159364 394052
rect 137336 394012 159364 394040
rect 137336 394000 137342 394012
rect 159358 394000 159364 394012
rect 159416 394000 159422 394052
rect 118602 393932 118608 393984
rect 118660 393972 118666 393984
rect 163866 393972 163872 393984
rect 118660 393944 163872 393972
rect 118660 393932 118666 393944
rect 163866 393932 163872 393944
rect 163924 393972 163930 393984
rect 171962 393972 171968 393984
rect 163924 393944 171968 393972
rect 163924 393932 163930 393944
rect 171962 393932 171968 393944
rect 172020 393932 172026 393984
rect 178678 393932 178684 393984
rect 178736 393972 178742 393984
rect 187970 393972 187976 393984
rect 178736 393944 187976 393972
rect 178736 393932 178742 393944
rect 187970 393932 187976 393944
rect 188028 393932 188034 393984
rect 256694 393932 256700 393984
rect 256752 393972 256758 393984
rect 278866 393972 278872 393984
rect 256752 393944 278872 393972
rect 256752 393932 256758 393944
rect 278866 393932 278872 393944
rect 278924 393932 278930 393984
rect 60550 393320 60556 393372
rect 60608 393360 60614 393372
rect 67726 393360 67732 393372
rect 60608 393332 67732 393360
rect 60608 393320 60614 393332
rect 67726 393320 67732 393332
rect 67784 393320 67790 393372
rect 166350 393320 166356 393372
rect 166408 393360 166414 393372
rect 177482 393360 177488 393372
rect 166408 393332 177488 393360
rect 166408 393320 166414 393332
rect 177482 393320 177488 393332
rect 177540 393320 177546 393372
rect 255406 393320 255412 393372
rect 255464 393360 255470 393372
rect 278866 393360 278872 393372
rect 255464 393332 278872 393360
rect 255464 393320 255470 393332
rect 278866 393320 278872 393332
rect 278924 393320 278930 393372
rect 115934 392708 115940 392760
rect 115992 392748 115998 392760
rect 117222 392748 117228 392760
rect 115992 392720 117228 392748
rect 115992 392708 115998 392720
rect 117222 392708 117228 392720
rect 117280 392708 117286 392760
rect 142982 392572 142988 392624
rect 143040 392612 143046 392624
rect 158530 392612 158536 392624
rect 143040 392584 158536 392612
rect 143040 392572 143046 392584
rect 158530 392572 158536 392584
rect 158588 392612 158594 392624
rect 179414 392612 179420 392624
rect 158588 392584 179420 392612
rect 158588 392572 158594 392584
rect 179414 392572 179420 392584
rect 179472 392572 179478 392624
rect 254026 392096 254032 392148
rect 254084 392136 254090 392148
rect 255498 392136 255504 392148
rect 254084 392108 255504 392136
rect 254084 392096 254090 392108
rect 255498 392096 255504 392108
rect 255556 392096 255562 392148
rect 60550 391960 60556 392012
rect 60608 392000 60614 392012
rect 66622 392000 66628 392012
rect 60608 391972 66628 392000
rect 60608 391960 60614 391972
rect 66622 391960 66628 391972
rect 66680 391960 66686 392012
rect 115842 391960 115848 392012
rect 115900 392000 115906 392012
rect 141602 392000 141608 392012
rect 115900 391972 141608 392000
rect 115900 391960 115906 391972
rect 141602 391960 141608 391972
rect 141660 391960 141666 392012
rect 168190 391960 168196 392012
rect 168248 392000 168254 392012
rect 186314 392000 186320 392012
rect 168248 391972 186320 392000
rect 168248 391960 168254 391972
rect 186314 391960 186320 391972
rect 186372 391960 186378 392012
rect 68554 391892 68560 391944
rect 68612 391932 68618 391944
rect 161198 391932 161204 391944
rect 68612 391904 161204 391932
rect 68612 391892 68618 391904
rect 161198 391892 161204 391904
rect 161256 391892 161262 391944
rect 177482 391280 177488 391332
rect 177540 391320 177546 391332
rect 193214 391320 193220 391332
rect 177540 391292 193220 391320
rect 177540 391280 177546 391292
rect 193214 391280 193220 391292
rect 193272 391280 193278 391332
rect 259270 391280 259276 391332
rect 259328 391320 259334 391332
rect 298186 391320 298192 391332
rect 259328 391292 298192 391320
rect 259328 391280 259334 391292
rect 298186 391280 298192 391292
rect 298244 391280 298250 391332
rect 43438 391212 43444 391264
rect 43496 391252 43502 391264
rect 43496 391224 80054 391252
rect 43496 391212 43502 391224
rect 80026 390980 80054 391224
rect 189718 391212 189724 391264
rect 189776 391252 189782 391264
rect 273898 391252 273904 391264
rect 189776 391224 200114 391252
rect 189776 391212 189782 391224
rect 93946 390980 93952 390992
rect 80026 390952 93952 390980
rect 93946 390940 93952 390952
rect 94004 390940 94010 390992
rect 193214 390940 193220 390992
rect 193272 390980 193278 390992
rect 194134 390980 194140 390992
rect 193272 390952 194140 390980
rect 193272 390940 193278 390952
rect 194134 390940 194140 390952
rect 194192 390940 194198 390992
rect 200086 390980 200114 391224
rect 258046 391224 273904 391252
rect 218330 390980 218336 390992
rect 200086 390952 218336 390980
rect 218330 390940 218336 390952
rect 218388 390980 218394 390992
rect 218790 390980 218796 390992
rect 218388 390952 218796 390980
rect 218388 390940 218394 390952
rect 218790 390940 218796 390952
rect 218848 390940 218854 390992
rect 251726 390940 251732 390992
rect 251784 390980 251790 390992
rect 258046 390980 258074 391224
rect 273898 391212 273904 391224
rect 273956 391212 273962 391264
rect 283558 391212 283564 391264
rect 283616 391252 283622 391264
rect 291470 391252 291476 391264
rect 283616 391224 291476 391252
rect 283616 391212 283622 391224
rect 291470 391212 291476 391224
rect 291528 391252 291534 391264
rect 582374 391252 582380 391264
rect 291528 391224 582380 391252
rect 291528 391212 291534 391224
rect 582374 391212 582380 391224
rect 582432 391212 582438 391264
rect 251784 390952 258074 390980
rect 251784 390940 251790 390952
rect 89898 390600 89904 390652
rect 89956 390640 89962 390652
rect 90450 390640 90456 390652
rect 89956 390612 90456 390640
rect 89956 390600 89962 390612
rect 90450 390600 90456 390612
rect 90508 390600 90514 390652
rect 100386 390532 100392 390584
rect 100444 390572 100450 390584
rect 179138 390572 179144 390584
rect 100444 390544 179144 390572
rect 100444 390532 100450 390544
rect 179138 390532 179144 390544
rect 179196 390572 179202 390584
rect 179506 390572 179512 390584
rect 179196 390544 179512 390572
rect 179196 390532 179202 390544
rect 179506 390532 179512 390544
rect 179564 390532 179570 390584
rect 67818 390124 67824 390176
rect 67876 390164 67882 390176
rect 68784 390164 68790 390176
rect 67876 390136 68790 390164
rect 67876 390124 67882 390136
rect 68784 390124 68790 390136
rect 68842 390124 68848 390176
rect 96706 390124 96712 390176
rect 96764 390164 96770 390176
rect 97856 390164 97862 390176
rect 96764 390136 97862 390164
rect 96764 390124 96770 390136
rect 97856 390124 97862 390136
rect 97914 390124 97920 390176
rect 100800 390124 100806 390176
rect 100858 390164 100864 390176
rect 101950 390164 101956 390176
rect 100858 390136 101956 390164
rect 100858 390124 100864 390136
rect 101950 390124 101956 390136
rect 102008 390124 102014 390176
rect 104802 389784 104808 389836
rect 104860 389824 104866 389836
rect 114830 389824 114836 389836
rect 104860 389796 114836 389824
rect 104860 389784 104866 389796
rect 114830 389784 114836 389796
rect 114888 389784 114894 389836
rect 156690 389784 156696 389836
rect 156748 389824 156754 389836
rect 168374 389824 168380 389836
rect 156748 389796 168380 389824
rect 156748 389784 156754 389796
rect 168374 389784 168380 389796
rect 168432 389784 168438 389836
rect 179230 389784 179236 389836
rect 179288 389824 179294 389836
rect 180886 389824 180892 389836
rect 179288 389796 180892 389824
rect 179288 389784 179294 389796
rect 180886 389784 180892 389796
rect 180944 389784 180950 389836
rect 277302 389784 277308 389836
rect 277360 389824 277366 389836
rect 281534 389824 281540 389836
rect 277360 389796 281540 389824
rect 277360 389784 277366 389796
rect 281534 389784 281540 389796
rect 281592 389784 281598 389836
rect 36538 389240 36544 389292
rect 36596 389280 36602 389292
rect 100754 389280 100760 389292
rect 36596 389252 100760 389280
rect 36596 389240 36602 389252
rect 100754 389240 100760 389252
rect 100812 389240 100818 389292
rect 168374 389240 168380 389292
rect 168432 389280 168438 389292
rect 169478 389280 169484 389292
rect 168432 389252 169484 389280
rect 168432 389240 168438 389252
rect 169478 389240 169484 389252
rect 169536 389280 169542 389292
rect 202046 389280 202052 389292
rect 169536 389252 202052 389280
rect 169536 389240 169542 389252
rect 202046 389240 202052 389252
rect 202104 389240 202110 389292
rect 230566 389240 230572 389292
rect 230624 389280 230630 389292
rect 256694 389280 256700 389292
rect 230624 389252 256700 389280
rect 230624 389240 230630 389252
rect 256694 389240 256700 389252
rect 256752 389240 256758 389292
rect 3510 389172 3516 389224
rect 3568 389212 3574 389224
rect 107654 389212 107660 389224
rect 3568 389184 107660 389212
rect 3568 389172 3574 389184
rect 107654 389172 107660 389184
rect 107712 389212 107718 389224
rect 118602 389212 118608 389224
rect 107712 389184 118608 389212
rect 107712 389172 107718 389184
rect 118602 389172 118608 389184
rect 118660 389172 118666 389224
rect 187970 389172 187976 389224
rect 188028 389212 188034 389224
rect 240134 389212 240140 389224
rect 188028 389184 240140 389212
rect 188028 389172 188034 389184
rect 240134 389172 240140 389184
rect 240192 389212 240198 389224
rect 241054 389212 241060 389224
rect 240192 389184 241060 389212
rect 240192 389172 240198 389184
rect 241054 389172 241060 389184
rect 241112 389172 241118 389224
rect 241514 389172 241520 389224
rect 241572 389212 241578 389224
rect 264238 389212 264244 389224
rect 241572 389184 264244 389212
rect 241572 389172 241578 389184
rect 264238 389172 264244 389184
rect 264296 389172 264302 389224
rect 157150 389104 157156 389156
rect 157208 389144 157214 389156
rect 161566 389144 161572 389156
rect 157208 389116 161572 389144
rect 157208 389104 157214 389116
rect 161566 389104 161572 389116
rect 161624 389104 161630 389156
rect 176378 389104 176384 389156
rect 176436 389144 176442 389156
rect 197262 389144 197268 389156
rect 176436 389116 197268 389144
rect 176436 389104 176442 389116
rect 197262 389104 197268 389116
rect 197320 389104 197326 389156
rect 250438 389104 250444 389156
rect 250496 389144 250502 389156
rect 281626 389144 281632 389156
rect 250496 389116 281632 389144
rect 250496 389104 250502 389116
rect 281626 389104 281632 389116
rect 281684 389104 281690 389156
rect 253382 389036 253388 389088
rect 253440 389076 253446 389088
rect 271966 389076 271972 389088
rect 253440 389048 271972 389076
rect 253440 389036 253446 389048
rect 271966 389036 271972 389048
rect 272024 389036 272030 389088
rect 59170 388424 59176 388476
rect 59228 388464 59234 388476
rect 71682 388464 71688 388476
rect 59228 388436 71688 388464
rect 59228 388424 59234 388436
rect 71682 388424 71688 388436
rect 71740 388424 71746 388476
rect 72326 388424 72332 388476
rect 72384 388464 72390 388476
rect 128354 388464 128360 388476
rect 72384 388436 128360 388464
rect 72384 388424 72390 388436
rect 128354 388424 128360 388436
rect 128412 388424 128418 388476
rect 180610 388424 180616 388476
rect 180668 388464 180674 388476
rect 184842 388464 184848 388476
rect 180668 388436 184848 388464
rect 180668 388424 180674 388436
rect 184842 388424 184848 388436
rect 184900 388424 184906 388476
rect 93946 388288 93952 388340
rect 94004 388328 94010 388340
rect 94222 388328 94228 388340
rect 94004 388300 94228 388328
rect 94004 388288 94010 388300
rect 94222 388288 94228 388300
rect 94280 388288 94286 388340
rect 232590 387948 232596 388000
rect 232648 387988 232654 388000
rect 236270 387988 236276 388000
rect 232648 387960 236276 387988
rect 232648 387948 232654 387960
rect 236270 387948 236276 387960
rect 236328 387948 236334 388000
rect 166258 387880 166264 387932
rect 166316 387920 166322 387932
rect 167730 387920 167736 387932
rect 166316 387892 167736 387920
rect 166316 387880 166322 387892
rect 167730 387880 167736 387892
rect 167788 387880 167794 387932
rect 231210 387880 231216 387932
rect 231268 387920 231274 387932
rect 234246 387920 234252 387932
rect 231268 387892 234252 387920
rect 231268 387880 231274 387892
rect 234246 387880 234252 387892
rect 234304 387880 234310 387932
rect 71682 387812 71688 387864
rect 71740 387852 71746 387864
rect 72510 387852 72516 387864
rect 71740 387824 72516 387852
rect 71740 387812 71746 387824
rect 72510 387812 72516 387824
rect 72568 387812 72574 387864
rect 128354 387812 128360 387864
rect 128412 387852 128418 387864
rect 128998 387852 129004 387864
rect 128412 387824 129004 387852
rect 128412 387812 128418 387824
rect 128998 387812 129004 387824
rect 129056 387852 129062 387864
rect 173618 387852 173624 387864
rect 129056 387824 173624 387852
rect 129056 387812 129062 387824
rect 173618 387812 173624 387824
rect 173676 387812 173682 387864
rect 196066 387812 196072 387864
rect 196124 387852 196130 387864
rect 197262 387852 197268 387864
rect 196124 387824 197268 387852
rect 196124 387812 196130 387824
rect 197262 387812 197268 387824
rect 197320 387812 197326 387864
rect 221458 387812 221464 387864
rect 221516 387852 221522 387864
rect 223942 387852 223948 387864
rect 221516 387824 223948 387852
rect 221516 387812 221522 387824
rect 223942 387812 223948 387824
rect 224000 387812 224006 387864
rect 233326 387812 233332 387864
rect 233384 387852 233390 387864
rect 235258 387852 235264 387864
rect 233384 387824 235264 387852
rect 233384 387812 233390 387824
rect 235258 387812 235264 387824
rect 235316 387812 235322 387864
rect 249150 387812 249156 387864
rect 249208 387852 249214 387864
rect 252278 387852 252284 387864
rect 249208 387824 252284 387852
rect 249208 387812 249214 387824
rect 252278 387812 252284 387824
rect 252336 387812 252342 387864
rect 103882 387744 103888 387796
rect 103940 387784 103946 387796
rect 126238 387784 126244 387796
rect 103940 387756 126244 387784
rect 103940 387744 103946 387756
rect 126238 387744 126244 387756
rect 126296 387744 126302 387796
rect 187418 387744 187424 387796
rect 187476 387784 187482 387796
rect 188430 387784 188436 387796
rect 187476 387756 188436 387784
rect 187476 387744 187482 387756
rect 188430 387744 188436 387756
rect 188488 387744 188494 387796
rect 188522 387744 188528 387796
rect 188580 387784 188586 387796
rect 215938 387784 215944 387796
rect 188580 387756 215944 387784
rect 188580 387744 188586 387756
rect 215938 387744 215944 387756
rect 215996 387744 216002 387796
rect 238110 387744 238116 387796
rect 238168 387784 238174 387796
rect 284294 387784 284300 387796
rect 238168 387756 284300 387784
rect 238168 387744 238174 387756
rect 284294 387744 284300 387756
rect 284352 387744 284358 387796
rect 184382 387676 184388 387728
rect 184440 387716 184446 387728
rect 184842 387716 184848 387728
rect 184440 387688 184848 387716
rect 184440 387676 184446 387688
rect 184842 387676 184848 387688
rect 184900 387716 184906 387728
rect 202966 387716 202972 387728
rect 184900 387688 202972 387716
rect 184900 387676 184906 387688
rect 202966 387676 202972 387688
rect 203024 387676 203030 387728
rect 149698 387132 149704 387184
rect 149756 387172 149762 387184
rect 168190 387172 168196 387184
rect 149756 387144 168196 387172
rect 149756 387132 149762 387144
rect 168190 387132 168196 387144
rect 168248 387132 168254 387184
rect 86862 387064 86868 387116
rect 86920 387104 86926 387116
rect 106182 387104 106188 387116
rect 86920 387076 106188 387104
rect 86920 387064 86926 387076
rect 106182 387064 106188 387076
rect 106240 387064 106246 387116
rect 110414 387064 110420 387116
rect 110472 387104 110478 387116
rect 187142 387104 187148 387116
rect 110472 387076 187148 387104
rect 110472 387064 110478 387076
rect 187142 387064 187148 387076
rect 187200 387064 187206 387116
rect 228358 387064 228364 387116
rect 228416 387104 228422 387116
rect 253382 387104 253388 387116
rect 228416 387076 253388 387104
rect 228416 387064 228422 387076
rect 253382 387064 253388 387076
rect 253440 387064 253446 387116
rect 265710 387064 265716 387116
rect 265768 387104 265774 387116
rect 582374 387104 582380 387116
rect 265768 387076 582380 387104
rect 265768 387064 265774 387076
rect 582374 387064 582380 387076
rect 582432 387064 582438 387116
rect 69014 386996 69020 387048
rect 69072 387036 69078 387048
rect 69750 387036 69756 387048
rect 69072 387008 69756 387036
rect 69072 386996 69078 387008
rect 69750 386996 69756 387008
rect 69808 386996 69814 387048
rect 70394 386996 70400 387048
rect 70452 387036 70458 387048
rect 71222 387036 71228 387048
rect 70452 387008 71228 387036
rect 70452 386996 70458 387008
rect 71222 386996 71228 387008
rect 71280 386996 71286 387048
rect 74534 386996 74540 387048
rect 74592 387036 74598 387048
rect 75270 387036 75276 387048
rect 74592 387008 75276 387036
rect 74592 386996 74598 387008
rect 75270 386996 75276 387008
rect 75328 386996 75334 387048
rect 78674 386996 78680 387048
rect 78732 387036 78738 387048
rect 79502 387036 79508 387048
rect 78732 387008 79508 387036
rect 78732 386996 78738 387008
rect 79502 386996 79508 387008
rect 79560 386996 79566 387048
rect 109034 386996 109040 387048
rect 109092 387036 109098 387048
rect 109494 387036 109500 387048
rect 109092 387008 109500 387036
rect 109092 386996 109098 387008
rect 109494 386996 109500 387008
rect 109552 386996 109558 387048
rect 205634 386996 205640 387048
rect 205692 387036 205698 387048
rect 206462 387036 206468 387048
rect 205692 387008 206468 387036
rect 205692 386996 205698 387008
rect 206462 386996 206468 387008
rect 206520 386996 206526 387048
rect 208394 386996 208400 387048
rect 208452 387036 208458 387048
rect 209222 387036 209228 387048
rect 208452 387008 209228 387036
rect 208452 386996 208458 387008
rect 209222 386996 209228 387008
rect 209280 386996 209286 387048
rect 83182 386928 83188 386980
rect 83240 386968 83246 386980
rect 84102 386968 84108 386980
rect 83240 386940 84108 386968
rect 83240 386928 83246 386940
rect 84102 386928 84108 386940
rect 84160 386928 84166 386980
rect 93946 386860 93952 386912
rect 94004 386900 94010 386912
rect 94774 386900 94780 386912
rect 94004 386872 94780 386900
rect 94004 386860 94010 386872
rect 94774 386860 94780 386872
rect 94832 386860 94838 386912
rect 124858 386356 124864 386368
rect 93826 386328 124864 386356
rect 85114 386248 85120 386300
rect 85172 386288 85178 386300
rect 93826 386288 93854 386328
rect 124858 386316 124864 386328
rect 124916 386316 124922 386368
rect 194134 386316 194140 386368
rect 194192 386356 194198 386368
rect 252554 386356 252560 386368
rect 194192 386328 252560 386356
rect 194192 386316 194198 386328
rect 252554 386316 252560 386328
rect 252612 386316 252618 386368
rect 85172 386260 93854 386288
rect 85172 386248 85178 386260
rect 224862 386248 224868 386300
rect 224920 386288 224926 386300
rect 258718 386288 258724 386300
rect 224920 386260 258724 386288
rect 224920 386248 224926 386260
rect 258718 386248 258724 386260
rect 258776 386248 258782 386300
rect 85390 385840 85396 385892
rect 85448 385880 85454 385892
rect 88426 385880 88432 385892
rect 85448 385852 88432 385880
rect 85448 385840 85454 385852
rect 88426 385840 88432 385852
rect 88484 385840 88490 385892
rect 77202 385772 77208 385824
rect 77260 385812 77266 385824
rect 78030 385812 78036 385824
rect 77260 385784 78036 385812
rect 77260 385772 77266 385784
rect 78030 385772 78036 385784
rect 78088 385772 78094 385824
rect 141970 385704 141976 385756
rect 142028 385744 142034 385756
rect 147030 385744 147036 385756
rect 142028 385716 147036 385744
rect 142028 385704 142034 385716
rect 147030 385704 147036 385716
rect 147088 385704 147094 385756
rect 99558 385636 99564 385688
rect 99616 385676 99622 385688
rect 170490 385676 170496 385688
rect 99616 385648 170496 385676
rect 99616 385636 99622 385648
rect 170490 385636 170496 385648
rect 170548 385636 170554 385688
rect 177390 385636 177396 385688
rect 177448 385676 177454 385688
rect 180058 385676 180064 385688
rect 177448 385648 180064 385676
rect 177448 385636 177454 385648
rect 180058 385636 180064 385648
rect 180116 385676 180122 385688
rect 195882 385676 195888 385688
rect 180116 385648 195888 385676
rect 180116 385636 180122 385648
rect 195882 385636 195888 385648
rect 195940 385636 195946 385688
rect 266998 385636 267004 385688
rect 267056 385676 267062 385688
rect 270494 385676 270500 385688
rect 267056 385648 270500 385676
rect 267056 385636 267062 385648
rect 270494 385636 270500 385648
rect 270552 385636 270558 385688
rect 188982 385364 188988 385416
rect 189040 385404 189046 385416
rect 191190 385404 191196 385416
rect 189040 385376 191196 385404
rect 189040 385364 189046 385376
rect 191190 385364 191196 385376
rect 191248 385364 191254 385416
rect 158070 385024 158076 385076
rect 158128 385064 158134 385076
rect 162118 385064 162124 385076
rect 158128 385036 162124 385064
rect 158128 385024 158134 385036
rect 162118 385024 162124 385036
rect 162176 385024 162182 385076
rect 185578 384956 185584 385008
rect 185636 384996 185642 385008
rect 215294 384996 215300 385008
rect 185636 384968 215300 384996
rect 185636 384956 185642 384968
rect 215294 384956 215300 384968
rect 215352 384956 215358 385008
rect 239398 384956 239404 385008
rect 239456 384996 239462 385008
rect 251726 384996 251732 385008
rect 239456 384968 251732 384996
rect 239456 384956 239462 384968
rect 251726 384956 251732 384968
rect 251784 384956 251790 385008
rect 251818 384956 251824 385008
rect 251876 384996 251882 385008
rect 254026 384996 254032 385008
rect 251876 384968 254032 384996
rect 251876 384956 251882 384968
rect 254026 384956 254032 384968
rect 254084 384956 254090 385008
rect 192570 384888 192576 384940
rect 192628 384928 192634 384940
rect 222838 384928 222844 384940
rect 192628 384900 222844 384928
rect 192628 384888 192634 384900
rect 222838 384888 222844 384900
rect 222896 384888 222902 384940
rect 226426 384344 226432 384396
rect 226484 384384 226490 384396
rect 227622 384384 227628 384396
rect 226484 384356 227628 384384
rect 226484 384344 226490 384356
rect 227622 384344 227628 384356
rect 227680 384344 227686 384396
rect 73798 384276 73804 384328
rect 73856 384316 73862 384328
rect 93118 384316 93124 384328
rect 73856 384288 93124 384316
rect 73856 384276 73862 384288
rect 93118 384276 93124 384288
rect 93176 384276 93182 384328
rect 215294 384276 215300 384328
rect 215352 384316 215358 384328
rect 216030 384316 216036 384328
rect 215352 384288 216036 384316
rect 215352 384276 215358 384288
rect 216030 384276 216036 384288
rect 216088 384276 216094 384328
rect 106182 383732 106188 383784
rect 106240 383772 106246 383784
rect 150434 383772 150440 383784
rect 106240 383744 150440 383772
rect 106240 383732 106246 383744
rect 150434 383732 150440 383744
rect 150492 383732 150498 383784
rect 3510 383664 3516 383716
rect 3568 383704 3574 383716
rect 113450 383704 113456 383716
rect 3568 383676 113456 383704
rect 3568 383664 3574 383676
rect 113450 383664 113456 383676
rect 113508 383664 113514 383716
rect 150250 383664 150256 383716
rect 150308 383704 150314 383716
rect 153930 383704 153936 383716
rect 150308 383676 153936 383704
rect 150308 383664 150314 383676
rect 153930 383664 153936 383676
rect 153988 383664 153994 383716
rect 227622 383664 227628 383716
rect 227680 383704 227686 383716
rect 280154 383704 280160 383716
rect 227680 383676 280160 383704
rect 227680 383664 227686 383676
rect 280154 383664 280160 383676
rect 280212 383664 280218 383716
rect 109126 382984 109132 383036
rect 109184 383024 109190 383036
rect 126238 383024 126244 383036
rect 109184 382996 126244 383024
rect 109184 382984 109190 382996
rect 126238 382984 126244 382996
rect 126296 382984 126302 383036
rect 175182 382984 175188 383036
rect 175240 383024 175246 383036
rect 182082 383024 182088 383036
rect 175240 382996 182088 383024
rect 175240 382984 175246 382996
rect 182082 382984 182088 382996
rect 182140 383024 182146 383036
rect 208486 383024 208492 383036
rect 182140 382996 208492 383024
rect 182140 382984 182146 382996
rect 208486 382984 208492 382996
rect 208544 382984 208550 383036
rect 252462 382984 252468 383036
rect 252520 383024 252526 383036
rect 263686 383024 263692 383036
rect 252520 382996 263692 383024
rect 252520 382984 252526 382996
rect 263686 382984 263692 382996
rect 263744 382984 263750 383036
rect 97718 382916 97724 382968
rect 97776 382956 97782 382968
rect 124214 382956 124220 382968
rect 97776 382928 124220 382956
rect 97776 382916 97782 382928
rect 124214 382916 124220 382928
rect 124272 382956 124278 382968
rect 231854 382956 231860 382968
rect 124272 382928 231860 382956
rect 124272 382916 124278 382928
rect 231854 382916 231860 382928
rect 231912 382956 231918 382968
rect 281626 382956 281632 382968
rect 231912 382928 281632 382956
rect 231912 382916 231918 382928
rect 281626 382916 281632 382928
rect 281684 382916 281690 382968
rect 67358 382168 67364 382220
rect 67416 382208 67422 382220
rect 150802 382208 150808 382220
rect 67416 382180 150808 382208
rect 67416 382168 67422 382180
rect 150802 382168 150808 382180
rect 150860 382208 150866 382220
rect 151078 382208 151084 382220
rect 150860 382180 151084 382208
rect 150860 382168 150866 382180
rect 151078 382168 151084 382180
rect 151136 382168 151142 382220
rect 177850 382168 177856 382220
rect 177908 382208 177914 382220
rect 211154 382208 211160 382220
rect 177908 382180 211160 382208
rect 177908 382168 177914 382180
rect 211154 382168 211160 382180
rect 211212 382168 211218 382220
rect 102042 381488 102048 381540
rect 102100 381528 102106 381540
rect 113358 381528 113364 381540
rect 102100 381500 113364 381528
rect 102100 381488 102106 381500
rect 113358 381488 113364 381500
rect 113416 381488 113422 381540
rect 150802 381488 150808 381540
rect 150860 381528 150866 381540
rect 158714 381528 158720 381540
rect 150860 381500 158720 381528
rect 150860 381488 150866 381500
rect 158714 381488 158720 381500
rect 158772 381488 158778 381540
rect 173618 381488 173624 381540
rect 173676 381528 173682 381540
rect 216674 381528 216680 381540
rect 173676 381500 216680 381528
rect 173676 381488 173682 381500
rect 216674 381488 216680 381500
rect 216732 381488 216738 381540
rect 227622 381488 227628 381540
rect 227680 381528 227686 381540
rect 256786 381528 256792 381540
rect 227680 381500 256792 381528
rect 227680 381488 227686 381500
rect 256786 381488 256792 381500
rect 256844 381488 256850 381540
rect 211154 380876 211160 380928
rect 211212 380916 211218 380928
rect 211798 380916 211804 380928
rect 211212 380888 211804 380916
rect 211212 380876 211218 380888
rect 211798 380876 211804 380888
rect 211856 380876 211862 380928
rect 231118 380876 231124 380928
rect 231176 380916 231182 380928
rect 277670 380916 277676 380928
rect 231176 380888 277676 380916
rect 231176 380876 231182 380888
rect 277670 380876 277676 380888
rect 277728 380876 277734 380928
rect 48130 380808 48136 380860
rect 48188 380848 48194 380860
rect 154022 380848 154028 380860
rect 48188 380820 154028 380848
rect 48188 380808 48194 380820
rect 154022 380808 154028 380820
rect 154080 380808 154086 380860
rect 236362 380808 236368 380860
rect 236420 380848 236426 380860
rect 236638 380848 236644 380860
rect 236420 380820 236644 380848
rect 236420 380808 236426 380820
rect 236638 380808 236644 380820
rect 236696 380848 236702 380860
rect 281718 380848 281724 380860
rect 236696 380820 281724 380848
rect 236696 380808 236702 380820
rect 281718 380808 281724 380820
rect 281776 380808 281782 380860
rect 77294 380740 77300 380792
rect 77352 380780 77358 380792
rect 130378 380780 130384 380792
rect 77352 380752 130384 380780
rect 77352 380740 77358 380752
rect 130378 380740 130384 380752
rect 130436 380740 130442 380792
rect 187694 380196 187700 380248
rect 187752 380236 187758 380248
rect 226426 380236 226432 380248
rect 187752 380208 226432 380236
rect 187752 380196 187758 380208
rect 226426 380196 226432 380208
rect 226484 380196 226490 380248
rect 129734 380128 129740 380180
rect 129792 380168 129798 380180
rect 138750 380168 138756 380180
rect 129792 380140 138756 380168
rect 129792 380128 129798 380140
rect 138750 380128 138756 380140
rect 138808 380168 138814 380180
rect 207014 380168 207020 380180
rect 138808 380140 207020 380168
rect 138808 380128 138814 380140
rect 207014 380128 207020 380140
rect 207072 380128 207078 380180
rect 221550 380128 221556 380180
rect 221608 380168 221614 380180
rect 269390 380168 269396 380180
rect 221608 380140 269396 380168
rect 221608 380128 221614 380140
rect 269390 380128 269396 380140
rect 269448 380168 269454 380180
rect 270678 380168 270684 380180
rect 269448 380140 270684 380168
rect 269448 380128 269454 380140
rect 270678 380128 270684 380140
rect 270736 380128 270742 380180
rect 67266 379448 67272 379500
rect 67324 379488 67330 379500
rect 157334 379488 157340 379500
rect 67324 379460 157340 379488
rect 67324 379448 67330 379460
rect 157334 379448 157340 379460
rect 157392 379448 157398 379500
rect 235258 379448 235264 379500
rect 235316 379488 235322 379500
rect 235902 379488 235908 379500
rect 235316 379460 235908 379488
rect 235316 379448 235322 379460
rect 235902 379448 235908 379460
rect 235960 379488 235966 379500
rect 291286 379488 291292 379500
rect 235960 379460 291292 379488
rect 235960 379448 235966 379460
rect 291286 379448 291292 379460
rect 291344 379448 291350 379500
rect 157334 378972 157340 379024
rect 157392 379012 157398 379024
rect 157978 379012 157984 379024
rect 157392 378984 157984 379012
rect 157392 378972 157398 378984
rect 157978 378972 157984 378984
rect 158036 378972 158042 379024
rect 188430 378836 188436 378888
rect 188488 378876 188494 378888
rect 197446 378876 197452 378888
rect 188488 378848 197452 378876
rect 188488 378836 188494 378848
rect 197446 378836 197452 378848
rect 197504 378836 197510 378888
rect 121638 378768 121644 378820
rect 121696 378808 121702 378820
rect 187694 378808 187700 378820
rect 121696 378780 187700 378808
rect 121696 378768 121702 378780
rect 187694 378768 187700 378780
rect 187752 378768 187758 378820
rect 241422 378768 241428 378820
rect 241480 378808 241486 378820
rect 253934 378808 253940 378820
rect 241480 378780 253940 378808
rect 241480 378768 241486 378780
rect 253934 378768 253940 378780
rect 253992 378768 253998 378820
rect 111978 378088 111984 378140
rect 112036 378128 112042 378140
rect 112438 378128 112444 378140
rect 112036 378100 112444 378128
rect 112036 378088 112042 378100
rect 112438 378088 112444 378100
rect 112496 378128 112502 378140
rect 112496 378100 219434 378128
rect 112496 378088 112502 378100
rect 179230 378020 179236 378072
rect 179288 378060 179294 378072
rect 205726 378060 205732 378072
rect 179288 378032 205732 378060
rect 179288 378020 179294 378032
rect 205726 378020 205732 378032
rect 205784 378020 205790 378072
rect 219406 378060 219434 378100
rect 227806 378088 227812 378140
rect 227864 378128 227870 378140
rect 283190 378128 283196 378140
rect 227864 378100 283196 378128
rect 227864 378088 227870 378100
rect 283190 378088 283196 378100
rect 283248 378088 283254 378140
rect 228358 378060 228364 378072
rect 219406 378032 228364 378060
rect 228358 378020 228364 378032
rect 228416 378020 228422 378072
rect 243078 378020 243084 378072
rect 243136 378060 243142 378072
rect 262214 378060 262220 378072
rect 243136 378032 262220 378060
rect 243136 378020 243142 378032
rect 262214 378020 262220 378032
rect 262272 378060 262278 378072
rect 262858 378060 262864 378072
rect 262272 378032 262864 378060
rect 262272 378020 262278 378032
rect 262858 378020 262864 378032
rect 262916 378020 262922 378072
rect 97626 377408 97632 377460
rect 97684 377448 97690 377460
rect 130378 377448 130384 377460
rect 97684 377420 130384 377448
rect 97684 377408 97690 377420
rect 130378 377408 130384 377420
rect 130436 377408 130442 377460
rect 94222 376660 94228 376712
rect 94280 376700 94286 376712
rect 121638 376700 121644 376712
rect 94280 376672 121644 376700
rect 94280 376660 94286 376672
rect 121638 376660 121644 376672
rect 121696 376660 121702 376712
rect 148962 376660 148968 376712
rect 149020 376700 149026 376712
rect 251266 376700 251272 376712
rect 149020 376672 251272 376700
rect 149020 376660 149026 376672
rect 251266 376660 251272 376672
rect 251324 376660 251330 376712
rect 108942 375980 108948 376032
rect 109000 376020 109006 376032
rect 116118 376020 116124 376032
rect 109000 375992 116124 376020
rect 109000 375980 109006 375992
rect 116118 375980 116124 375992
rect 116176 375980 116182 376032
rect 245746 375408 245752 375420
rect 245659 375380 245752 375408
rect 88242 375300 88248 375352
rect 88300 375340 88306 375352
rect 91922 375340 91928 375352
rect 88300 375312 91928 375340
rect 88300 375300 88306 375312
rect 91922 375300 91928 375312
rect 91980 375340 91986 375352
rect 213178 375340 213184 375352
rect 91980 375312 213184 375340
rect 91980 375300 91986 375312
rect 213178 375300 213184 375312
rect 213236 375300 213242 375352
rect 245672 375340 245700 375380
rect 245746 375368 245752 375380
rect 245804 375408 245810 375420
rect 263962 375408 263968 375420
rect 245804 375380 263968 375408
rect 245804 375368 245810 375380
rect 263962 375368 263968 375380
rect 264020 375368 264026 375420
rect 238726 375312 245700 375340
rect 171962 375232 171968 375284
rect 172020 375272 172026 375284
rect 238726 375272 238754 375312
rect 172020 375244 238754 375272
rect 172020 375232 172026 375244
rect 218054 374008 218060 374060
rect 218112 374048 218118 374060
rect 265158 374048 265164 374060
rect 218112 374020 265164 374048
rect 218112 374008 218118 374020
rect 265158 374008 265164 374020
rect 265216 374008 265222 374060
rect 82814 373940 82820 373992
rect 82872 373980 82878 373992
rect 82872 373952 142154 373980
rect 82872 373940 82878 373952
rect 142126 373912 142154 373952
rect 187142 373940 187148 373992
rect 187200 373980 187206 373992
rect 250438 373980 250444 373992
rect 187200 373952 250444 373980
rect 187200 373940 187206 373952
rect 250438 373940 250444 373952
rect 250496 373940 250502 373992
rect 161566 373912 161572 373924
rect 142126 373884 161572 373912
rect 161566 373872 161572 373884
rect 161624 373912 161630 373924
rect 162762 373912 162768 373924
rect 161624 373884 162768 373912
rect 161624 373872 161630 373884
rect 162762 373872 162768 373884
rect 162820 373912 162826 373924
rect 213914 373912 213920 373924
rect 162820 373884 213920 373912
rect 162820 373872 162826 373884
rect 213914 373872 213920 373884
rect 213972 373872 213978 373924
rect 187142 373396 187148 373448
rect 187200 373436 187206 373448
rect 187602 373436 187608 373448
rect 187200 373408 187608 373436
rect 187200 373396 187206 373408
rect 187602 373396 187608 373408
rect 187660 373396 187666 373448
rect 107562 373260 107568 373312
rect 107620 373300 107626 373312
rect 115934 373300 115940 373312
rect 107620 373272 115940 373300
rect 107620 373260 107626 373272
rect 115934 373260 115940 373272
rect 115992 373260 115998 373312
rect 242342 373260 242348 373312
rect 242400 373300 242406 373312
rect 263778 373300 263784 373312
rect 242400 373272 263784 373300
rect 242400 373260 242406 373272
rect 263778 373260 263784 373272
rect 263836 373260 263842 373312
rect 137830 372716 137836 372768
rect 137888 372756 137894 372768
rect 141510 372756 141516 372768
rect 137888 372728 141516 372756
rect 137888 372716 137894 372728
rect 141510 372716 141516 372728
rect 141568 372716 141574 372768
rect 61930 372512 61936 372564
rect 61988 372552 61994 372564
rect 169754 372552 169760 372564
rect 61988 372524 169760 372552
rect 61988 372512 61994 372524
rect 169754 372512 169760 372524
rect 169812 372512 169818 372564
rect 188338 372512 188344 372564
rect 188396 372552 188402 372564
rect 273254 372552 273260 372564
rect 188396 372524 273260 372552
rect 188396 372512 188402 372524
rect 273254 372512 273260 372524
rect 273312 372512 273318 372564
rect 93946 372444 93952 372496
rect 94004 372484 94010 372496
rect 141234 372484 141240 372496
rect 94004 372456 141240 372484
rect 94004 372444 94010 372456
rect 141234 372444 141240 372456
rect 141292 372444 141298 372496
rect 141234 371832 141240 371884
rect 141292 371872 141298 371884
rect 142062 371872 142068 371884
rect 141292 371844 142068 371872
rect 141292 371832 141298 371844
rect 142062 371832 142068 371844
rect 142120 371872 142126 371884
rect 178770 371872 178776 371884
rect 142120 371844 178776 371872
rect 142120 371832 142126 371844
rect 178770 371832 178776 371844
rect 178828 371872 178834 371884
rect 182818 371872 182824 371884
rect 178828 371844 182824 371872
rect 178828 371832 178834 371844
rect 182818 371832 182824 371844
rect 182876 371832 182882 371884
rect 187050 371832 187056 371884
rect 187108 371872 187114 371884
rect 209038 371872 209044 371884
rect 187108 371844 209044 371872
rect 187108 371832 187114 371844
rect 209038 371832 209044 371844
rect 209096 371832 209102 371884
rect 234522 371832 234528 371884
rect 234580 371872 234586 371884
rect 298094 371872 298100 371884
rect 234580 371844 298100 371872
rect 234580 371832 234586 371844
rect 298094 371832 298100 371844
rect 298152 371832 298158 371884
rect 169754 371220 169760 371272
rect 169812 371260 169818 371272
rect 170398 371260 170404 371272
rect 169812 371232 170404 371260
rect 169812 371220 169818 371232
rect 170398 371220 170404 371232
rect 170456 371220 170462 371272
rect 67818 371152 67824 371204
rect 67876 371192 67882 371204
rect 158070 371192 158076 371204
rect 67876 371164 158076 371192
rect 67876 371152 67882 371164
rect 158070 371152 158076 371164
rect 158128 371152 158134 371204
rect 161382 371152 161388 371204
rect 161440 371192 161446 371204
rect 231210 371192 231216 371204
rect 161440 371164 231216 371192
rect 161440 371152 161446 371164
rect 231210 371152 231216 371164
rect 231268 371152 231274 371204
rect 150342 371084 150348 371136
rect 150400 371124 150406 371136
rect 218054 371124 218060 371136
rect 150400 371096 218060 371124
rect 150400 371084 150406 371096
rect 218054 371084 218060 371096
rect 218112 371084 218118 371136
rect 232498 370472 232504 370524
rect 232556 370512 232562 370524
rect 265250 370512 265256 370524
rect 232556 370484 265256 370512
rect 232556 370472 232562 370484
rect 265250 370472 265256 370484
rect 265308 370472 265314 370524
rect 101950 369792 101956 369844
rect 102008 369832 102014 369844
rect 236638 369832 236644 369844
rect 102008 369804 236644 369832
rect 102008 369792 102014 369804
rect 236638 369792 236644 369804
rect 236696 369792 236702 369844
rect 110414 369724 110420 369776
rect 110472 369764 110478 369776
rect 111058 369764 111064 369776
rect 110472 369736 111064 369764
rect 110472 369724 110478 369736
rect 111058 369724 111064 369736
rect 111116 369764 111122 369776
rect 148962 369764 148968 369776
rect 111116 369736 148968 369764
rect 111116 369724 111122 369736
rect 148962 369724 148968 369736
rect 149020 369724 149026 369776
rect 151170 369724 151176 369776
rect 151228 369764 151234 369776
rect 255406 369764 255412 369776
rect 151228 369736 255412 369764
rect 151228 369724 151234 369736
rect 255406 369724 255412 369736
rect 255464 369724 255470 369776
rect 114462 368432 114468 368484
rect 114520 368472 114526 368484
rect 281810 368472 281816 368484
rect 114520 368444 281816 368472
rect 114520 368432 114526 368444
rect 281810 368432 281816 368444
rect 281868 368432 281874 368484
rect 69106 368364 69112 368416
rect 69164 368404 69170 368416
rect 165706 368404 165712 368416
rect 69164 368376 165712 368404
rect 69164 368364 69170 368376
rect 165706 368364 165712 368376
rect 165764 368404 165770 368416
rect 166350 368404 166356 368416
rect 165764 368376 166356 368404
rect 165764 368364 165770 368376
rect 166350 368364 166356 368376
rect 166408 368364 166414 368416
rect 168282 368364 168288 368416
rect 168340 368404 168346 368416
rect 227714 368404 227720 368416
rect 168340 368376 227720 368404
rect 168340 368364 168346 368376
rect 227714 368364 227720 368376
rect 227772 368404 227778 368416
rect 228542 368404 228548 368416
rect 227772 368376 228548 368404
rect 227772 368364 227778 368376
rect 228542 368364 228548 368376
rect 228600 368364 228606 368416
rect 98362 367752 98368 367804
rect 98420 367792 98426 367804
rect 113358 367792 113364 367804
rect 98420 367764 113364 367792
rect 98420 367752 98426 367764
rect 113358 367752 113364 367764
rect 113416 367792 113422 367804
rect 114462 367792 114468 367804
rect 113416 367764 114468 367792
rect 113416 367752 113422 367764
rect 114462 367752 114468 367764
rect 114520 367752 114526 367804
rect 228358 367752 228364 367804
rect 228416 367792 228422 367804
rect 288434 367792 288440 367804
rect 228416 367764 288440 367792
rect 228416 367752 228422 367764
rect 288434 367752 288440 367764
rect 288492 367752 288498 367804
rect 67726 367004 67732 367056
rect 67784 367044 67790 367056
rect 180794 367044 180800 367056
rect 67784 367016 180800 367044
rect 67784 367004 67790 367016
rect 180794 367004 180800 367016
rect 180852 367044 180858 367056
rect 181530 367044 181536 367056
rect 180852 367016 181536 367044
rect 180852 367004 180858 367016
rect 181530 367004 181536 367016
rect 181588 367004 181594 367056
rect 97258 366936 97264 366988
rect 97316 366976 97322 366988
rect 161474 366976 161480 366988
rect 97316 366948 161480 366976
rect 97316 366936 97322 366948
rect 161474 366936 161480 366948
rect 161532 366976 161538 366988
rect 162210 366976 162216 366988
rect 161532 366948 162216 366976
rect 161532 366936 161538 366948
rect 162210 366936 162216 366948
rect 162268 366936 162274 366988
rect 183370 366324 183376 366376
rect 183428 366364 183434 366376
rect 190546 366364 190552 366376
rect 183428 366336 190552 366364
rect 183428 366324 183434 366336
rect 190546 366324 190552 366336
rect 190604 366324 190610 366376
rect 218698 366324 218704 366376
rect 218756 366364 218762 366376
rect 263594 366364 263600 366376
rect 218756 366336 263600 366364
rect 218756 366324 218762 366336
rect 263594 366324 263600 366336
rect 263652 366324 263658 366376
rect 93118 365644 93124 365696
rect 93176 365684 93182 365696
rect 171226 365684 171232 365696
rect 93176 365656 171232 365684
rect 93176 365644 93182 365656
rect 171226 365644 171232 365656
rect 171284 365684 171290 365696
rect 171870 365684 171876 365696
rect 171284 365656 171876 365684
rect 171284 365644 171290 365656
rect 171870 365644 171876 365656
rect 171928 365644 171934 365696
rect 163866 365576 163872 365628
rect 163924 365616 163930 365628
rect 221458 365616 221464 365628
rect 163924 365588 221464 365616
rect 163924 365576 163930 365588
rect 221458 365576 221464 365588
rect 221516 365576 221522 365628
rect 249702 365100 249708 365152
rect 249760 365140 249766 365152
rect 252554 365140 252560 365152
rect 249760 365112 252560 365140
rect 249760 365100 249766 365112
rect 252554 365100 252560 365112
rect 252612 365100 252618 365152
rect 211798 364964 211804 365016
rect 211856 365004 211862 365016
rect 256786 365004 256792 365016
rect 211856 364976 256792 365004
rect 211856 364964 211862 364976
rect 256786 364964 256792 364976
rect 256844 364964 256850 365016
rect 241514 364392 241520 364404
rect 241486 364352 241520 364392
rect 241572 364392 241578 364404
rect 249058 364392 249064 364404
rect 241572 364364 249064 364392
rect 241572 364352 241578 364364
rect 249058 364352 249064 364364
rect 249116 364352 249122 364404
rect 104710 364284 104716 364336
rect 104768 364324 104774 364336
rect 241486 364324 241514 364352
rect 104768 364296 241514 364324
rect 104768 364284 104774 364296
rect 60550 364216 60556 364268
rect 60608 364256 60614 364268
rect 142982 364256 142988 364268
rect 60608 364228 142988 364256
rect 60608 364216 60614 364228
rect 142982 364216 142988 364228
rect 143040 364216 143046 364268
rect 153010 364216 153016 364268
rect 153068 364256 153074 364268
rect 272150 364256 272156 364268
rect 153068 364228 272156 364256
rect 153068 364216 153074 364228
rect 272150 364216 272156 364228
rect 272208 364216 272214 364268
rect 123478 362856 123484 362908
rect 123536 362896 123542 362908
rect 226334 362896 226340 362908
rect 123536 362868 226340 362896
rect 123536 362856 123542 362868
rect 226334 362856 226340 362868
rect 226392 362856 226398 362908
rect 240134 362244 240140 362296
rect 240192 362284 240198 362296
rect 263594 362284 263600 362296
rect 240192 362256 263600 362284
rect 240192 362244 240198 362256
rect 263594 362244 263600 362256
rect 263652 362244 263658 362296
rect 93854 362176 93860 362228
rect 93912 362216 93918 362228
rect 103514 362216 103520 362228
rect 93912 362188 103520 362216
rect 93912 362176 93918 362188
rect 103514 362176 103520 362188
rect 103572 362176 103578 362228
rect 212810 362176 212816 362228
rect 212868 362216 212874 362228
rect 247770 362216 247776 362228
rect 212868 362188 247776 362216
rect 212868 362176 212874 362188
rect 247770 362176 247776 362188
rect 247828 362176 247834 362228
rect 226334 361564 226340 361616
rect 226392 361604 226398 361616
rect 226978 361604 226984 361616
rect 226392 361576 226984 361604
rect 226392 361564 226398 361576
rect 226978 361564 226984 361576
rect 227036 361564 227042 361616
rect 155218 361496 155224 361548
rect 155276 361536 155282 361548
rect 249150 361536 249156 361548
rect 155276 361508 249156 361536
rect 155276 361496 155282 361508
rect 249150 361496 249156 361508
rect 249208 361536 249214 361548
rect 249610 361536 249616 361548
rect 249208 361508 249616 361536
rect 249208 361496 249214 361508
rect 249610 361496 249616 361508
rect 249668 361496 249674 361548
rect 74626 361428 74632 361480
rect 74684 361468 74690 361480
rect 156690 361468 156696 361480
rect 74684 361440 156696 361468
rect 74684 361428 74690 361440
rect 156690 361428 156696 361440
rect 156748 361428 156754 361480
rect 231210 360816 231216 360868
rect 231268 360856 231274 360868
rect 253198 360856 253204 360868
rect 231268 360828 253204 360856
rect 231268 360816 231274 360828
rect 253198 360816 253204 360828
rect 253256 360816 253262 360868
rect 156046 360612 156052 360664
rect 156104 360652 156110 360664
rect 156690 360652 156696 360664
rect 156104 360624 156696 360652
rect 156104 360612 156110 360624
rect 156690 360612 156696 360624
rect 156748 360612 156754 360664
rect 141602 360136 141608 360188
rect 141660 360176 141666 360188
rect 255498 360176 255504 360188
rect 141660 360148 255504 360176
rect 141660 360136 141666 360148
rect 255498 360136 255504 360148
rect 255556 360136 255562 360188
rect 84102 360068 84108 360120
rect 84160 360108 84166 360120
rect 155862 360108 155868 360120
rect 84160 360080 155868 360108
rect 84160 360068 84166 360080
rect 155862 360068 155868 360080
rect 155920 360108 155926 360120
rect 179506 360108 179512 360120
rect 155920 360080 179512 360108
rect 155920 360068 155926 360080
rect 179506 360068 179512 360080
rect 179564 360068 179570 360120
rect 179506 359660 179512 359712
rect 179564 359700 179570 359712
rect 180150 359700 180156 359712
rect 179564 359672 180156 359700
rect 179564 359660 179570 359672
rect 180150 359660 180156 359672
rect 180208 359660 180214 359712
rect 255498 359660 255504 359712
rect 255556 359700 255562 359712
rect 255958 359700 255964 359712
rect 255556 359672 255964 359700
rect 255556 359660 255562 359672
rect 255958 359660 255964 359672
rect 256016 359660 256022 359712
rect 195974 359456 195980 359508
rect 196032 359496 196038 359508
rect 240134 359496 240140 359508
rect 196032 359468 240140 359496
rect 196032 359456 196038 359468
rect 240134 359456 240140 359468
rect 240192 359456 240198 359508
rect 69014 358708 69020 358760
rect 69072 358748 69078 358760
rect 69658 358748 69664 358760
rect 69072 358720 69664 358748
rect 69072 358708 69078 358720
rect 69658 358708 69664 358720
rect 69716 358748 69722 358760
rect 69716 358720 74534 358748
rect 69716 358708 69722 358720
rect 74506 358680 74534 358720
rect 142798 358708 142804 358760
rect 142856 358748 142862 358760
rect 285858 358748 285864 358760
rect 142856 358720 285864 358748
rect 142856 358708 142862 358720
rect 285858 358708 285864 358720
rect 285916 358708 285922 358760
rect 194594 358680 194600 358692
rect 74506 358652 194600 358680
rect 194594 358640 194600 358652
rect 194652 358640 194658 358692
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4798 358476 4804 358488
rect 2832 358448 4804 358476
rect 2832 358436 2838 358448
rect 4798 358436 4804 358448
rect 4856 358436 4862 358488
rect 247770 358028 247776 358080
rect 247828 358068 247834 358080
rect 253934 358068 253940 358080
rect 247828 358040 253940 358068
rect 247828 358028 247834 358040
rect 253934 358028 253940 358040
rect 253992 358028 253998 358080
rect 103422 356668 103428 356720
rect 103480 356708 103486 356720
rect 110414 356708 110420 356720
rect 103480 356680 110420 356708
rect 103480 356668 103486 356680
rect 110414 356668 110420 356680
rect 110472 356668 110478 356720
rect 126238 356668 126244 356720
rect 126296 356708 126302 356720
rect 155862 356708 155868 356720
rect 126296 356680 155868 356708
rect 126296 356668 126302 356680
rect 155862 356668 155868 356680
rect 155920 356708 155926 356720
rect 212810 356708 212816 356720
rect 155920 356680 212816 356708
rect 155920 356668 155926 356680
rect 212810 356668 212816 356680
rect 212868 356668 212874 356720
rect 242158 356668 242164 356720
rect 242216 356708 242222 356720
rect 292574 356708 292580 356720
rect 242216 356680 292580 356708
rect 242216 356668 242222 356680
rect 292574 356668 292580 356680
rect 292632 356668 292638 356720
rect 110414 356056 110420 356108
rect 110472 356096 110478 356108
rect 239398 356096 239404 356108
rect 110472 356068 239404 356096
rect 110472 356056 110478 356068
rect 239398 356056 239404 356068
rect 239456 356056 239462 356108
rect 75914 355988 75920 356040
rect 75972 356028 75978 356040
rect 76558 356028 76564 356040
rect 75972 356000 76564 356028
rect 75972 355988 75978 356000
rect 76558 355988 76564 356000
rect 76616 356028 76622 356040
rect 202966 356028 202972 356040
rect 76616 356000 202972 356028
rect 76616 355988 76622 356000
rect 202966 355988 202972 356000
rect 203024 355988 203030 356040
rect 102226 355920 102232 355972
rect 102284 355960 102290 355972
rect 103422 355960 103428 355972
rect 102284 355932 103428 355960
rect 102284 355920 102290 355932
rect 103422 355920 103428 355932
rect 103480 355960 103486 355972
rect 218790 355960 218796 355972
rect 103480 355932 218796 355960
rect 103480 355920 103486 355932
rect 218790 355920 218796 355932
rect 218848 355920 218854 355972
rect 222838 355308 222844 355360
rect 222896 355348 222902 355360
rect 244918 355348 244924 355360
rect 222896 355320 244924 355348
rect 222896 355308 222902 355320
rect 244918 355308 244924 355320
rect 244976 355308 244982 355360
rect 249610 355308 249616 355360
rect 249668 355348 249674 355360
rect 260374 355348 260380 355360
rect 249668 355320 260380 355348
rect 249668 355308 249674 355320
rect 260374 355308 260380 355320
rect 260432 355308 260438 355360
rect 137278 354628 137284 354680
rect 137336 354668 137342 354680
rect 205634 354668 205640 354680
rect 137336 354640 205640 354668
rect 137336 354628 137342 354640
rect 205634 354628 205640 354640
rect 205692 354628 205698 354680
rect 100754 353948 100760 354000
rect 100812 353988 100818 354000
rect 118786 353988 118792 354000
rect 100812 353960 118792 353988
rect 100812 353948 100818 353960
rect 118786 353948 118792 353960
rect 118844 353948 118850 354000
rect 236638 353948 236644 354000
rect 236696 353988 236702 354000
rect 262398 353988 262404 354000
rect 236696 353960 262404 353988
rect 236696 353948 236702 353960
rect 262398 353948 262404 353960
rect 262456 353948 262462 354000
rect 118786 353268 118792 353320
rect 118844 353308 118850 353320
rect 238110 353308 238116 353320
rect 118844 353280 238116 353308
rect 118844 353268 118850 353280
rect 238110 353268 238116 353280
rect 238168 353268 238174 353320
rect 74534 353200 74540 353252
rect 74592 353240 74598 353252
rect 184290 353240 184296 353252
rect 74592 353212 184296 353240
rect 74592 353200 74598 353212
rect 184290 353200 184296 353212
rect 184348 353200 184354 353252
rect 205634 352588 205640 352640
rect 205692 352628 205698 352640
rect 252830 352628 252836 352640
rect 205692 352600 252836 352628
rect 205692 352588 205698 352600
rect 252830 352588 252836 352600
rect 252888 352588 252894 352640
rect 108942 352520 108948 352572
rect 109000 352560 109006 352572
rect 280338 352560 280344 352572
rect 109000 352532 280344 352560
rect 109000 352520 109006 352532
rect 280338 352520 280344 352532
rect 280396 352520 280402 352572
rect 119982 351840 119988 351892
rect 120040 351880 120046 351892
rect 274818 351880 274824 351892
rect 120040 351852 274824 351880
rect 120040 351840 120046 351852
rect 274818 351840 274824 351852
rect 274876 351840 274882 351892
rect 172330 351160 172336 351212
rect 172388 351200 172394 351212
rect 181438 351200 181444 351212
rect 172388 351172 181444 351200
rect 172388 351160 172394 351172
rect 181438 351160 181444 351172
rect 181496 351160 181502 351212
rect 204990 351160 204996 351212
rect 205048 351200 205054 351212
rect 222930 351200 222936 351212
rect 205048 351172 222936 351200
rect 205048 351160 205054 351172
rect 222930 351160 222936 351172
rect 222988 351160 222994 351212
rect 180702 349868 180708 349920
rect 180760 349908 180766 349920
rect 254578 349908 254584 349920
rect 180760 349880 254584 349908
rect 180760 349868 180766 349880
rect 254578 349868 254584 349880
rect 254636 349868 254642 349920
rect 107562 349800 107568 349852
rect 107620 349840 107626 349852
rect 278866 349840 278872 349852
rect 107620 349812 278872 349840
rect 107620 349800 107626 349812
rect 278866 349800 278872 349812
rect 278924 349800 278930 349852
rect 130378 349052 130384 349104
rect 130436 349092 130442 349104
rect 130654 349092 130660 349104
rect 130436 349064 130660 349092
rect 130436 349052 130442 349064
rect 130654 349052 130660 349064
rect 130712 349092 130718 349104
rect 231118 349092 231124 349104
rect 130712 349064 231124 349092
rect 130712 349052 130718 349064
rect 231118 349052 231124 349064
rect 231176 349052 231182 349104
rect 188982 348372 188988 348424
rect 189040 348412 189046 348424
rect 253474 348412 253480 348424
rect 189040 348384 253480 348412
rect 189040 348372 189046 348384
rect 253474 348372 253480 348384
rect 253532 348372 253538 348424
rect 259362 347692 259368 347744
rect 259420 347732 259426 347744
rect 261110 347732 261116 347744
rect 259420 347704 261116 347732
rect 259420 347692 259426 347704
rect 261110 347692 261116 347704
rect 261168 347692 261174 347744
rect 216030 347080 216036 347132
rect 216088 347120 216094 347132
rect 261202 347120 261208 347132
rect 216088 347092 261208 347120
rect 216088 347080 216094 347092
rect 261202 347080 261208 347092
rect 261260 347080 261266 347132
rect 180150 347012 180156 347064
rect 180208 347052 180214 347064
rect 242342 347052 242348 347064
rect 180208 347024 242348 347052
rect 180208 347012 180214 347024
rect 242342 347012 242348 347024
rect 242400 347012 242406 347064
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 42702 346372 42708 346384
rect 3200 346344 42708 346372
rect 3200 346332 3206 346344
rect 42702 346332 42708 346344
rect 42760 346332 42766 346384
rect 42702 345856 42708 345908
rect 42760 345896 42766 345908
rect 43438 345896 43444 345908
rect 42760 345868 43444 345896
rect 42760 345856 42766 345868
rect 43438 345856 43444 345868
rect 43496 345856 43502 345908
rect 72510 345720 72516 345772
rect 72568 345760 72574 345772
rect 73062 345760 73068 345772
rect 72568 345732 73068 345760
rect 72568 345720 72574 345732
rect 73062 345720 73068 345732
rect 73120 345720 73126 345772
rect 175550 345108 175556 345160
rect 175608 345148 175614 345160
rect 198734 345148 198740 345160
rect 175608 345120 198740 345148
rect 175608 345108 175614 345120
rect 198734 345108 198740 345120
rect 198792 345108 198798 345160
rect 72510 345040 72516 345092
rect 72568 345080 72574 345092
rect 231118 345080 231124 345092
rect 72568 345052 231124 345080
rect 72568 345040 72574 345052
rect 231118 345040 231124 345052
rect 231176 345040 231182 345092
rect 247678 344292 247684 344344
rect 247736 344332 247742 344344
rect 251910 344332 251916 344344
rect 247736 344304 251916 344332
rect 247736 344292 247742 344304
rect 251910 344292 251916 344304
rect 251968 344292 251974 344344
rect 130378 343680 130384 343732
rect 130436 343720 130442 343732
rect 228450 343720 228456 343732
rect 130436 343692 228456 343720
rect 130436 343680 130442 343692
rect 228450 343680 228456 343692
rect 228508 343680 228514 343732
rect 129090 343612 129096 343664
rect 129148 343652 129154 343664
rect 129642 343652 129648 343664
rect 129148 343624 129648 343652
rect 129148 343612 129154 343624
rect 129642 343612 129648 343624
rect 129700 343652 129706 343664
rect 246482 343652 246488 343664
rect 129700 343624 246488 343652
rect 129700 343612 129706 343624
rect 246482 343612 246488 343624
rect 246540 343612 246546 343664
rect 209130 342864 209136 342916
rect 209188 342904 209194 342916
rect 277394 342904 277400 342916
rect 209188 342876 277400 342904
rect 209188 342864 209194 342876
rect 277394 342864 277400 342876
rect 277452 342864 277458 342916
rect 175090 342320 175096 342372
rect 175148 342360 175154 342372
rect 202138 342360 202144 342372
rect 175148 342332 202144 342360
rect 175148 342320 175154 342332
rect 202138 342320 202144 342332
rect 202196 342320 202202 342372
rect 95142 342252 95148 342304
rect 95200 342292 95206 342304
rect 294046 342292 294052 342304
rect 95200 342264 294052 342292
rect 95200 342252 95206 342264
rect 294046 342252 294052 342264
rect 294104 342252 294110 342304
rect 143442 341572 143448 341624
rect 143500 341612 143506 341624
rect 155402 341612 155408 341624
rect 143500 341584 155408 341612
rect 143500 341572 143506 341584
rect 155402 341572 155408 341584
rect 155460 341572 155466 341624
rect 177942 341572 177948 341624
rect 178000 341612 178006 341624
rect 253290 341612 253296 341624
rect 178000 341584 253296 341612
rect 178000 341572 178006 341584
rect 253290 341572 253296 341584
rect 253348 341572 253354 341624
rect 101398 341504 101404 341556
rect 101456 341544 101462 341556
rect 268010 341544 268016 341556
rect 101456 341516 268016 341544
rect 101456 341504 101462 341516
rect 268010 341504 268016 341516
rect 268068 341504 268074 341556
rect 183186 340144 183192 340196
rect 183244 340184 183250 340196
rect 246390 340184 246396 340196
rect 183244 340156 246396 340184
rect 183244 340144 183250 340156
rect 246390 340144 246396 340156
rect 246448 340144 246454 340196
rect 67542 339464 67548 339516
rect 67600 339504 67606 339516
rect 291470 339504 291476 339516
rect 67600 339476 291476 339504
rect 67600 339464 67606 339476
rect 291470 339464 291476 339476
rect 291528 339464 291534 339516
rect 239398 339396 239404 339448
rect 239456 339436 239462 339448
rect 246298 339436 246304 339448
rect 239456 339408 246304 339436
rect 239456 339396 239462 339408
rect 246298 339396 246304 339408
rect 246356 339396 246362 339448
rect 215938 338784 215944 338836
rect 215996 338824 216002 338836
rect 243538 338824 243544 338836
rect 215996 338796 243544 338824
rect 215996 338784 216002 338796
rect 243538 338784 243544 338796
rect 243596 338784 243602 338836
rect 33134 338716 33140 338768
rect 33192 338756 33198 338768
rect 175090 338756 175096 338768
rect 33192 338728 175096 338756
rect 33192 338716 33198 338728
rect 175090 338716 175096 338728
rect 175148 338716 175154 338768
rect 191742 338716 191748 338768
rect 191800 338756 191806 338768
rect 222194 338756 222200 338768
rect 191800 338728 222200 338756
rect 191800 338716 191806 338728
rect 222194 338716 222200 338728
rect 222252 338716 222258 338768
rect 246942 338716 246948 338768
rect 247000 338756 247006 338768
rect 258074 338756 258080 338768
rect 247000 338728 258080 338756
rect 247000 338716 247006 338728
rect 258074 338716 258080 338728
rect 258132 338716 258138 338768
rect 148870 338104 148876 338156
rect 148928 338144 148934 338156
rect 150434 338144 150440 338156
rect 148928 338116 150440 338144
rect 148928 338104 148934 338116
rect 150434 338104 150440 338116
rect 150492 338144 150498 338156
rect 215294 338144 215300 338156
rect 150492 338116 215300 338144
rect 150492 338104 150498 338116
rect 215294 338104 215300 338116
rect 215352 338104 215358 338156
rect 142798 337356 142804 337408
rect 142856 337396 142862 337408
rect 188890 337396 188896 337408
rect 142856 337368 188896 337396
rect 142856 337356 142862 337368
rect 188890 337356 188896 337368
rect 188948 337396 188954 337408
rect 215570 337396 215576 337408
rect 188948 337368 215576 337396
rect 188948 337356 188954 337368
rect 215570 337356 215576 337368
rect 215628 337356 215634 337408
rect 221458 337356 221464 337408
rect 221516 337396 221522 337408
rect 274634 337396 274640 337408
rect 221516 337368 274640 337396
rect 221516 337356 221522 337368
rect 274634 337356 274640 337368
rect 274692 337356 274698 337408
rect 141602 336744 141608 336796
rect 141660 336784 141666 336796
rect 247770 336784 247776 336796
rect 141660 336756 247776 336784
rect 141660 336744 141666 336756
rect 247770 336744 247776 336756
rect 247828 336744 247834 336796
rect 165522 335996 165528 336048
rect 165580 336036 165586 336048
rect 215478 336036 215484 336048
rect 165580 336008 215484 336036
rect 165580 335996 165586 336008
rect 215478 335996 215484 336008
rect 215536 335996 215542 336048
rect 244274 335792 244280 335844
rect 244332 335832 244338 335844
rect 245010 335832 245016 335844
rect 244332 335804 245016 335832
rect 244332 335792 244338 335804
rect 245010 335792 245016 335804
rect 245068 335792 245074 335844
rect 143074 335316 143080 335368
rect 143132 335356 143138 335368
rect 244274 335356 244280 335368
rect 143132 335328 244280 335356
rect 143132 335316 143138 335328
rect 244274 335316 244280 335328
rect 244332 335316 244338 335368
rect 222286 334636 222292 334688
rect 222344 334676 222350 334688
rect 260834 334676 260840 334688
rect 222344 334648 260840 334676
rect 222344 334636 222350 334648
rect 260834 334636 260840 334648
rect 260892 334636 260898 334688
rect 151630 334568 151636 334620
rect 151688 334608 151694 334620
rect 160186 334608 160192 334620
rect 151688 334580 160192 334608
rect 151688 334568 151694 334580
rect 160186 334568 160192 334580
rect 160244 334568 160250 334620
rect 177390 334568 177396 334620
rect 177448 334608 177454 334620
rect 187510 334608 187516 334620
rect 177448 334580 187516 334608
rect 177448 334568 177454 334580
rect 187510 334568 187516 334580
rect 187568 334608 187574 334620
rect 242894 334608 242900 334620
rect 187568 334580 242900 334608
rect 187568 334568 187574 334580
rect 242894 334568 242900 334580
rect 242952 334568 242958 334620
rect 160186 333956 160192 334008
rect 160244 333996 160250 334008
rect 160738 333996 160744 334008
rect 160244 333968 160744 333996
rect 160244 333956 160250 333968
rect 160738 333956 160744 333968
rect 160796 333996 160802 334008
rect 205634 333996 205640 334008
rect 160796 333968 205640 333996
rect 160796 333956 160802 333968
rect 205634 333956 205640 333968
rect 205692 333956 205698 334008
rect 205634 333276 205640 333328
rect 205692 333316 205698 333328
rect 245746 333316 245752 333328
rect 205692 333288 245752 333316
rect 205692 333276 205698 333288
rect 245746 333276 245752 333288
rect 245804 333276 245810 333328
rect 246482 333276 246488 333328
rect 246540 333316 246546 333328
rect 273530 333316 273536 333328
rect 246540 333288 273536 333316
rect 246540 333276 246546 333288
rect 273530 333276 273536 333288
rect 273588 333276 273594 333328
rect 30374 333208 30380 333260
rect 30432 333248 30438 333260
rect 154022 333248 154028 333260
rect 30432 333220 154028 333248
rect 30432 333208 30438 333220
rect 154022 333208 154028 333220
rect 154080 333208 154086 333260
rect 172422 333208 172428 333260
rect 172480 333248 172486 333260
rect 190362 333248 190368 333260
rect 172480 333220 190368 333248
rect 172480 333208 172486 333220
rect 190362 333208 190368 333220
rect 190420 333248 190426 333260
rect 247034 333248 247040 333260
rect 190420 333220 247040 333248
rect 190420 333208 190426 333220
rect 247034 333208 247040 333220
rect 247092 333208 247098 333260
rect 234614 332528 234620 332580
rect 234672 332568 234678 332580
rect 240778 332568 240784 332580
rect 234672 332540 240784 332568
rect 234672 332528 234678 332540
rect 240778 332528 240784 332540
rect 240836 332528 240842 332580
rect 158070 331848 158076 331900
rect 158128 331888 158134 331900
rect 173710 331888 173716 331900
rect 158128 331860 173716 331888
rect 158128 331848 158134 331860
rect 173710 331848 173716 331860
rect 173768 331888 173774 331900
rect 243170 331888 243176 331900
rect 173768 331860 243176 331888
rect 173768 331848 173774 331860
rect 243170 331848 243176 331860
rect 243228 331848 243234 331900
rect 148502 331236 148508 331288
rect 148560 331276 148566 331288
rect 234614 331276 234620 331288
rect 148560 331248 234620 331276
rect 148560 331236 148566 331248
rect 234614 331236 234620 331248
rect 234672 331236 234678 331288
rect 94498 330488 94504 330540
rect 94556 330528 94562 330540
rect 153194 330528 153200 330540
rect 94556 330500 153200 330528
rect 94556 330488 94562 330500
rect 153194 330488 153200 330500
rect 153252 330488 153258 330540
rect 172238 329876 172244 329928
rect 172296 329916 172302 329928
rect 201586 329916 201592 329928
rect 172296 329888 201592 329916
rect 172296 329876 172302 329888
rect 201586 329876 201592 329888
rect 201644 329876 201650 329928
rect 166258 329808 166264 329860
rect 166316 329848 166322 329860
rect 233878 329848 233884 329860
rect 166316 329820 233884 329848
rect 166316 329808 166322 329820
rect 233878 329808 233884 329820
rect 233936 329808 233942 329860
rect 252370 329740 252376 329792
rect 252428 329780 252434 329792
rect 254026 329780 254032 329792
rect 252428 329752 254032 329780
rect 252428 329740 252434 329752
rect 254026 329740 254032 329752
rect 254084 329740 254090 329792
rect 164878 328516 164884 328568
rect 164936 328556 164942 328568
rect 240134 328556 240140 328568
rect 164936 328528 240140 328556
rect 164936 328516 164942 328528
rect 240134 328516 240140 328528
rect 240192 328516 240198 328568
rect 116670 328448 116676 328500
rect 116728 328488 116734 328500
rect 252370 328488 252376 328500
rect 116728 328460 252376 328488
rect 116728 328448 116734 328460
rect 252370 328448 252376 328460
rect 252428 328448 252434 328500
rect 218146 328380 218152 328432
rect 218204 328420 218210 328432
rect 218698 328420 218704 328432
rect 218204 328392 218704 328420
rect 218204 328380 218210 328392
rect 218698 328380 218704 328392
rect 218756 328380 218762 328432
rect 260374 328380 260380 328432
rect 260432 328420 260438 328432
rect 266722 328420 266728 328432
rect 260432 328392 266728 328420
rect 260432 328380 260438 328392
rect 266722 328380 266728 328392
rect 266780 328380 266786 328432
rect 209774 327700 209780 327752
rect 209832 327740 209838 327752
rect 266354 327740 266360 327752
rect 209832 327712 266360 327740
rect 209832 327700 209838 327712
rect 266354 327700 266360 327712
rect 266412 327700 266418 327752
rect 190362 327156 190368 327208
rect 190420 327196 190426 327208
rect 192478 327196 192484 327208
rect 190420 327168 192484 327196
rect 190420 327156 190426 327168
rect 192478 327156 192484 327168
rect 192536 327156 192542 327208
rect 121454 327088 121460 327140
rect 121512 327128 121518 327140
rect 218146 327128 218152 327140
rect 121512 327100 218152 327128
rect 121512 327088 121518 327100
rect 218146 327088 218152 327100
rect 218204 327088 218210 327140
rect 123570 326340 123576 326392
rect 123628 326380 123634 326392
rect 154482 326380 154488 326392
rect 123628 326352 154488 326380
rect 123628 326340 123634 326352
rect 154482 326340 154488 326352
rect 154540 326340 154546 326392
rect 160922 326340 160928 326392
rect 160980 326380 160986 326392
rect 169386 326380 169392 326392
rect 160980 326352 169392 326380
rect 160980 326340 160986 326352
rect 169386 326340 169392 326352
rect 169444 326380 169450 326392
rect 241514 326380 241520 326392
rect 169444 326352 241520 326380
rect 169444 326340 169450 326352
rect 241514 326340 241520 326352
rect 241572 326340 241578 326392
rect 242250 326340 242256 326392
rect 242308 326380 242314 326392
rect 256694 326380 256700 326392
rect 242308 326352 256700 326380
rect 242308 326340 242314 326352
rect 256694 326340 256700 326352
rect 256752 326340 256758 326392
rect 96706 325660 96712 325712
rect 96764 325700 96770 325712
rect 250438 325700 250444 325712
rect 96764 325672 250444 325700
rect 96764 325660 96770 325672
rect 250438 325660 250444 325672
rect 250496 325660 250502 325712
rect 232590 324912 232596 324964
rect 232648 324952 232654 324964
rect 271874 324952 271880 324964
rect 232648 324924 271880 324952
rect 232648 324912 232654 324924
rect 271874 324912 271880 324924
rect 271932 324912 271938 324964
rect 138658 324368 138664 324420
rect 138716 324408 138722 324420
rect 209774 324408 209780 324420
rect 138716 324380 209780 324408
rect 138716 324368 138722 324380
rect 209774 324368 209780 324380
rect 209832 324408 209838 324420
rect 210234 324408 210240 324420
rect 209832 324380 210240 324408
rect 209832 324368 209838 324380
rect 210234 324368 210240 324380
rect 210292 324368 210298 324420
rect 41230 324300 41236 324352
rect 41288 324340 41294 324352
rect 154482 324340 154488 324352
rect 41288 324312 154488 324340
rect 41288 324300 41294 324312
rect 154482 324300 154488 324312
rect 154540 324300 154546 324352
rect 175918 324300 175924 324352
rect 175976 324340 175982 324352
rect 176470 324340 176476 324352
rect 175976 324312 176476 324340
rect 175976 324300 175982 324312
rect 176470 324300 176476 324312
rect 176528 324340 176534 324352
rect 258718 324340 258724 324352
rect 176528 324312 258724 324340
rect 176528 324300 176534 324312
rect 258718 324300 258724 324312
rect 258776 324300 258782 324352
rect 260834 323756 260840 323808
rect 260892 323796 260898 323808
rect 261202 323796 261208 323808
rect 260892 323768 261208 323796
rect 260892 323756 260898 323768
rect 261202 323756 261208 323768
rect 261260 323756 261266 323808
rect 151170 323008 151176 323060
rect 151228 323048 151234 323060
rect 260834 323048 260840 323060
rect 151228 323020 260840 323048
rect 151228 323008 151234 323020
rect 260834 323008 260840 323020
rect 260892 323008 260898 323060
rect 155310 322940 155316 322992
rect 155368 322980 155374 322992
rect 269298 322980 269304 322992
rect 155368 322952 269304 322980
rect 155368 322940 155374 322952
rect 269298 322940 269304 322952
rect 269356 322940 269362 322992
rect 35894 322328 35900 322380
rect 35952 322368 35958 322380
rect 153286 322368 153292 322380
rect 35952 322340 153292 322368
rect 35952 322328 35958 322340
rect 153286 322328 153292 322340
rect 153344 322328 153350 322380
rect 157058 322260 157064 322312
rect 157116 322300 157122 322312
rect 233602 322300 233608 322312
rect 157116 322272 233608 322300
rect 157116 322260 157122 322272
rect 233602 322260 233608 322272
rect 233660 322260 233666 322312
rect 104802 322192 104808 322244
rect 104860 322232 104866 322244
rect 277394 322232 277400 322244
rect 104860 322204 277400 322232
rect 104860 322192 104866 322204
rect 277394 322192 277400 322204
rect 277452 322232 277458 322244
rect 277762 322232 277768 322244
rect 277452 322204 277768 322232
rect 277452 322192 277458 322204
rect 277762 322192 277768 322204
rect 277820 322192 277826 322244
rect 153838 321580 153844 321632
rect 153896 321620 153902 321632
rect 157058 321620 157064 321632
rect 153896 321592 157064 321620
rect 153896 321580 153902 321592
rect 157058 321580 157064 321592
rect 157116 321580 157122 321632
rect 154482 320832 154488 320884
rect 154540 320872 154546 320884
rect 292574 320872 292580 320884
rect 154540 320844 292580 320872
rect 154540 320832 154546 320844
rect 292574 320832 292580 320844
rect 292632 320832 292638 320884
rect 185578 320152 185584 320204
rect 185636 320192 185642 320204
rect 259730 320192 259736 320204
rect 185636 320164 259736 320192
rect 185636 320152 185642 320164
rect 259730 320152 259736 320164
rect 259788 320152 259794 320204
rect 84838 320084 84844 320136
rect 84896 320124 84902 320136
rect 85482 320124 85488 320136
rect 84896 320096 85488 320124
rect 84896 320084 84902 320096
rect 85482 320084 85488 320096
rect 85540 320124 85546 320136
rect 150158 320124 150164 320136
rect 85540 320096 150164 320124
rect 85540 320084 85546 320096
rect 150158 320084 150164 320096
rect 150216 320124 150222 320136
rect 247126 320124 247132 320136
rect 150216 320096 247132 320124
rect 150216 320084 150222 320096
rect 247126 320084 247132 320096
rect 247184 320084 247190 320136
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 41230 319444 41236 319456
rect 4120 319416 41236 319444
rect 4120 319404 4126 319416
rect 41230 319404 41236 319416
rect 41288 319404 41294 319456
rect 252278 319404 252284 319456
rect 252336 319444 252342 319456
rect 292666 319444 292672 319456
rect 252336 319416 292672 319444
rect 252336 319404 252342 319416
rect 292666 319404 292672 319416
rect 292724 319404 292730 319456
rect 188430 318792 188436 318844
rect 188488 318832 188494 318844
rect 266630 318832 266636 318844
rect 188488 318804 266636 318832
rect 188488 318792 188494 318804
rect 266630 318792 266636 318804
rect 266688 318792 266694 318844
rect 44266 318044 44272 318096
rect 44324 318084 44330 318096
rect 94498 318084 94504 318096
rect 44324 318056 94504 318084
rect 44324 318044 44330 318056
rect 94498 318044 94504 318056
rect 94556 318044 94562 318096
rect 178678 317500 178684 317552
rect 178736 317540 178742 317552
rect 179322 317540 179328 317552
rect 178736 317512 179328 317540
rect 178736 317500 178742 317512
rect 179322 317500 179328 317512
rect 179380 317540 179386 317552
rect 249150 317540 249156 317552
rect 179380 317512 249156 317540
rect 179380 317500 179386 317512
rect 249150 317500 249156 317512
rect 249208 317500 249214 317552
rect 176010 317432 176016 317484
rect 176068 317472 176074 317484
rect 266538 317472 266544 317484
rect 176068 317444 266544 317472
rect 176068 317432 176074 317444
rect 266538 317432 266544 317444
rect 266596 317432 266602 317484
rect 280246 317364 280252 317416
rect 280304 317404 280310 317416
rect 280430 317404 280436 317416
rect 280304 317376 280436 317404
rect 280304 317364 280310 317376
rect 280430 317364 280436 317376
rect 280488 317364 280494 317416
rect 87598 316752 87604 316804
rect 87656 316792 87662 316804
rect 88242 316792 88248 316804
rect 87656 316764 88248 316792
rect 87656 316752 87662 316764
rect 88242 316752 88248 316764
rect 88300 316752 88306 316804
rect 34422 316684 34428 316736
rect 34480 316724 34486 316736
rect 165430 316724 165436 316736
rect 34480 316696 165436 316724
rect 34480 316684 34486 316696
rect 165430 316684 165436 316696
rect 165488 316724 165494 316736
rect 264974 316724 264980 316736
rect 165488 316696 264980 316724
rect 165488 316684 165494 316696
rect 264974 316684 264980 316696
rect 265032 316684 265038 316736
rect 87598 316004 87604 316056
rect 87656 316044 87662 316056
rect 116578 316044 116584 316056
rect 87656 316016 116584 316044
rect 87656 316004 87662 316016
rect 116578 316004 116584 316016
rect 116636 316004 116642 316056
rect 148870 316004 148876 316056
rect 148928 316044 148934 316056
rect 149790 316044 149796 316056
rect 148928 316016 149796 316044
rect 148928 316004 148934 316016
rect 149790 316004 149796 316016
rect 149848 316004 149854 316056
rect 188338 316004 188344 316056
rect 188396 316044 188402 316056
rect 280430 316044 280436 316056
rect 188396 316016 280436 316044
rect 188396 316004 188402 316016
rect 280430 316004 280436 316016
rect 280488 316004 280494 316056
rect 155402 315460 155408 315512
rect 155460 315500 155466 315512
rect 162210 315500 162216 315512
rect 155460 315472 162216 315500
rect 155460 315460 155466 315472
rect 162210 315460 162216 315472
rect 162268 315460 162274 315512
rect 154022 315324 154028 315376
rect 154080 315364 154086 315376
rect 188430 315364 188436 315376
rect 154080 315336 188436 315364
rect 154080 315324 154086 315336
rect 188430 315324 188436 315336
rect 188488 315324 188494 315376
rect 40034 315256 40040 315308
rect 40092 315296 40098 315308
rect 154114 315296 154120 315308
rect 40092 315268 154120 315296
rect 40092 315256 40098 315268
rect 154114 315256 154120 315268
rect 154172 315256 154178 315308
rect 231118 315256 231124 315308
rect 231176 315296 231182 315308
rect 262858 315296 262864 315308
rect 231176 315268 262864 315296
rect 231176 315256 231182 315268
rect 262858 315256 262864 315268
rect 262916 315256 262922 315308
rect 170582 314712 170588 314764
rect 170640 314752 170646 314764
rect 224218 314752 224224 314764
rect 170640 314724 224224 314752
rect 170640 314712 170646 314724
rect 224218 314712 224224 314724
rect 224276 314712 224282 314764
rect 187786 314644 187792 314696
rect 187844 314684 187850 314696
rect 281534 314684 281540 314696
rect 187844 314656 281540 314684
rect 187844 314644 187850 314656
rect 281534 314644 281540 314656
rect 281592 314684 281598 314696
rect 281810 314684 281816 314696
rect 281592 314656 281816 314684
rect 281592 314644 281598 314656
rect 281810 314644 281816 314656
rect 281868 314644 281874 314696
rect 184198 313352 184204 313404
rect 184256 313392 184262 313404
rect 240778 313392 240784 313404
rect 184256 313364 240784 313392
rect 184256 313352 184262 313364
rect 240778 313352 240784 313364
rect 240836 313352 240842 313404
rect 135990 313284 135996 313336
rect 136048 313324 136054 313336
rect 260926 313324 260932 313336
rect 136048 313296 260932 313324
rect 136048 313284 136054 313296
rect 260926 313284 260932 313296
rect 260984 313284 260990 313336
rect 104158 312604 104164 312656
rect 104216 312644 104222 312656
rect 116026 312644 116032 312656
rect 104216 312616 116032 312644
rect 104216 312604 104222 312616
rect 116026 312604 116032 312616
rect 116084 312644 116090 312656
rect 126882 312644 126888 312656
rect 116084 312616 126888 312644
rect 116084 312604 116090 312616
rect 126882 312604 126888 312616
rect 126940 312604 126946 312656
rect 92474 312536 92480 312588
rect 92532 312576 92538 312588
rect 188338 312576 188344 312588
rect 92532 312548 188344 312576
rect 92532 312536 92538 312548
rect 188338 312536 188344 312548
rect 188396 312536 188402 312588
rect 187694 311924 187700 311976
rect 187752 311964 187758 311976
rect 256878 311964 256884 311976
rect 187752 311936 256884 311964
rect 187752 311924 187758 311936
rect 256878 311924 256884 311936
rect 256936 311924 256942 311976
rect 126330 311856 126336 311908
rect 126388 311896 126394 311908
rect 126882 311896 126888 311908
rect 126388 311868 126888 311896
rect 126388 311856 126394 311868
rect 126882 311856 126888 311868
rect 126940 311896 126946 311908
rect 263870 311896 263876 311908
rect 126940 311868 263876 311896
rect 126940 311856 126946 311868
rect 263870 311856 263876 311868
rect 263928 311856 263934 311908
rect 71038 311176 71044 311228
rect 71096 311216 71102 311228
rect 77478 311216 77484 311228
rect 71096 311188 77484 311216
rect 71096 311176 71102 311188
rect 77478 311176 77484 311188
rect 77536 311176 77542 311228
rect 108206 311176 108212 311228
rect 108264 311216 108270 311228
rect 118694 311216 118700 311228
rect 108264 311188 118700 311216
rect 108264 311176 108270 311188
rect 118694 311176 118700 311188
rect 118752 311216 118758 311228
rect 127618 311216 127624 311228
rect 118752 311188 127624 311216
rect 118752 311176 118758 311188
rect 127618 311176 127624 311188
rect 127676 311176 127682 311228
rect 67726 311108 67732 311160
rect 67784 311148 67790 311160
rect 158714 311148 158720 311160
rect 67784 311120 158720 311148
rect 67784 311108 67790 311120
rect 158714 311108 158720 311120
rect 158772 311148 158778 311160
rect 259546 311148 259552 311160
rect 158772 311120 259552 311148
rect 158772 311108 158778 311120
rect 259546 311108 259552 311120
rect 259604 311108 259610 311160
rect 127618 310496 127624 310548
rect 127676 310536 127682 310548
rect 251910 310536 251916 310548
rect 127676 310508 251916 310536
rect 127676 310496 127682 310508
rect 251910 310496 251916 310508
rect 251968 310496 251974 310548
rect 174722 309748 174728 309800
rect 174780 309788 174786 309800
rect 187694 309788 187700 309800
rect 174780 309760 187700 309788
rect 174780 309748 174786 309760
rect 187694 309748 187700 309760
rect 187752 309748 187758 309800
rect 224862 309748 224868 309800
rect 224920 309788 224926 309800
rect 255314 309788 255320 309800
rect 224920 309760 255320 309788
rect 224920 309748 224926 309760
rect 255314 309748 255320 309760
rect 255372 309748 255378 309800
rect 192478 309544 192484 309596
rect 192536 309584 192542 309596
rect 198826 309584 198832 309596
rect 192536 309556 198832 309584
rect 192536 309544 192542 309556
rect 198826 309544 198832 309556
rect 198884 309584 198890 309596
rect 199378 309584 199384 309596
rect 198884 309556 199384 309584
rect 198884 309544 198890 309556
rect 199378 309544 199384 309556
rect 199436 309544 199442 309596
rect 116578 309136 116584 309188
rect 116636 309176 116642 309188
rect 274910 309176 274916 309188
rect 116636 309148 274916 309176
rect 116636 309136 116642 309148
rect 274910 309136 274916 309148
rect 274968 309136 274974 309188
rect 52270 309068 52276 309120
rect 52328 309108 52334 309120
rect 187694 309108 187700 309120
rect 52328 309080 187700 309108
rect 52328 309068 52334 309080
rect 187694 309068 187700 309080
rect 187752 309068 187758 309120
rect 97258 308388 97264 308440
rect 97316 308428 97322 308440
rect 108206 308428 108212 308440
rect 97316 308400 108212 308428
rect 97316 308388 97322 308400
rect 108206 308388 108212 308400
rect 108264 308388 108270 308440
rect 147582 308388 147588 308440
rect 147640 308428 147646 308440
rect 172514 308428 172520 308440
rect 147640 308400 172520 308428
rect 147640 308388 147646 308400
rect 172514 308388 172520 308400
rect 172572 308388 172578 308440
rect 188890 308388 188896 308440
rect 188948 308428 188954 308440
rect 195238 308428 195244 308440
rect 188948 308400 195244 308428
rect 188948 308388 188954 308400
rect 195238 308388 195244 308400
rect 195296 308388 195302 308440
rect 230474 308388 230480 308440
rect 230532 308428 230538 308440
rect 252738 308428 252744 308440
rect 230532 308400 252744 308428
rect 230532 308388 230538 308400
rect 252738 308388 252744 308400
rect 252796 308388 252802 308440
rect 111794 307776 111800 307828
rect 111852 307816 111858 307828
rect 129090 307816 129096 307828
rect 111852 307788 129096 307816
rect 111852 307776 111858 307788
rect 129090 307776 129096 307788
rect 129148 307776 129154 307828
rect 172514 307776 172520 307828
rect 172572 307816 172578 307828
rect 210050 307816 210056 307828
rect 172572 307788 210056 307816
rect 172572 307776 172578 307788
rect 210050 307776 210056 307788
rect 210108 307776 210114 307828
rect 242802 307776 242808 307828
rect 242860 307816 242866 307828
rect 259454 307816 259460 307828
rect 242860 307788 259460 307816
rect 242860 307776 242866 307788
rect 259454 307776 259460 307788
rect 259512 307776 259518 307828
rect 202138 307708 202144 307760
rect 202196 307748 202202 307760
rect 203978 307748 203984 307760
rect 202196 307720 203984 307748
rect 202196 307708 202202 307720
rect 203978 307708 203984 307720
rect 204036 307708 204042 307760
rect 282914 307708 282920 307760
rect 282972 307748 282978 307760
rect 283098 307748 283104 307760
rect 282972 307720 283104 307748
rect 282972 307708 282978 307720
rect 283098 307708 283104 307720
rect 283156 307708 283162 307760
rect 99190 307096 99196 307148
rect 99248 307136 99254 307148
rect 111794 307136 111800 307148
rect 99248 307108 111800 307136
rect 99248 307096 99254 307108
rect 111794 307096 111800 307108
rect 111852 307096 111858 307148
rect 93118 307028 93124 307080
rect 93176 307068 93182 307080
rect 187786 307068 187792 307080
rect 93176 307040 187792 307068
rect 93176 307028 93182 307040
rect 187786 307028 187792 307040
rect 187844 307028 187850 307080
rect 235902 307028 235908 307080
rect 235960 307068 235966 307080
rect 252554 307068 252560 307080
rect 235960 307040 252560 307068
rect 235960 307028 235966 307040
rect 252554 307028 252560 307040
rect 252612 307028 252618 307080
rect 115198 306416 115204 306468
rect 115256 306456 115262 306468
rect 193858 306456 193864 306468
rect 115256 306428 193864 306456
rect 115256 306416 115262 306428
rect 193858 306416 193864 306428
rect 193916 306416 193922 306468
rect 188062 306348 188068 306400
rect 188120 306388 188126 306400
rect 282914 306388 282920 306400
rect 188120 306360 282920 306388
rect 188120 306348 188126 306360
rect 282914 306348 282920 306360
rect 282972 306348 282978 306400
rect 3418 306280 3424 306332
rect 3476 306320 3482 306332
rect 34422 306320 34428 306332
rect 3476 306292 34428 306320
rect 3476 306280 3482 306292
rect 34422 306280 34428 306292
rect 34480 306280 34486 306332
rect 262858 306144 262864 306196
rect 262916 306184 262922 306196
rect 265066 306184 265072 306196
rect 262916 306156 265072 306184
rect 262916 306144 262922 306156
rect 265066 306144 265072 306156
rect 265124 306144 265130 306196
rect 224218 305668 224224 305720
rect 224276 305708 224282 305720
rect 258074 305708 258080 305720
rect 224276 305680 258080 305708
rect 224276 305668 224282 305680
rect 258074 305668 258080 305680
rect 258132 305668 258138 305720
rect 76282 305600 76288 305652
rect 76340 305640 76346 305652
rect 84838 305640 84844 305652
rect 76340 305612 84844 305640
rect 76340 305600 76346 305612
rect 84838 305600 84844 305612
rect 84896 305600 84902 305652
rect 92382 305600 92388 305652
rect 92440 305640 92446 305652
rect 104158 305640 104164 305652
rect 92440 305612 104164 305640
rect 92440 305600 92446 305612
rect 104158 305600 104164 305612
rect 104216 305600 104222 305652
rect 104710 305600 104716 305652
rect 104768 305640 104774 305652
rect 114646 305640 114652 305652
rect 104768 305612 114652 305640
rect 104768 305600 104774 305612
rect 114646 305600 114652 305612
rect 114704 305600 114710 305652
rect 195422 305600 195428 305652
rect 195480 305640 195486 305652
rect 230382 305640 230388 305652
rect 195480 305612 230388 305640
rect 195480 305600 195486 305612
rect 230382 305600 230388 305612
rect 230440 305600 230446 305652
rect 242434 305600 242440 305652
rect 242492 305640 242498 305652
rect 260098 305640 260104 305652
rect 242492 305612 260104 305640
rect 242492 305600 242498 305612
rect 260098 305600 260104 305612
rect 260156 305640 260162 305652
rect 276290 305640 276296 305652
rect 260156 305612 276296 305640
rect 260156 305600 260162 305612
rect 276290 305600 276296 305612
rect 276348 305600 276354 305652
rect 197354 305192 197360 305244
rect 197412 305232 197418 305244
rect 198366 305232 198372 305244
rect 197412 305204 198372 305232
rect 197412 305192 197418 305204
rect 198366 305192 198372 305204
rect 198424 305192 198430 305244
rect 144730 305056 144736 305108
rect 144788 305096 144794 305108
rect 197354 305096 197360 305108
rect 144788 305068 197360 305096
rect 144788 305056 144794 305068
rect 197354 305056 197360 305068
rect 197412 305056 197418 305108
rect 34422 304988 34428 305040
rect 34480 305028 34486 305040
rect 35158 305028 35164 305040
rect 34480 305000 35164 305028
rect 34480 304988 34486 305000
rect 35158 304988 35164 305000
rect 35216 304988 35222 305040
rect 101490 304988 101496 305040
rect 101548 305028 101554 305040
rect 102042 305028 102048 305040
rect 101548 305000 102048 305028
rect 101548 304988 101554 305000
rect 102042 304988 102048 305000
rect 102100 305028 102106 305040
rect 186314 305028 186320 305040
rect 102100 305000 186320 305028
rect 102100 304988 102106 305000
rect 186314 304988 186320 305000
rect 186372 304988 186378 305040
rect 187510 304988 187516 305040
rect 187568 305028 187574 305040
rect 194410 305028 194416 305040
rect 187568 305000 194416 305028
rect 187568 304988 187574 305000
rect 194410 304988 194416 305000
rect 194468 304988 194474 305040
rect 227622 304716 227628 304768
rect 227680 304756 227686 304768
rect 229186 304756 229192 304768
rect 227680 304728 229192 304756
rect 227680 304716 227686 304728
rect 229186 304716 229192 304728
rect 229244 304716 229250 304768
rect 246298 304648 246304 304700
rect 246356 304688 246362 304700
rect 250162 304688 250168 304700
rect 246356 304660 250168 304688
rect 246356 304648 246362 304660
rect 250162 304648 250168 304660
rect 250220 304648 250226 304700
rect 230382 304308 230388 304360
rect 230440 304348 230446 304360
rect 246574 304348 246580 304360
rect 230440 304320 246580 304348
rect 230440 304308 230446 304320
rect 246574 304308 246580 304320
rect 246632 304308 246638 304360
rect 97166 304240 97172 304292
rect 97224 304280 97230 304292
rect 160186 304280 160192 304292
rect 97224 304252 160192 304280
rect 97224 304240 97230 304252
rect 160186 304240 160192 304252
rect 160244 304240 160250 304292
rect 213178 304240 213184 304292
rect 213236 304280 213242 304292
rect 232774 304280 232780 304292
rect 213236 304252 232780 304280
rect 213236 304240 213242 304252
rect 232774 304240 232780 304252
rect 232832 304240 232838 304292
rect 249150 304240 249156 304292
rect 249208 304280 249214 304292
rect 258166 304280 258172 304292
rect 249208 304252 258172 304280
rect 249208 304240 249214 304252
rect 258166 304240 258172 304252
rect 258224 304240 258230 304292
rect 259454 304240 259460 304292
rect 259512 304280 259518 304292
rect 277578 304280 277584 304292
rect 259512 304252 277584 304280
rect 259512 304240 259518 304252
rect 277578 304240 277584 304252
rect 277636 304280 277642 304292
rect 289998 304280 290004 304292
rect 277636 304252 290004 304280
rect 277636 304240 277642 304252
rect 289998 304240 290004 304252
rect 290056 304240 290062 304292
rect 244734 304036 244740 304088
rect 244792 304076 244798 304088
rect 246942 304076 246948 304088
rect 244792 304048 246948 304076
rect 244792 304036 244798 304048
rect 246942 304036 246948 304048
rect 247000 304036 247006 304088
rect 213822 303832 213828 303884
rect 213880 303872 213886 303884
rect 222010 303872 222016 303884
rect 213880 303844 222016 303872
rect 213880 303832 213886 303844
rect 222010 303832 222016 303844
rect 222068 303832 222074 303884
rect 189810 303696 189816 303748
rect 189868 303736 189874 303748
rect 195606 303736 195612 303748
rect 189868 303708 195612 303736
rect 189868 303696 189874 303708
rect 195606 303696 195612 303708
rect 195664 303696 195670 303748
rect 198734 303696 198740 303748
rect 198792 303736 198798 303748
rect 201034 303736 201040 303748
rect 198792 303708 201040 303736
rect 198792 303696 198798 303708
rect 201034 303696 201040 303708
rect 201092 303696 201098 303748
rect 151078 303628 151084 303680
rect 151136 303668 151142 303680
rect 212074 303668 212080 303680
rect 151136 303640 212080 303668
rect 151136 303628 151142 303640
rect 212074 303628 212080 303640
rect 212132 303628 212138 303680
rect 213914 303628 213920 303680
rect 213972 303668 213978 303680
rect 214558 303668 214564 303680
rect 213972 303640 214564 303668
rect 213972 303628 213978 303640
rect 214558 303628 214564 303640
rect 214616 303628 214622 303680
rect 219434 303628 219440 303680
rect 219492 303668 219498 303680
rect 219894 303668 219900 303680
rect 219492 303640 219900 303668
rect 219492 303628 219498 303640
rect 219894 303628 219900 303640
rect 219952 303628 219958 303680
rect 224954 303628 224960 303680
rect 225012 303668 225018 303680
rect 225230 303668 225236 303680
rect 225012 303640 225236 303668
rect 225012 303628 225018 303640
rect 225230 303628 225236 303640
rect 225288 303628 225294 303680
rect 232222 303628 232228 303680
rect 232280 303668 232286 303680
rect 233142 303668 233148 303680
rect 232280 303640 233148 303668
rect 232280 303628 232286 303640
rect 233142 303628 233148 303640
rect 233200 303628 233206 303680
rect 233878 303628 233884 303680
rect 233936 303668 233942 303680
rect 234614 303668 234620 303680
rect 233936 303640 234620 303668
rect 233936 303628 233942 303640
rect 234614 303628 234620 303640
rect 234672 303628 234678 303680
rect 239398 303628 239404 303680
rect 239456 303668 239462 303680
rect 242802 303668 242808 303680
rect 239456 303640 242808 303668
rect 239456 303628 239462 303640
rect 242802 303628 242808 303640
rect 242860 303628 242866 303680
rect 242894 303628 242900 303680
rect 242952 303668 242958 303680
rect 243814 303668 243820 303680
rect 242952 303640 243820 303668
rect 242952 303628 242958 303640
rect 243814 303628 243820 303640
rect 243872 303628 243878 303680
rect 248414 303628 248420 303680
rect 248472 303668 248478 303680
rect 249610 303668 249616 303680
rect 248472 303640 249616 303668
rect 248472 303628 248478 303640
rect 249610 303628 249616 303640
rect 249668 303628 249674 303680
rect 250806 303628 250812 303680
rect 250864 303668 250870 303680
rect 262490 303668 262496 303680
rect 250864 303640 262496 303668
rect 250864 303628 250870 303640
rect 262490 303628 262496 303640
rect 262548 303628 262554 303680
rect 195974 303560 195980 303612
rect 196032 303600 196038 303612
rect 196710 303600 196716 303612
rect 196032 303572 196716 303600
rect 196032 303560 196038 303572
rect 196710 303560 196716 303572
rect 196768 303560 196774 303612
rect 201494 303560 201500 303612
rect 201552 303600 201558 303612
rect 201862 303600 201868 303612
rect 201552 303572 201868 303600
rect 201552 303560 201558 303572
rect 201862 303560 201868 303572
rect 201920 303560 201926 303612
rect 72694 302880 72700 302932
rect 72752 302920 72758 302932
rect 175182 302920 175188 302932
rect 72752 302892 175188 302920
rect 72752 302880 72758 302892
rect 175182 302880 175188 302892
rect 175240 302880 175246 302932
rect 220814 302880 220820 302932
rect 220872 302920 220878 302932
rect 232498 302920 232504 302932
rect 220872 302892 232504 302920
rect 220872 302880 220878 302892
rect 232498 302880 232504 302892
rect 232556 302880 232562 302932
rect 187694 302268 187700 302320
rect 187752 302308 187758 302320
rect 218422 302308 218428 302320
rect 187752 302280 218428 302308
rect 187752 302268 187758 302280
rect 218422 302268 218428 302280
rect 218480 302308 218486 302320
rect 219342 302308 219348 302320
rect 218480 302280 219348 302308
rect 218480 302268 218486 302280
rect 219342 302268 219348 302280
rect 219400 302268 219406 302320
rect 240594 302268 240600 302320
rect 240652 302308 240658 302320
rect 241422 302308 241428 302320
rect 240652 302280 241428 302308
rect 240652 302268 240658 302280
rect 241422 302268 241428 302280
rect 241480 302308 241486 302320
rect 268010 302308 268016 302320
rect 241480 302280 268016 302308
rect 241480 302268 241486 302280
rect 268010 302268 268016 302280
rect 268068 302268 268074 302320
rect 171778 302200 171784 302252
rect 171836 302240 171842 302252
rect 172238 302240 172244 302252
rect 171836 302212 172244 302240
rect 171836 302200 171842 302212
rect 172238 302200 172244 302212
rect 172296 302240 172302 302252
rect 227438 302240 227444 302252
rect 172296 302212 227444 302240
rect 172296 302200 172302 302212
rect 227438 302200 227444 302212
rect 227496 302200 227502 302252
rect 240042 302200 240048 302252
rect 240100 302240 240106 302252
rect 271966 302240 271972 302252
rect 240100 302212 271972 302240
rect 240100 302200 240106 302212
rect 271966 302200 271972 302212
rect 272024 302200 272030 302252
rect 186314 302132 186320 302184
rect 186372 302172 186378 302184
rect 191466 302172 191472 302184
rect 186372 302144 191472 302172
rect 186372 302132 186378 302144
rect 191466 302132 191472 302144
rect 191524 302132 191530 302184
rect 228450 302132 228456 302184
rect 228508 302172 228514 302184
rect 231026 302172 231032 302184
rect 228508 302144 231032 302172
rect 228508 302132 228514 302144
rect 231026 302132 231032 302144
rect 231084 302132 231090 302184
rect 92290 301520 92296 301572
rect 92348 301560 92354 301572
rect 96614 301560 96620 301572
rect 92348 301532 96620 301560
rect 92348 301520 92354 301532
rect 96614 301520 96620 301532
rect 96672 301520 96678 301572
rect 250438 301520 250444 301572
rect 250496 301560 250502 301572
rect 256786 301560 256792 301572
rect 250496 301532 256792 301560
rect 250496 301520 250502 301532
rect 256786 301520 256792 301532
rect 256844 301520 256850 301572
rect 94590 301452 94596 301504
rect 94648 301492 94654 301504
rect 135990 301492 135996 301504
rect 94648 301464 135996 301492
rect 94648 301452 94654 301464
rect 135990 301452 135996 301464
rect 136048 301452 136054 301504
rect 193122 300908 193128 300960
rect 193180 300948 193186 300960
rect 197630 300948 197636 300960
rect 193180 300920 197636 300948
rect 193180 300908 193186 300920
rect 197630 300908 197636 300920
rect 197688 300908 197694 300960
rect 237374 300948 237380 300960
rect 219406 300920 237380 300948
rect 175642 300840 175648 300892
rect 175700 300880 175706 300892
rect 219406 300880 219434 300920
rect 237374 300908 237380 300920
rect 237432 300948 237438 300960
rect 238662 300948 238668 300960
rect 237432 300920 238668 300948
rect 237432 300908 237438 300920
rect 238662 300908 238668 300920
rect 238720 300908 238726 300960
rect 175700 300852 219434 300880
rect 175700 300840 175706 300852
rect 252370 300840 252376 300892
rect 252428 300880 252434 300892
rect 252830 300880 252836 300892
rect 252428 300852 252836 300880
rect 252428 300840 252434 300852
rect 252830 300840 252836 300852
rect 252888 300840 252894 300892
rect 255590 300840 255596 300892
rect 255648 300880 255654 300892
rect 255958 300880 255964 300892
rect 255648 300852 255964 300880
rect 255648 300840 255654 300852
rect 255958 300840 255964 300852
rect 256016 300880 256022 300892
rect 288618 300880 288624 300892
rect 256016 300852 288624 300880
rect 256016 300840 256022 300852
rect 288618 300840 288624 300852
rect 288676 300840 288682 300892
rect 170398 300772 170404 300824
rect 170456 300812 170462 300824
rect 172238 300812 172244 300824
rect 170456 300784 172244 300812
rect 170456 300772 170462 300784
rect 172238 300772 172244 300784
rect 172296 300772 172302 300824
rect 183462 300772 183468 300824
rect 183520 300812 183526 300824
rect 186958 300812 186964 300824
rect 183520 300784 186964 300812
rect 183520 300772 183526 300784
rect 186958 300772 186964 300784
rect 187016 300772 187022 300824
rect 259270 300160 259276 300212
rect 259328 300200 259334 300212
rect 281534 300200 281540 300212
rect 259328 300172 281540 300200
rect 259328 300160 259334 300172
rect 281534 300160 281540 300172
rect 281592 300160 281598 300212
rect 169202 300092 169208 300144
rect 169260 300132 169266 300144
rect 187694 300132 187700 300144
rect 169260 300104 187700 300132
rect 169260 300092 169266 300104
rect 187694 300092 187700 300104
rect 187752 300092 187758 300144
rect 262122 300092 262128 300144
rect 262180 300132 262186 300144
rect 287054 300132 287060 300144
rect 262180 300104 287060 300132
rect 262180 300092 262186 300104
rect 287054 300092 287060 300104
rect 287112 300132 287118 300144
rect 303614 300132 303620 300144
rect 287112 300104 303620 300132
rect 287112 300092 287118 300104
rect 303614 300092 303620 300104
rect 303672 300092 303678 300144
rect 255498 300024 255504 300076
rect 255556 300064 255562 300076
rect 259270 300064 259276 300076
rect 255556 300036 259276 300064
rect 255556 300024 255562 300036
rect 259270 300024 259276 300036
rect 259328 300024 259334 300076
rect 188338 299616 188344 299668
rect 188396 299656 188402 299668
rect 193674 299656 193680 299668
rect 188396 299628 193680 299656
rect 188396 299616 188402 299628
rect 193674 299616 193680 299628
rect 193732 299616 193738 299668
rect 162210 299412 162216 299464
rect 162268 299452 162274 299464
rect 185670 299452 185676 299464
rect 162268 299424 185676 299452
rect 162268 299412 162274 299424
rect 185670 299412 185676 299424
rect 185728 299412 185734 299464
rect 255498 299412 255504 299464
rect 255556 299452 255562 299464
rect 262122 299452 262128 299464
rect 255556 299424 262128 299452
rect 255556 299412 255562 299424
rect 262122 299412 262128 299424
rect 262180 299412 262186 299464
rect 129182 298800 129188 298852
rect 129240 298840 129246 298852
rect 159358 298840 159364 298852
rect 129240 298812 159364 298840
rect 129240 298800 129246 298812
rect 159358 298800 159364 298812
rect 159416 298800 159422 298852
rect 148318 298732 148324 298784
rect 148376 298772 148382 298784
rect 187786 298772 187792 298784
rect 148376 298744 187792 298772
rect 148376 298732 148382 298744
rect 187786 298732 187792 298744
rect 187844 298732 187850 298784
rect 187602 298120 187608 298172
rect 187660 298160 187666 298172
rect 191466 298160 191472 298172
rect 187660 298132 191472 298160
rect 187660 298120 187666 298132
rect 191466 298120 191472 298132
rect 191524 298120 191530 298172
rect 255498 298120 255504 298172
rect 255556 298160 255562 298172
rect 271138 298160 271144 298172
rect 255556 298132 271144 298160
rect 255556 298120 255562 298132
rect 271138 298120 271144 298132
rect 271196 298120 271202 298172
rect 118694 297372 118700 297424
rect 118752 297412 118758 297424
rect 175642 297412 175648 297424
rect 118752 297384 175648 297412
rect 118752 297372 118758 297384
rect 175642 297372 175648 297384
rect 175700 297372 175706 297424
rect 265618 297372 265624 297424
rect 265676 297412 265682 297424
rect 296806 297412 296812 297424
rect 265676 297384 296812 297412
rect 265676 297372 265682 297384
rect 296806 297372 296812 297384
rect 296864 297372 296870 297424
rect 255498 296760 255504 296812
rect 255556 296800 255562 296812
rect 263778 296800 263784 296812
rect 255556 296772 263784 296800
rect 255556 296760 255562 296772
rect 263778 296760 263784 296772
rect 263836 296760 263842 296812
rect 171134 296692 171140 296744
rect 171192 296732 171198 296744
rect 191466 296732 191472 296744
rect 171192 296704 191472 296732
rect 171192 296692 171198 296704
rect 191466 296692 191472 296704
rect 191524 296692 191530 296744
rect 256050 296692 256056 296744
rect 256108 296732 256114 296744
rect 276198 296732 276204 296744
rect 256108 296704 276204 296732
rect 256108 296692 256114 296704
rect 276198 296692 276204 296704
rect 276256 296692 276262 296744
rect 255498 296556 255504 296608
rect 255556 296596 255562 296608
rect 259822 296596 259828 296608
rect 255556 296568 259828 296596
rect 255556 296556 255562 296568
rect 259822 296556 259828 296568
rect 259880 296596 259886 296608
rect 260742 296596 260748 296608
rect 259880 296568 260748 296596
rect 259880 296556 259886 296568
rect 260742 296556 260748 296568
rect 260800 296556 260806 296608
rect 86954 296012 86960 296064
rect 87012 296052 87018 296064
rect 116670 296052 116676 296064
rect 87012 296024 116676 296052
rect 87012 296012 87018 296024
rect 116670 296012 116676 296024
rect 116728 296012 116734 296064
rect 117222 296012 117228 296064
rect 117280 296052 117286 296064
rect 175918 296052 175924 296064
rect 117280 296024 175924 296052
rect 117280 296012 117286 296024
rect 175918 296012 175924 296024
rect 175976 296012 175982 296064
rect 67266 295944 67272 295996
rect 67324 295984 67330 295996
rect 166442 295984 166448 295996
rect 67324 295956 166448 295984
rect 67324 295944 67330 295956
rect 166442 295944 166448 295956
rect 166500 295984 166506 295996
rect 174538 295984 174544 295996
rect 166500 295956 174544 295984
rect 166500 295944 166506 295956
rect 174538 295944 174544 295956
rect 174596 295984 174602 295996
rect 189994 295984 190000 295996
rect 174596 295956 190000 295984
rect 174596 295944 174602 295956
rect 189994 295944 190000 295956
rect 190052 295944 190058 295996
rect 253934 295604 253940 295656
rect 253992 295644 253998 295656
rect 259454 295644 259460 295656
rect 253992 295616 259460 295644
rect 253992 295604 253998 295616
rect 259454 295604 259460 295616
rect 259512 295604 259518 295656
rect 260742 295332 260748 295384
rect 260800 295372 260806 295384
rect 288434 295372 288440 295384
rect 260800 295344 288440 295372
rect 260800 295332 260806 295344
rect 288434 295332 288440 295344
rect 288492 295332 288498 295384
rect 255314 295264 255320 295316
rect 255372 295304 255378 295316
rect 272150 295304 272156 295316
rect 255372 295276 272156 295304
rect 255372 295264 255378 295276
rect 272150 295264 272156 295276
rect 272208 295264 272214 295316
rect 156598 294652 156604 294704
rect 156656 294692 156662 294704
rect 184842 294692 184848 294704
rect 156656 294664 184848 294692
rect 156656 294652 156662 294664
rect 184842 294652 184848 294664
rect 184900 294652 184906 294704
rect 186222 294652 186228 294704
rect 186280 294692 186286 294704
rect 191466 294692 191472 294704
rect 186280 294664 191472 294692
rect 186280 294652 186286 294664
rect 191466 294652 191472 294664
rect 191524 294652 191530 294704
rect 65886 294584 65892 294636
rect 65944 294624 65950 294636
rect 160094 294624 160100 294636
rect 65944 294596 160100 294624
rect 65944 294584 65950 294596
rect 160094 294584 160100 294596
rect 160152 294624 160158 294636
rect 163590 294624 163596 294636
rect 160152 294596 163596 294624
rect 160152 294584 160158 294596
rect 163590 294584 163596 294596
rect 163648 294584 163654 294636
rect 272150 294584 272156 294636
rect 272208 294624 272214 294636
rect 285950 294624 285956 294636
rect 272208 294596 285956 294624
rect 272208 294584 272214 294596
rect 285950 294584 285956 294596
rect 286008 294584 286014 294636
rect 176194 293972 176200 294024
rect 176252 294012 176258 294024
rect 178862 294012 178868 294024
rect 176252 293984 178868 294012
rect 176252 293972 176258 293984
rect 178862 293972 178868 293984
rect 178920 293972 178926 294024
rect 184842 293972 184848 294024
rect 184900 294012 184906 294024
rect 186222 294012 186228 294024
rect 184900 293984 186228 294012
rect 184900 293972 184906 293984
rect 186222 293972 186228 293984
rect 186280 293972 186286 294024
rect 255406 293972 255412 294024
rect 255464 294012 255470 294024
rect 298094 294012 298100 294024
rect 255464 293984 298100 294012
rect 255464 293972 255470 293984
rect 298094 293972 298100 293984
rect 298152 293972 298158 294024
rect 92566 293904 92572 293956
rect 92624 293944 92630 293956
rect 93762 293944 93768 293956
rect 92624 293916 93768 293944
rect 92624 293904 92630 293916
rect 93762 293904 93768 293916
rect 93820 293944 93826 293956
rect 133782 293944 133788 293956
rect 93820 293916 133788 293944
rect 93820 293904 93826 293916
rect 133782 293904 133788 293916
rect 133840 293904 133846 293956
rect 171134 293332 171140 293344
rect 161446 293304 171140 293332
rect 133782 293224 133788 293276
rect 133840 293264 133846 293276
rect 159358 293264 159364 293276
rect 133840 293236 159364 293264
rect 133840 293224 133846 293236
rect 159358 293224 159364 293236
rect 159416 293264 159422 293276
rect 161446 293264 161474 293304
rect 171134 293292 171140 293304
rect 171192 293292 171198 293344
rect 256694 293292 256700 293344
rect 256752 293332 256758 293344
rect 289906 293332 289912 293344
rect 256752 293304 289912 293332
rect 256752 293292 256758 293304
rect 289906 293292 289912 293304
rect 289964 293292 289970 293344
rect 159416 293236 161474 293264
rect 159416 293224 159422 293236
rect 171778 293224 171784 293276
rect 171836 293264 171842 293276
rect 187602 293264 187608 293276
rect 171836 293236 187608 293264
rect 171836 293224 171842 293236
rect 187602 293224 187608 293236
rect 187660 293224 187666 293276
rect 255406 293224 255412 293276
rect 255464 293264 255470 293276
rect 259362 293264 259368 293276
rect 255464 293236 259368 293264
rect 255464 293224 255470 293236
rect 259362 293224 259368 293236
rect 259420 293264 259426 293276
rect 299474 293264 299480 293276
rect 259420 293236 299480 293264
rect 259420 293224 259426 293236
rect 299474 293224 299480 293236
rect 299532 293224 299538 293276
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 14458 292584 14464 292596
rect 3476 292556 14464 292584
rect 3476 292544 3482 292556
rect 14458 292544 14464 292556
rect 14516 292544 14522 292596
rect 82170 292544 82176 292596
rect 82228 292584 82234 292596
rect 82630 292584 82636 292596
rect 82228 292556 82636 292584
rect 82228 292544 82234 292556
rect 82630 292544 82636 292556
rect 82688 292584 82694 292596
rect 113818 292584 113824 292596
rect 82688 292556 113824 292584
rect 82688 292544 82694 292556
rect 113818 292544 113824 292556
rect 113876 292544 113882 292596
rect 191466 292584 191472 292596
rect 184676 292556 191472 292584
rect 157242 292476 157248 292528
rect 157300 292516 157306 292528
rect 164050 292516 164056 292528
rect 157300 292488 164056 292516
rect 157300 292476 157306 292488
rect 164050 292476 164056 292488
rect 164108 292516 164114 292528
rect 184676 292516 184704 292556
rect 191466 292544 191472 292556
rect 191524 292544 191530 292596
rect 164108 292488 184704 292516
rect 164108 292476 164114 292488
rect 176102 292408 176108 292460
rect 176160 292448 176166 292460
rect 180058 292448 180064 292460
rect 176160 292420 180064 292448
rect 176160 292408 176166 292420
rect 180058 292408 180064 292420
rect 180116 292448 180122 292460
rect 191466 292448 191472 292460
rect 180116 292420 191472 292448
rect 180116 292408 180122 292420
rect 191466 292408 191472 292420
rect 191524 292408 191530 292460
rect 256602 291864 256608 291916
rect 256660 291904 256666 291916
rect 263594 291904 263600 291916
rect 256660 291876 263600 291904
rect 256660 291864 256666 291876
rect 263594 291864 263600 291876
rect 263652 291864 263658 291916
rect 262858 291796 262864 291848
rect 262916 291836 262922 291848
rect 280246 291836 280252 291848
rect 262916 291808 280252 291836
rect 262916 291796 262922 291808
rect 280246 291796 280252 291808
rect 280304 291796 280310 291848
rect 86218 291592 86224 291644
rect 86276 291632 86282 291644
rect 93118 291632 93124 291644
rect 86276 291604 93124 291632
rect 86276 291592 86282 291604
rect 93118 291592 93124 291604
rect 93176 291592 93182 291644
rect 98270 291184 98276 291236
rect 98328 291224 98334 291236
rect 99282 291224 99288 291236
rect 98328 291196 99288 291224
rect 98328 291184 98334 291196
rect 99282 291184 99288 291196
rect 99340 291224 99346 291236
rect 157242 291224 157248 291236
rect 99340 291196 157248 291224
rect 99340 291184 99346 291196
rect 157242 291184 157248 291196
rect 157300 291184 157306 291236
rect 67542 291116 67548 291168
rect 67600 291156 67606 291168
rect 68554 291156 68560 291168
rect 67600 291128 68560 291156
rect 67600 291116 67606 291128
rect 68554 291116 68560 291128
rect 68612 291156 68618 291168
rect 131114 291156 131120 291168
rect 68612 291128 131120 291156
rect 68612 291116 68618 291128
rect 131114 291116 131120 291128
rect 131172 291116 131178 291168
rect 256510 291048 256516 291100
rect 256568 291088 256574 291100
rect 260834 291088 260840 291100
rect 256568 291060 260840 291088
rect 256568 291048 256574 291060
rect 260834 291048 260840 291060
rect 260892 291048 260898 291100
rect 131114 290436 131120 290488
rect 131172 290476 131178 290488
rect 132402 290476 132408 290488
rect 131172 290448 132408 290476
rect 131172 290436 131178 290448
rect 132402 290436 132408 290448
rect 132460 290476 132466 290488
rect 163682 290476 163688 290488
rect 132460 290448 163688 290476
rect 132460 290436 132466 290448
rect 163682 290436 163688 290448
rect 163740 290436 163746 290488
rect 261478 290436 261484 290488
rect 261536 290476 261542 290488
rect 265066 290476 265072 290488
rect 261536 290448 265072 290476
rect 261536 290436 261542 290448
rect 265066 290436 265072 290448
rect 265124 290436 265130 290488
rect 186038 289960 186044 290012
rect 186096 290000 186102 290012
rect 190822 290000 190828 290012
rect 186096 289972 190828 290000
rect 186096 289960 186102 289972
rect 190822 289960 190828 289972
rect 190880 289960 190886 290012
rect 170490 289892 170496 289944
rect 170548 289932 170554 289944
rect 191466 289932 191472 289944
rect 170548 289904 191472 289932
rect 170548 289892 170554 289904
rect 191466 289892 191472 289904
rect 191524 289892 191530 289944
rect 84562 289824 84568 289876
rect 84620 289864 84626 289876
rect 177390 289864 177396 289876
rect 84620 289836 177396 289864
rect 84620 289824 84626 289836
rect 177390 289824 177396 289836
rect 177448 289824 177454 289876
rect 256510 289824 256516 289876
rect 256568 289864 256574 289876
rect 582558 289864 582564 289876
rect 256568 289836 582564 289864
rect 256568 289824 256574 289836
rect 582558 289824 582564 289836
rect 582616 289824 582622 289876
rect 256602 289756 256608 289808
rect 256660 289796 256666 289808
rect 267734 289796 267740 289808
rect 256660 289768 267740 289796
rect 256660 289756 256666 289768
rect 267734 289756 267740 289768
rect 267792 289756 267798 289808
rect 71590 289144 71596 289196
rect 71648 289184 71654 289196
rect 117222 289184 117228 289196
rect 71648 289156 117228 289184
rect 71648 289144 71654 289156
rect 117222 289144 117228 289156
rect 117280 289144 117286 289196
rect 164970 289144 164976 289196
rect 165028 289184 165034 289196
rect 187602 289184 187608 289196
rect 165028 289156 187608 289184
rect 165028 289144 165034 289156
rect 187602 289144 187608 289156
rect 187660 289144 187666 289196
rect 78950 289076 78956 289128
rect 79008 289116 79014 289128
rect 79962 289116 79968 289128
rect 79008 289088 79968 289116
rect 79008 289076 79014 289088
rect 79962 289076 79968 289088
rect 80020 289116 80026 289128
rect 159450 289116 159456 289128
rect 80020 289088 159456 289116
rect 80020 289076 80026 289088
rect 159450 289076 159456 289088
rect 159508 289116 159514 289128
rect 160002 289116 160008 289128
rect 159508 289088 160008 289116
rect 159508 289076 159514 289088
rect 160002 289076 160008 289088
rect 160060 289116 160066 289128
rect 191466 289116 191472 289128
rect 160060 289088 191472 289116
rect 160060 289076 160066 289088
rect 191466 289076 191472 289088
rect 191524 289076 191530 289128
rect 256510 289076 256516 289128
rect 256568 289116 256574 289128
rect 259454 289116 259460 289128
rect 256568 289088 259460 289116
rect 256568 289076 256574 289088
rect 259454 289076 259460 289088
rect 259512 289116 259518 289128
rect 269298 289116 269304 289128
rect 259512 289088 269304 289116
rect 259512 289076 259518 289088
rect 269298 289076 269304 289088
rect 269356 289076 269362 289128
rect 56410 288396 56416 288448
rect 56468 288436 56474 288448
rect 72510 288436 72516 288448
rect 56468 288408 72516 288436
rect 56468 288396 56474 288408
rect 72510 288396 72516 288408
rect 72568 288436 72574 288448
rect 72786 288436 72792 288448
rect 72568 288408 72792 288436
rect 72568 288396 72574 288408
rect 72786 288396 72792 288408
rect 72844 288396 72850 288448
rect 80054 288328 80060 288380
rect 80112 288368 80118 288380
rect 80698 288368 80704 288380
rect 80112 288340 80704 288368
rect 80112 288328 80118 288340
rect 80698 288328 80704 288340
rect 80756 288328 80762 288380
rect 255866 288328 255872 288380
rect 255924 288368 255930 288380
rect 277394 288368 277400 288380
rect 255924 288340 277400 288368
rect 255924 288328 255930 288340
rect 277394 288328 277400 288340
rect 277452 288328 277458 288380
rect 85850 287920 85856 287972
rect 85908 287960 85914 287972
rect 86770 287960 86776 287972
rect 85908 287932 86776 287960
rect 85908 287920 85914 287932
rect 86770 287920 86776 287932
rect 86828 287920 86834 287972
rect 92474 287716 92480 287768
rect 92532 287756 92538 287768
rect 92934 287756 92940 287768
rect 92532 287728 92940 287756
rect 92532 287716 92538 287728
rect 92934 287716 92940 287728
rect 92992 287716 92998 287768
rect 104618 287716 104624 287768
rect 104676 287756 104682 287768
rect 115198 287756 115204 287768
rect 104676 287728 115204 287756
rect 104676 287716 104682 287728
rect 115198 287716 115204 287728
rect 115256 287716 115262 287768
rect 115290 287716 115296 287768
rect 115348 287756 115354 287768
rect 169662 287756 169668 287768
rect 115348 287728 169668 287756
rect 115348 287716 115354 287728
rect 169662 287716 169668 287728
rect 169720 287756 169726 287768
rect 184750 287756 184756 287768
rect 169720 287728 184756 287756
rect 169720 287716 169726 287728
rect 184750 287716 184756 287728
rect 184808 287756 184814 287768
rect 191466 287756 191472 287768
rect 184808 287728 191472 287756
rect 184808 287716 184814 287728
rect 191466 287716 191472 287728
rect 191524 287716 191530 287768
rect 255958 287716 255964 287768
rect 256016 287756 256022 287768
rect 259546 287756 259552 287768
rect 256016 287728 259552 287756
rect 256016 287716 256022 287728
rect 259546 287716 259552 287728
rect 259604 287716 259610 287768
rect 43438 287648 43444 287700
rect 43496 287688 43502 287700
rect 70486 287688 70492 287700
rect 43496 287660 70492 287688
rect 43496 287648 43502 287660
rect 70486 287648 70492 287660
rect 70544 287648 70550 287700
rect 78582 287648 78588 287700
rect 78640 287688 78646 287700
rect 184198 287688 184204 287700
rect 78640 287660 184204 287688
rect 78640 287648 78646 287660
rect 184198 287648 184204 287660
rect 184256 287648 184262 287700
rect 271138 287648 271144 287700
rect 271196 287688 271202 287700
rect 284938 287688 284944 287700
rect 271196 287660 284944 287688
rect 271196 287648 271202 287660
rect 284938 287648 284944 287660
rect 284996 287688 285002 287700
rect 302234 287688 302240 287700
rect 284996 287660 302240 287688
rect 284996 287648 285002 287660
rect 302234 287648 302240 287660
rect 302292 287648 302298 287700
rect 73890 287036 73896 287088
rect 73948 287076 73954 287088
rect 80054 287076 80060 287088
rect 73948 287048 80060 287076
rect 73948 287036 73954 287048
rect 80054 287036 80060 287048
rect 80112 287036 80118 287088
rect 86770 287036 86776 287088
rect 86828 287076 86834 287088
rect 102134 287076 102140 287088
rect 86828 287048 102140 287076
rect 86828 287036 86834 287048
rect 102134 287036 102140 287048
rect 102192 287036 102198 287088
rect 91922 286968 91928 287020
rect 91980 287008 91986 287020
rect 92382 287008 92388 287020
rect 91980 286980 92388 287008
rect 91980 286968 91986 286980
rect 92382 286968 92388 286980
rect 92440 286968 92446 287020
rect 142890 286968 142896 287020
rect 142948 287008 142954 287020
rect 185578 287008 185584 287020
rect 142948 286980 185584 287008
rect 142948 286968 142954 286980
rect 185578 286968 185584 286980
rect 185636 286968 185642 287020
rect 255866 286968 255872 287020
rect 255924 287008 255930 287020
rect 294046 287008 294052 287020
rect 255924 286980 294052 287008
rect 255924 286968 255930 286980
rect 294046 286968 294052 286980
rect 294104 286968 294110 287020
rect 95326 286696 95332 286748
rect 95384 286736 95390 286748
rect 97258 286736 97264 286748
rect 95384 286708 97264 286736
rect 95384 286696 95390 286708
rect 97258 286696 97264 286708
rect 97316 286696 97322 286748
rect 74718 286396 74724 286408
rect 64846 286368 74724 286396
rect 52086 286288 52092 286340
rect 52144 286328 52150 286340
rect 60642 286328 60648 286340
rect 52144 286300 60648 286328
rect 52144 286288 52150 286300
rect 60642 286288 60648 286300
rect 60700 286328 60706 286340
rect 64846 286328 64874 286368
rect 74718 286356 74724 286368
rect 74776 286356 74782 286408
rect 60700 286300 64874 286328
rect 60700 286288 60706 286300
rect 75730 286288 75736 286340
rect 75788 286328 75794 286340
rect 142890 286328 142896 286340
rect 75788 286300 142896 286328
rect 75788 286288 75794 286300
rect 142890 286288 142896 286300
rect 142948 286288 142954 286340
rect 173618 286288 173624 286340
rect 173676 286328 173682 286340
rect 186314 286328 186320 286340
rect 173676 286300 186320 286328
rect 173676 286288 173682 286300
rect 186314 286288 186320 286300
rect 186372 286328 186378 286340
rect 191466 286328 191472 286340
rect 186372 286300 191472 286328
rect 186372 286288 186378 286300
rect 191466 286288 191472 286300
rect 191524 286288 191530 286340
rect 82354 286220 82360 286272
rect 82412 286260 82418 286272
rect 83458 286260 83464 286272
rect 82412 286232 83464 286260
rect 82412 286220 82418 286232
rect 83458 286220 83464 286232
rect 83516 286220 83522 286272
rect 91370 285880 91376 285932
rect 91428 285920 91434 285932
rect 94590 285920 94596 285932
rect 91428 285892 94596 285920
rect 91428 285880 91434 285892
rect 94590 285880 94596 285892
rect 94648 285880 94654 285932
rect 187602 285880 187608 285932
rect 187660 285920 187666 285932
rect 191374 285920 191380 285932
rect 187660 285892 191380 285920
rect 187660 285880 187666 285892
rect 191374 285880 191380 285892
rect 191432 285880 191438 285932
rect 80974 285784 80980 285796
rect 64846 285756 80980 285784
rect 60366 285676 60372 285728
rect 60424 285716 60430 285728
rect 64846 285716 64874 285756
rect 80974 285744 80980 285756
rect 81032 285744 81038 285796
rect 60424 285688 64874 285716
rect 60424 285676 60430 285688
rect 80882 285676 80888 285728
rect 80940 285716 80946 285728
rect 82170 285716 82176 285728
rect 80940 285688 82176 285716
rect 80940 285676 80946 285688
rect 82170 285676 82176 285688
rect 82228 285676 82234 285728
rect 84286 285676 84292 285728
rect 84344 285716 84350 285728
rect 90358 285716 90364 285728
rect 84344 285688 90364 285716
rect 84344 285676 84350 285688
rect 90358 285676 90364 285688
rect 90416 285676 90422 285728
rect 163498 285676 163504 285728
rect 163556 285716 163562 285728
rect 170582 285716 170588 285728
rect 163556 285688 170588 285716
rect 163556 285676 163562 285688
rect 170582 285676 170588 285688
rect 170640 285676 170646 285728
rect 256510 285676 256516 285728
rect 256568 285716 256574 285728
rect 259730 285716 259736 285728
rect 256568 285688 259736 285716
rect 256568 285676 256574 285688
rect 259730 285676 259736 285688
rect 259788 285716 259794 285728
rect 263594 285716 263600 285728
rect 259788 285688 263600 285716
rect 259788 285676 259794 285688
rect 263594 285676 263600 285688
rect 263652 285676 263658 285728
rect 171042 285608 171048 285660
rect 171100 285648 171106 285660
rect 189902 285648 189908 285660
rect 171100 285620 189908 285648
rect 171100 285608 171106 285620
rect 189902 285608 189908 285620
rect 189960 285608 189966 285660
rect 256602 285608 256608 285660
rect 256660 285648 256666 285660
rect 263870 285648 263876 285660
rect 256660 285620 263876 285648
rect 256660 285608 256666 285620
rect 263870 285608 263876 285620
rect 263928 285608 263934 285660
rect 135990 284928 135996 284980
rect 136048 284968 136054 284980
rect 148502 284968 148508 284980
rect 136048 284940 148508 284968
rect 136048 284928 136054 284940
rect 148502 284928 148508 284940
rect 148560 284928 148566 284980
rect 262214 284928 262220 284980
rect 262272 284968 262278 284980
rect 291470 284968 291476 284980
rect 262272 284940 291476 284968
rect 262272 284928 262278 284940
rect 291470 284928 291476 284940
rect 291528 284928 291534 284980
rect 50982 284384 50988 284436
rect 51040 284424 51046 284436
rect 69014 284424 69020 284436
rect 51040 284396 69020 284424
rect 51040 284384 51046 284396
rect 69014 284384 69020 284396
rect 69072 284384 69078 284436
rect 78214 284384 78220 284436
rect 78272 284424 78278 284436
rect 100018 284424 100024 284436
rect 78272 284396 100024 284424
rect 78272 284384 78278 284396
rect 100018 284384 100024 284396
rect 100076 284384 100082 284436
rect 70302 284316 70308 284368
rect 70360 284356 70366 284368
rect 99098 284356 99104 284368
rect 70360 284328 99104 284356
rect 70360 284316 70366 284328
rect 99098 284316 99104 284328
rect 99156 284316 99162 284368
rect 166350 284316 166356 284368
rect 166408 284356 166414 284368
rect 191466 284356 191472 284368
rect 166408 284328 191472 284356
rect 166408 284316 166414 284328
rect 191466 284316 191472 284328
rect 191524 284316 191530 284368
rect 125594 284248 125600 284300
rect 125652 284288 125658 284300
rect 156598 284288 156604 284300
rect 125652 284260 156604 284288
rect 125652 284248 125658 284260
rect 156598 284248 156604 284260
rect 156656 284248 156662 284300
rect 167638 284248 167644 284300
rect 167696 284288 167702 284300
rect 193122 284288 193128 284300
rect 167696 284260 193128 284288
rect 167696 284248 167702 284260
rect 193122 284248 193128 284260
rect 193180 284248 193186 284300
rect 256418 284248 256424 284300
rect 256476 284288 256482 284300
rect 266538 284288 266544 284300
rect 256476 284260 266544 284288
rect 256476 284248 256482 284260
rect 266538 284248 266544 284260
rect 266596 284248 266602 284300
rect 255774 283840 255780 283892
rect 255832 283880 255838 283892
rect 258166 283880 258172 283892
rect 255832 283852 258172 283880
rect 255832 283840 255838 283852
rect 258166 283840 258172 283852
rect 258224 283840 258230 283892
rect 76144 283704 76150 283756
rect 76202 283744 76208 283756
rect 76650 283744 76656 283756
rect 76202 283716 76656 283744
rect 76202 283704 76208 283716
rect 76650 283704 76656 283716
rect 76708 283704 76714 283756
rect 100938 283568 100944 283620
rect 100996 283608 101002 283620
rect 125594 283608 125600 283620
rect 100996 283580 125600 283608
rect 100996 283568 101002 283580
rect 125594 283568 125600 283580
rect 125652 283568 125658 283620
rect 126422 283568 126428 283620
rect 126480 283608 126486 283620
rect 137278 283608 137284 283620
rect 126480 283580 137284 283608
rect 126480 283568 126486 283580
rect 137278 283568 137284 283580
rect 137336 283568 137342 283620
rect 140130 283568 140136 283620
rect 140188 283608 140194 283620
rect 148686 283608 148692 283620
rect 140188 283580 148692 283608
rect 140188 283568 140194 283580
rect 148686 283568 148692 283580
rect 148744 283568 148750 283620
rect 259270 283568 259276 283620
rect 259328 283608 259334 283620
rect 273530 283608 273536 283620
rect 259328 283580 273536 283608
rect 259328 283568 259334 283580
rect 273530 283568 273536 283580
rect 273588 283568 273594 283620
rect 70366 283104 80054 283132
rect 68830 283024 68836 283076
rect 68888 283064 68894 283076
rect 69198 283064 69204 283076
rect 68888 283036 69204 283064
rect 68888 283024 68894 283036
rect 69198 283024 69204 283036
rect 69256 283024 69262 283076
rect 58986 282956 58992 283008
rect 59044 282996 59050 283008
rect 70366 282996 70394 283104
rect 59044 282968 70394 282996
rect 59044 282956 59050 282968
rect 70762 282956 70768 283008
rect 70820 282956 70826 283008
rect 80026 282996 80054 283104
rect 98730 282996 98736 283008
rect 80026 282968 98736 282996
rect 98730 282956 98736 282968
rect 98788 282956 98794 283008
rect 70780 282928 70808 282956
rect 99374 282928 99380 282940
rect 70780 282900 99380 282928
rect 99374 282888 99380 282900
rect 99432 282888 99438 282940
rect 175918 282888 175924 282940
rect 175976 282928 175982 282940
rect 178678 282928 178684 282940
rect 175976 282900 178684 282928
rect 175976 282888 175982 282900
rect 178678 282888 178684 282900
rect 178736 282888 178742 282940
rect 255498 282820 255504 282872
rect 255556 282860 255562 282872
rect 271874 282860 271880 282872
rect 255556 282832 271880 282860
rect 255556 282820 255562 282832
rect 271874 282820 271880 282832
rect 271932 282820 271938 282872
rect 255406 282752 255412 282804
rect 255464 282792 255470 282804
rect 264974 282792 264980 282804
rect 255464 282764 264980 282792
rect 255464 282752 255470 282764
rect 264974 282752 264980 282764
rect 265032 282752 265038 282804
rect 271874 282412 271880 282464
rect 271932 282452 271938 282464
rect 273346 282452 273352 282464
rect 271932 282424 273352 282452
rect 271932 282412 271938 282424
rect 273346 282412 273352 282424
rect 273404 282412 273410 282464
rect 100754 281596 100760 281648
rect 100812 281636 100818 281648
rect 115198 281636 115204 281648
rect 100812 281608 115204 281636
rect 100812 281596 100818 281608
rect 115198 281596 115204 281608
rect 115256 281596 115262 281648
rect 160830 281596 160836 281648
rect 160888 281636 160894 281648
rect 191466 281636 191472 281648
rect 160888 281608 191472 281636
rect 160888 281596 160894 281608
rect 191466 281596 191472 281608
rect 191524 281596 191530 281648
rect 100846 281528 100852 281580
rect 100904 281568 100910 281580
rect 189902 281568 189908 281580
rect 100904 281540 189908 281568
rect 100904 281528 100910 281540
rect 189902 281528 189908 281540
rect 189960 281528 189966 281580
rect 99374 281460 99380 281512
rect 99432 281500 99438 281512
rect 140590 281500 140596 281512
rect 99432 281472 140596 281500
rect 99432 281460 99438 281472
rect 140590 281460 140596 281472
rect 140648 281500 140654 281512
rect 182818 281500 182824 281512
rect 140648 281472 182824 281500
rect 140648 281460 140654 281472
rect 182818 281460 182824 281472
rect 182876 281460 182882 281512
rect 255406 281460 255412 281512
rect 255464 281500 255470 281512
rect 292574 281500 292580 281512
rect 255464 281472 292580 281500
rect 255464 281460 255470 281472
rect 292574 281460 292580 281472
rect 292632 281460 292638 281512
rect 255498 281392 255504 281444
rect 255556 281432 255562 281444
rect 281718 281432 281724 281444
rect 255556 281404 281724 281432
rect 255556 281392 255562 281404
rect 281718 281392 281724 281404
rect 281776 281392 281782 281444
rect 126238 280848 126244 280900
rect 126296 280888 126302 280900
rect 137462 280888 137468 280900
rect 126296 280860 137468 280888
rect 126296 280848 126302 280860
rect 137462 280848 137468 280860
rect 137520 280848 137526 280900
rect 137278 280780 137284 280832
rect 137336 280820 137342 280832
rect 162118 280820 162124 280832
rect 137336 280792 162124 280820
rect 137336 280780 137342 280792
rect 162118 280780 162124 280792
rect 162176 280780 162182 280832
rect 163682 280780 163688 280832
rect 163740 280820 163746 280832
rect 173802 280820 173808 280832
rect 163740 280792 173808 280820
rect 163740 280780 163746 280792
rect 173802 280780 173808 280792
rect 173860 280820 173866 280832
rect 176010 280820 176016 280832
rect 173860 280792 176016 280820
rect 173860 280780 173866 280792
rect 176010 280780 176016 280792
rect 176068 280780 176074 280832
rect 179230 280780 179236 280832
rect 179288 280820 179294 280832
rect 191466 280820 191472 280832
rect 179288 280792 191472 280820
rect 179288 280780 179294 280792
rect 191466 280780 191472 280792
rect 191524 280780 191530 280832
rect 184290 280236 184296 280288
rect 184348 280276 184354 280288
rect 191466 280276 191472 280288
rect 184348 280248 191472 280276
rect 184348 280236 184354 280248
rect 191466 280236 191472 280248
rect 191524 280236 191530 280288
rect 43438 280168 43444 280220
rect 43496 280208 43502 280220
rect 67266 280208 67272 280220
rect 43496 280180 67272 280208
rect 43496 280168 43502 280180
rect 67266 280168 67272 280180
rect 67324 280168 67330 280220
rect 98730 280100 98736 280152
rect 98788 280140 98794 280152
rect 176194 280140 176200 280152
rect 98788 280112 176200 280140
rect 98788 280100 98794 280112
rect 176194 280100 176200 280112
rect 176252 280100 176258 280152
rect 263962 280100 263968 280152
rect 264020 280140 264026 280152
rect 264974 280140 264980 280152
rect 264020 280112 264980 280140
rect 264020 280100 264026 280112
rect 264974 280100 264980 280112
rect 265032 280100 265038 280152
rect 100754 280032 100760 280084
rect 100812 280072 100818 280084
rect 155310 280072 155316 280084
rect 100812 280044 155316 280072
rect 100812 280032 100818 280044
rect 155310 280032 155316 280044
rect 155368 280032 155374 280084
rect 163590 280032 163596 280084
rect 163648 280072 163654 280084
rect 164050 280072 164056 280084
rect 163648 280044 164056 280072
rect 163648 280032 163654 280044
rect 164050 280032 164056 280044
rect 164108 280032 164114 280084
rect 4062 279420 4068 279472
rect 4120 279460 4126 279472
rect 52454 279460 52460 279472
rect 4120 279432 52460 279460
rect 4120 279420 4126 279432
rect 52454 279420 52460 279432
rect 52512 279420 52518 279472
rect 164050 279420 164056 279472
rect 164108 279460 164114 279472
rect 191466 279460 191472 279472
rect 164108 279432 191472 279460
rect 164108 279420 164114 279432
rect 191466 279420 191472 279432
rect 191524 279420 191530 279472
rect 255406 279420 255412 279472
rect 255464 279460 255470 279472
rect 259270 279460 259276 279472
rect 255464 279432 259276 279460
rect 255464 279420 255470 279432
rect 259270 279420 259276 279432
rect 259328 279420 259334 279472
rect 52454 278740 52460 278792
rect 52512 278780 52518 278792
rect 53558 278780 53564 278792
rect 52512 278752 53564 278780
rect 52512 278740 52518 278752
rect 53558 278740 53564 278752
rect 53616 278780 53622 278792
rect 66806 278780 66812 278792
rect 53616 278752 66812 278780
rect 53616 278740 53622 278752
rect 66806 278740 66812 278752
rect 66864 278740 66870 278792
rect 53466 278672 53472 278724
rect 53524 278712 53530 278724
rect 67542 278712 67548 278724
rect 53524 278684 67548 278712
rect 53524 278672 53530 278684
rect 67542 278672 67548 278684
rect 67600 278672 67606 278724
rect 255498 278672 255504 278724
rect 255556 278712 255562 278724
rect 280154 278712 280160 278724
rect 255556 278684 280160 278712
rect 255556 278672 255562 278684
rect 280154 278672 280160 278684
rect 280212 278672 280218 278724
rect 258350 278604 258356 278656
rect 258408 278644 258414 278656
rect 262398 278644 262404 278656
rect 258408 278616 262404 278644
rect 258408 278604 258414 278616
rect 262398 278604 262404 278616
rect 262456 278604 262462 278656
rect 100846 278060 100852 278112
rect 100904 278100 100910 278112
rect 127710 278100 127716 278112
rect 100904 278072 127716 278100
rect 100904 278060 100910 278072
rect 127710 278060 127716 278072
rect 127768 278060 127774 278112
rect 105630 277992 105636 278044
rect 105688 278032 105694 278044
rect 156046 278032 156052 278044
rect 105688 278004 156052 278032
rect 105688 277992 105694 278004
rect 156046 277992 156052 278004
rect 156104 278032 156110 278044
rect 183462 278032 183468 278044
rect 156104 278004 183468 278032
rect 156104 277992 156110 278004
rect 183462 277992 183468 278004
rect 183520 277992 183526 278044
rect 255406 277992 255412 278044
rect 255464 278032 255470 278044
rect 258350 278032 258356 278044
rect 255464 278004 258356 278032
rect 255464 277992 255470 278004
rect 258350 277992 258356 278004
rect 258408 277992 258414 278044
rect 262858 277992 262864 278044
rect 262916 278032 262922 278044
rect 291378 278032 291384 278044
rect 262916 278004 291384 278032
rect 262916 277992 262922 278004
rect 291378 277992 291384 278004
rect 291436 278032 291442 278044
rect 580166 278032 580172 278044
rect 291436 278004 580172 278032
rect 291436 277992 291442 278004
rect 580166 277992 580172 278004
rect 580224 277992 580230 278044
rect 67266 277924 67272 277976
rect 67324 277964 67330 277976
rect 67542 277964 67548 277976
rect 67324 277936 67548 277964
rect 67324 277924 67330 277936
rect 67542 277924 67548 277936
rect 67600 277924 67606 277976
rect 183462 277380 183468 277432
rect 183520 277420 183526 277432
rect 191466 277420 191472 277432
rect 183520 277392 191472 277420
rect 183520 277380 183526 277392
rect 191466 277380 191472 277392
rect 191524 277380 191530 277432
rect 52270 277312 52276 277364
rect 52328 277352 52334 277364
rect 66898 277352 66904 277364
rect 52328 277324 66904 277352
rect 52328 277312 52334 277324
rect 66898 277312 66904 277324
rect 66956 277312 66962 277364
rect 100846 277312 100852 277364
rect 100904 277352 100910 277364
rect 154022 277352 154028 277364
rect 100904 277324 154028 277352
rect 100904 277312 100910 277324
rect 154022 277312 154028 277324
rect 154080 277312 154086 277364
rect 255406 277312 255412 277364
rect 255464 277352 255470 277364
rect 278866 277352 278872 277364
rect 255464 277324 278872 277352
rect 255464 277312 255470 277324
rect 278866 277312 278872 277324
rect 278924 277312 278930 277364
rect 100202 277244 100208 277296
rect 100260 277284 100266 277296
rect 150526 277284 150532 277296
rect 100260 277256 150532 277284
rect 100260 277244 100266 277256
rect 150526 277244 150532 277256
rect 150584 277284 150590 277296
rect 151262 277284 151268 277296
rect 150584 277256 151268 277284
rect 150584 277244 150590 277256
rect 151262 277244 151268 277256
rect 151320 277244 151326 277296
rect 155310 276632 155316 276684
rect 155368 276672 155374 276684
rect 177482 276672 177488 276684
rect 155368 276644 177488 276672
rect 155368 276632 155374 276644
rect 177482 276632 177488 276644
rect 177540 276632 177546 276684
rect 272334 276632 272340 276684
rect 272392 276672 272398 276684
rect 281810 276672 281816 276684
rect 272392 276644 281816 276672
rect 272392 276632 272398 276644
rect 281810 276632 281816 276644
rect 281868 276632 281874 276684
rect 66162 276020 66168 276072
rect 66220 276060 66226 276072
rect 67818 276060 67824 276072
rect 66220 276032 67824 276060
rect 66220 276020 66226 276032
rect 67818 276020 67824 276032
rect 67876 276020 67882 276072
rect 155494 276020 155500 276072
rect 155552 276060 155558 276072
rect 190638 276060 190644 276072
rect 155552 276032 190644 276060
rect 155552 276020 155558 276032
rect 190638 276020 190644 276032
rect 190696 276020 190702 276072
rect 255498 276020 255504 276072
rect 255556 276060 255562 276072
rect 271874 276060 271880 276072
rect 255556 276032 271880 276060
rect 255556 276020 255562 276032
rect 271874 276020 271880 276032
rect 271932 276060 271938 276072
rect 272334 276060 272340 276072
rect 271932 276032 272340 276060
rect 271932 276020 271938 276032
rect 272334 276020 272340 276032
rect 272392 276020 272398 276072
rect 255406 275952 255412 276004
rect 255464 275992 255470 276004
rect 277670 275992 277676 276004
rect 255464 275964 277676 275992
rect 255464 275952 255470 275964
rect 277670 275952 277676 275964
rect 277728 275952 277734 276004
rect 255498 275612 255504 275664
rect 255556 275652 255562 275664
rect 258074 275652 258080 275664
rect 255556 275624 258080 275652
rect 255556 275612 255562 275624
rect 258074 275612 258080 275624
rect 258132 275612 258138 275664
rect 155770 275340 155776 275392
rect 155828 275380 155834 275392
rect 177390 275380 177396 275392
rect 155828 275352 177396 275380
rect 155828 275340 155834 275352
rect 177390 275340 177396 275352
rect 177448 275340 177454 275392
rect 56226 275272 56232 275324
rect 56284 275312 56290 275324
rect 65702 275312 65708 275324
rect 56284 275284 65708 275312
rect 56284 275272 56290 275284
rect 65702 275272 65708 275284
rect 65760 275312 65766 275324
rect 66438 275312 66444 275324
rect 65760 275284 66444 275312
rect 65760 275272 65766 275284
rect 66438 275272 66444 275284
rect 66496 275272 66502 275324
rect 136542 275272 136548 275324
rect 136600 275312 136606 275324
rect 184198 275312 184204 275324
rect 136600 275284 184204 275312
rect 136600 275272 136606 275284
rect 184198 275272 184204 275284
rect 184256 275272 184262 275324
rect 188430 275000 188436 275052
rect 188488 275040 188494 275052
rect 191558 275040 191564 275052
rect 188488 275012 191564 275040
rect 188488 275000 188494 275012
rect 191558 275000 191564 275012
rect 191616 275000 191622 275052
rect 100938 274660 100944 274712
rect 100996 274700 101002 274712
rect 152826 274700 152832 274712
rect 100996 274672 152832 274700
rect 100996 274660 101002 274672
rect 152826 274660 152832 274672
rect 152884 274660 152890 274712
rect 100846 274592 100852 274644
rect 100904 274632 100910 274644
rect 120718 274632 120724 274644
rect 100904 274604 120724 274632
rect 100904 274592 100910 274604
rect 120718 274592 120724 274604
rect 120776 274592 120782 274644
rect 255498 274592 255504 274644
rect 255556 274632 255562 274644
rect 281626 274632 281632 274644
rect 255556 274604 281632 274632
rect 255556 274592 255562 274604
rect 281626 274592 281632 274604
rect 281684 274592 281690 274644
rect 156598 273980 156604 274032
rect 156656 274020 156662 274032
rect 188890 274020 188896 274032
rect 156656 273992 188896 274020
rect 156656 273980 156662 273992
rect 188890 273980 188896 273992
rect 188948 274020 188954 274032
rect 190822 274020 190828 274032
rect 188948 273992 190828 274020
rect 188948 273980 188954 273992
rect 190822 273980 190828 273992
rect 190880 273980 190886 274032
rect 100110 273912 100116 273964
rect 100168 273952 100174 273964
rect 120166 273952 120172 273964
rect 100168 273924 120172 273952
rect 100168 273912 100174 273924
rect 120166 273912 120172 273924
rect 120224 273912 120230 273964
rect 124950 273912 124956 273964
rect 125008 273952 125014 273964
rect 171778 273952 171784 273964
rect 125008 273924 171784 273952
rect 125008 273912 125014 273924
rect 171778 273912 171784 273924
rect 171836 273912 171842 273964
rect 255406 273912 255412 273964
rect 255464 273952 255470 273964
rect 260926 273952 260932 273964
rect 255464 273924 260932 273952
rect 255464 273912 255470 273924
rect 260926 273912 260932 273924
rect 260984 273912 260990 273964
rect 56502 273300 56508 273352
rect 56560 273340 56566 273352
rect 61102 273340 61108 273352
rect 56560 273312 61108 273340
rect 56560 273300 56566 273312
rect 61102 273300 61108 273312
rect 61160 273300 61166 273352
rect 64690 273232 64696 273284
rect 64748 273272 64754 273284
rect 66622 273272 66628 273284
rect 64748 273244 66628 273272
rect 64748 273232 64754 273244
rect 66622 273232 66628 273244
rect 66680 273232 66686 273284
rect 172330 273164 172336 273216
rect 172388 273204 172394 273216
rect 191558 273204 191564 273216
rect 172388 273176 191564 273204
rect 172388 273164 172394 273176
rect 191558 273164 191564 273176
rect 191616 273164 191622 273216
rect 255498 273164 255504 273216
rect 255556 273204 255562 273216
rect 261478 273204 261484 273216
rect 255556 273176 261484 273204
rect 255556 273164 255562 273176
rect 261478 273164 261484 273176
rect 261536 273164 261542 273216
rect 157978 272552 157984 272604
rect 158036 272592 158042 272604
rect 172330 272592 172336 272604
rect 158036 272564 172336 272592
rect 158036 272552 158042 272564
rect 172330 272552 172336 272564
rect 172388 272552 172394 272604
rect 48222 272484 48228 272536
rect 48280 272524 48286 272536
rect 59078 272524 59084 272536
rect 48280 272496 59084 272524
rect 48280 272484 48286 272496
rect 59078 272484 59084 272496
rect 59136 272484 59142 272536
rect 100846 272484 100852 272536
rect 100904 272524 100910 272536
rect 100904 272496 103514 272524
rect 100904 272484 100910 272496
rect 103486 271844 103514 272496
rect 118050 272484 118056 272536
rect 118108 272524 118114 272536
rect 174722 272524 174728 272536
rect 118108 272496 174728 272524
rect 118108 272484 118114 272496
rect 174722 272484 174728 272496
rect 174780 272484 174786 272536
rect 272058 272484 272064 272536
rect 272116 272524 272122 272536
rect 281626 272524 281632 272536
rect 272116 272496 281632 272524
rect 272116 272484 272122 272496
rect 281626 272484 281632 272496
rect 281684 272484 281690 272536
rect 113174 271872 113180 271924
rect 113232 271872 113238 271924
rect 113192 271844 113220 271872
rect 180150 271844 180156 271856
rect 103486 271816 180156 271844
rect 180150 271804 180156 271816
rect 180208 271804 180214 271856
rect 262398 271804 262404 271856
rect 262456 271844 262462 271856
rect 267826 271844 267832 271856
rect 262456 271816 267832 271844
rect 262456 271804 262462 271816
rect 267826 271804 267832 271816
rect 267884 271804 267890 271856
rect 49510 271124 49516 271176
rect 49568 271164 49574 271176
rect 65794 271164 65800 271176
rect 49568 271136 65800 271164
rect 49568 271124 49574 271136
rect 65794 271124 65800 271136
rect 65852 271164 65858 271176
rect 66530 271164 66536 271176
rect 65852 271136 66536 271164
rect 65852 271124 65858 271136
rect 66530 271124 66536 271136
rect 66588 271124 66594 271176
rect 147030 271124 147036 271176
rect 147088 271164 147094 271176
rect 180794 271164 180800 271176
rect 147088 271136 180800 271164
rect 147088 271124 147094 271136
rect 180794 271124 180800 271136
rect 180852 271164 180858 271176
rect 181714 271164 181720 271176
rect 180852 271136 181720 271164
rect 180852 271124 180858 271136
rect 181714 271124 181720 271136
rect 181772 271124 181778 271176
rect 255406 270784 255412 270836
rect 255464 270824 255470 270836
rect 259362 270824 259368 270836
rect 255464 270796 259368 270824
rect 255464 270784 255470 270796
rect 259362 270784 259368 270796
rect 259420 270784 259426 270836
rect 181714 270512 181720 270564
rect 181772 270552 181778 270564
rect 191558 270552 191564 270564
rect 181772 270524 191564 270552
rect 181772 270512 181778 270524
rect 191558 270512 191564 270524
rect 191616 270512 191622 270564
rect 57606 270444 57612 270496
rect 57664 270484 57670 270496
rect 57882 270484 57888 270496
rect 57664 270456 57888 270484
rect 57664 270444 57670 270456
rect 57882 270444 57888 270456
rect 57940 270484 57946 270496
rect 66806 270484 66812 270496
rect 57940 270456 66812 270484
rect 57940 270444 57946 270456
rect 66806 270444 66812 270456
rect 66864 270444 66870 270496
rect 100846 270444 100852 270496
rect 100904 270484 100910 270496
rect 114554 270484 114560 270496
rect 100904 270456 114560 270484
rect 100904 270444 100910 270456
rect 114554 270444 114560 270456
rect 114612 270484 114618 270496
rect 119338 270484 119344 270496
rect 114612 270456 119344 270484
rect 114612 270444 114618 270456
rect 119338 270444 119344 270456
rect 119396 270444 119402 270496
rect 255406 270444 255412 270496
rect 255464 270484 255470 270496
rect 280338 270484 280344 270496
rect 255464 270456 280344 270484
rect 255464 270444 255470 270456
rect 280338 270444 280344 270456
rect 280396 270444 280402 270496
rect 154022 269832 154028 269884
rect 154080 269872 154086 269884
rect 169110 269872 169116 269884
rect 154080 269844 169116 269872
rect 154080 269832 154086 269844
rect 169110 269832 169116 269844
rect 169168 269832 169174 269884
rect 43990 269764 43996 269816
rect 44048 269804 44054 269816
rect 57882 269804 57888 269816
rect 44048 269776 57888 269804
rect 44048 269764 44054 269776
rect 57882 269764 57888 269776
rect 57940 269764 57946 269816
rect 98822 269764 98828 269816
rect 98880 269804 98886 269816
rect 165062 269804 165068 269816
rect 98880 269776 165068 269804
rect 98880 269764 98886 269776
rect 165062 269764 165068 269776
rect 165120 269764 165126 269816
rect 259362 269764 259368 269816
rect 259420 269804 259426 269816
rect 280338 269804 280344 269816
rect 259420 269776 280344 269804
rect 259420 269764 259426 269776
rect 280338 269764 280344 269776
rect 280396 269764 280402 269816
rect 184198 269356 184204 269408
rect 184256 269396 184262 269408
rect 191558 269396 191564 269408
rect 184256 269368 191564 269396
rect 184256 269356 184262 269368
rect 191558 269356 191564 269368
rect 191616 269356 191622 269408
rect 181990 269016 181996 269068
rect 182048 269056 182054 269068
rect 191558 269056 191564 269068
rect 182048 269028 191564 269056
rect 182048 269016 182054 269028
rect 191558 269016 191564 269028
rect 191616 269016 191622 269068
rect 141418 268404 141424 268456
rect 141476 268444 141482 268456
rect 181990 268444 181996 268456
rect 141476 268416 181996 268444
rect 141476 268404 141482 268416
rect 181990 268404 181996 268416
rect 182048 268404 182054 268456
rect 57790 268336 57796 268388
rect 57848 268376 57854 268388
rect 59262 268376 59268 268388
rect 57848 268348 59268 268376
rect 57848 268336 57854 268348
rect 59262 268336 59268 268348
rect 59320 268376 59326 268388
rect 66806 268376 66812 268388
rect 59320 268348 66812 268376
rect 59320 268336 59326 268348
rect 66806 268336 66812 268348
rect 66864 268336 66870 268388
rect 104158 268336 104164 268388
rect 104216 268376 104222 268388
rect 163498 268376 163504 268388
rect 104216 268348 163504 268376
rect 104216 268336 104222 268348
rect 163498 268336 163504 268348
rect 163556 268336 163562 268388
rect 168282 268336 168288 268388
rect 168340 268376 168346 268388
rect 176654 268376 176660 268388
rect 168340 268348 176660 268376
rect 168340 268336 168346 268348
rect 176654 268336 176660 268348
rect 176712 268336 176718 268388
rect 269022 268336 269028 268388
rect 269080 268376 269086 268388
rect 280430 268376 280436 268388
rect 269080 268348 280436 268376
rect 269080 268336 269086 268348
rect 280430 268336 280436 268348
rect 280488 268336 280494 268388
rect 104802 268200 104808 268252
rect 104860 268240 104866 268252
rect 105538 268240 105544 268252
rect 104860 268212 105544 268240
rect 104860 268200 104866 268212
rect 105538 268200 105544 268212
rect 105596 268200 105602 268252
rect 255406 267792 255412 267844
rect 255464 267832 255470 267844
rect 268102 267832 268108 267844
rect 255464 267804 268108 267832
rect 255464 267792 255470 267804
rect 268102 267792 268108 267804
rect 268160 267832 268166 267844
rect 269022 267832 269028 267844
rect 268160 267804 269028 267832
rect 268160 267792 268166 267804
rect 269022 267792 269028 267804
rect 269080 267792 269086 267844
rect 100846 267724 100852 267776
rect 100904 267764 100910 267776
rect 104802 267764 104808 267776
rect 100904 267736 104808 267764
rect 100904 267724 100910 267736
rect 104802 267724 104808 267736
rect 104860 267724 104866 267776
rect 255498 267724 255504 267776
rect 255556 267764 255562 267776
rect 269390 267764 269396 267776
rect 255556 267736 269396 267764
rect 255556 267724 255562 267736
rect 269390 267724 269396 267736
rect 269448 267724 269454 267776
rect 100018 267656 100024 267708
rect 100076 267696 100082 267708
rect 135162 267696 135168 267708
rect 100076 267668 135168 267696
rect 100076 267656 100082 267668
rect 135162 267656 135168 267668
rect 135220 267656 135226 267708
rect 255406 267656 255412 267708
rect 255464 267696 255470 267708
rect 267918 267696 267924 267708
rect 255464 267668 267924 267696
rect 255464 267656 255470 267668
rect 267918 267656 267924 267668
rect 267976 267656 267982 267708
rect 282914 267112 282920 267164
rect 282972 267152 282978 267164
rect 284478 267152 284484 267164
rect 282972 267124 284484 267152
rect 282972 267112 282978 267124
rect 284478 267112 284484 267124
rect 284536 267112 284542 267164
rect 54938 267044 54944 267096
rect 54996 267084 55002 267096
rect 65978 267084 65984 267096
rect 54996 267056 65984 267084
rect 54996 267044 55002 267056
rect 65978 267044 65984 267056
rect 66036 267044 66042 267096
rect 135162 267044 135168 267096
rect 135220 267084 135226 267096
rect 169110 267084 169116 267096
rect 135220 267056 169116 267084
rect 135220 267044 135226 267056
rect 169110 267044 169116 267056
rect 169168 267044 169174 267096
rect 44082 266976 44088 267028
rect 44140 267016 44146 267028
rect 58342 267016 58348 267028
rect 44140 266988 58348 267016
rect 44140 266976 44146 266988
rect 58342 266976 58348 266988
rect 58400 266976 58406 267028
rect 101398 266976 101404 267028
rect 101456 267016 101462 267028
rect 141694 267016 141700 267028
rect 101456 266988 141700 267016
rect 101456 266976 101462 266988
rect 141694 266976 141700 266988
rect 141752 266976 141758 267028
rect 166442 266976 166448 267028
rect 166500 267016 166506 267028
rect 174630 267016 174636 267028
rect 166500 266988 174636 267016
rect 166500 266976 166506 266988
rect 174630 266976 174636 266988
rect 174688 266976 174694 267028
rect 186130 266976 186136 267028
rect 186188 267016 186194 267028
rect 192570 267016 192576 267028
rect 186188 266988 192576 267016
rect 186188 266976 186194 266988
rect 192570 266976 192576 266988
rect 192628 266976 192634 267028
rect 259362 266364 259368 266416
rect 259420 266404 259426 266416
rect 282914 266404 282920 266416
rect 259420 266376 282920 266404
rect 259420 266364 259426 266376
rect 282914 266364 282920 266376
rect 282972 266364 282978 266416
rect 111794 266296 111800 266348
rect 111852 266336 111858 266348
rect 113082 266336 113088 266348
rect 111852 266308 113088 266336
rect 111852 266296 111858 266308
rect 113082 266296 113088 266308
rect 113140 266336 113146 266348
rect 160830 266336 160836 266348
rect 113140 266308 160836 266336
rect 113140 266296 113146 266308
rect 160830 266296 160836 266308
rect 160888 266296 160894 266348
rect 168190 266296 168196 266348
rect 168248 266336 168254 266348
rect 191650 266336 191656 266348
rect 168248 266308 191656 266336
rect 168248 266296 168254 266308
rect 191650 266296 191656 266308
rect 191708 266296 191714 266348
rect 255406 266160 255412 266212
rect 255464 266200 255470 266212
rect 260098 266200 260104 266212
rect 255464 266172 260104 266200
rect 255464 266160 255470 266172
rect 260098 266160 260104 266172
rect 260156 266160 260162 266212
rect 101122 265616 101128 265668
rect 101180 265656 101186 265668
rect 111794 265656 111800 265668
rect 101180 265628 111800 265656
rect 101180 265616 101186 265628
rect 111794 265616 111800 265628
rect 111852 265616 111858 265668
rect 153930 265616 153936 265668
rect 153988 265656 153994 265668
rect 184934 265656 184940 265668
rect 153988 265628 184940 265656
rect 153988 265616 153994 265628
rect 184934 265616 184940 265628
rect 184992 265656 184998 265668
rect 190638 265656 190644 265668
rect 184992 265628 190644 265656
rect 184992 265616 184998 265628
rect 190638 265616 190644 265628
rect 190696 265616 190702 265668
rect 63126 264936 63132 264988
rect 63184 264976 63190 264988
rect 66806 264976 66812 264988
rect 63184 264948 66812 264976
rect 63184 264936 63190 264948
rect 66806 264936 66812 264948
rect 66864 264936 66870 264988
rect 100846 264936 100852 264988
rect 100904 264976 100910 264988
rect 133230 264976 133236 264988
rect 100904 264948 133236 264976
rect 100904 264936 100910 264948
rect 133230 264936 133236 264948
rect 133288 264936 133294 264988
rect 164970 264936 164976 264988
rect 165028 264976 165034 264988
rect 168190 264976 168196 264988
rect 165028 264948 168196 264976
rect 165028 264936 165034 264948
rect 168190 264936 168196 264948
rect 168248 264936 168254 264988
rect 255314 264936 255320 264988
rect 255372 264976 255378 264988
rect 295426 264976 295432 264988
rect 255372 264948 295432 264976
rect 255372 264936 255378 264948
rect 295426 264936 295432 264948
rect 295484 264936 295490 264988
rect 137462 264256 137468 264308
rect 137520 264296 137526 264308
rect 169202 264296 169208 264308
rect 137520 264268 169208 264296
rect 137520 264256 137526 264268
rect 169202 264256 169208 264268
rect 169260 264256 169266 264308
rect 98730 264188 98736 264240
rect 98788 264228 98794 264240
rect 153930 264228 153936 264240
rect 98788 264200 153936 264228
rect 98788 264188 98794 264200
rect 153930 264188 153936 264200
rect 153988 264188 153994 264240
rect 276014 264188 276020 264240
rect 276072 264228 276078 264240
rect 285766 264228 285772 264240
rect 276072 264200 285772 264228
rect 276072 264188 276078 264200
rect 285766 264188 285772 264200
rect 285824 264188 285830 264240
rect 255406 264120 255412 264172
rect 255464 264160 255470 264172
rect 259362 264160 259368 264172
rect 255464 264132 259368 264160
rect 255464 264120 255470 264132
rect 259362 264120 259368 264132
rect 259420 264120 259426 264172
rect 255498 263712 255504 263764
rect 255556 263752 255562 263764
rect 259730 263752 259736 263764
rect 255556 263724 259736 263752
rect 255556 263712 255562 263724
rect 259730 263712 259736 263724
rect 259788 263712 259794 263764
rect 59262 263576 59268 263628
rect 59320 263616 59326 263628
rect 63218 263616 63224 263628
rect 59320 263588 63224 263616
rect 59320 263576 59326 263588
rect 63218 263576 63224 263588
rect 63276 263616 63282 263628
rect 66622 263616 66628 263628
rect 63276 263588 66628 263616
rect 63276 263576 63282 263588
rect 66622 263576 66628 263588
rect 66680 263576 66686 263628
rect 100938 263576 100944 263628
rect 100996 263616 101002 263628
rect 120718 263616 120724 263628
rect 100996 263588 120724 263616
rect 100996 263576 101002 263588
rect 120718 263576 120724 263588
rect 120776 263576 120782 263628
rect 160830 263576 160836 263628
rect 160888 263616 160894 263628
rect 192018 263616 192024 263628
rect 160888 263588 192024 263616
rect 160888 263576 160894 263588
rect 192018 263576 192024 263588
rect 192076 263576 192082 263628
rect 260742 263576 260748 263628
rect 260800 263616 260806 263628
rect 287238 263616 287244 263628
rect 260800 263588 287244 263616
rect 260800 263576 260806 263588
rect 287238 263576 287244 263588
rect 287296 263576 287302 263628
rect 100846 263508 100852 263560
rect 100904 263548 100910 263560
rect 141602 263548 141608 263560
rect 100904 263520 141608 263548
rect 100904 263508 100910 263520
rect 141602 263508 141608 263520
rect 141660 263508 141666 263560
rect 142890 262964 142896 263016
rect 142948 263004 142954 263016
rect 152734 263004 152740 263016
rect 142948 262976 152740 263004
rect 142948 262964 142954 262976
rect 152734 262964 152740 262976
rect 152792 262964 152798 263016
rect 152550 262896 152556 262948
rect 152608 262936 152614 262948
rect 172514 262936 172520 262948
rect 152608 262908 172520 262936
rect 152608 262896 152614 262908
rect 172514 262896 172520 262908
rect 172572 262896 172578 262948
rect 54846 262828 54852 262880
rect 54904 262868 54910 262880
rect 66254 262868 66260 262880
rect 54904 262840 66260 262868
rect 54904 262828 54910 262840
rect 66254 262828 66260 262840
rect 66312 262828 66318 262880
rect 141510 262828 141516 262880
rect 141568 262868 141574 262880
rect 179414 262868 179420 262880
rect 141568 262840 179420 262868
rect 141568 262828 141574 262840
rect 179414 262828 179420 262840
rect 179472 262828 179478 262880
rect 255498 262284 255504 262336
rect 255556 262324 255562 262336
rect 263870 262324 263876 262336
rect 255556 262296 263876 262324
rect 255556 262284 255562 262296
rect 263870 262284 263876 262296
rect 263928 262284 263934 262336
rect 22738 262216 22744 262268
rect 22796 262256 22802 262268
rect 63218 262256 63224 262268
rect 22796 262228 63224 262256
rect 22796 262216 22802 262228
rect 63218 262216 63224 262228
rect 63276 262256 63282 262268
rect 66898 262256 66904 262268
rect 63276 262228 66904 262256
rect 63276 262216 63282 262228
rect 66898 262216 66904 262228
rect 66956 262216 66962 262268
rect 179414 262216 179420 262268
rect 179472 262256 179478 262268
rect 191650 262256 191656 262268
rect 179472 262228 191656 262256
rect 179472 262216 179478 262228
rect 191650 262216 191656 262228
rect 191708 262216 191714 262268
rect 255406 262216 255412 262268
rect 255464 262256 255470 262268
rect 267826 262256 267832 262268
rect 255464 262228 267832 262256
rect 255464 262216 255470 262228
rect 267826 262216 267832 262228
rect 267884 262256 267890 262268
rect 268286 262256 268292 262268
rect 267884 262228 268292 262256
rect 267884 262216 267890 262228
rect 268286 262216 268292 262228
rect 268344 262216 268350 262268
rect 164142 262148 164148 262200
rect 164200 262188 164206 262200
rect 168374 262188 168380 262200
rect 164200 262160 168380 262188
rect 164200 262148 164206 262160
rect 168374 262148 168380 262160
rect 168432 262148 168438 262200
rect 104802 262080 104808 262132
rect 104860 262120 104866 262132
rect 111058 262120 111064 262132
rect 104860 262092 111064 262120
rect 104860 262080 104866 262092
rect 111058 262080 111064 262092
rect 111116 262080 111122 262132
rect 7558 261468 7564 261520
rect 7616 261508 7622 261520
rect 67082 261508 67088 261520
rect 7616 261480 67088 261508
rect 7616 261468 7622 261480
rect 67082 261468 67088 261480
rect 67140 261468 67146 261520
rect 100846 261468 100852 261520
rect 100904 261508 100910 261520
rect 104618 261508 104624 261520
rect 100904 261480 104624 261508
rect 100904 261468 100910 261480
rect 104618 261468 104624 261480
rect 104676 261508 104682 261520
rect 134610 261508 134616 261520
rect 104676 261480 134616 261508
rect 104676 261468 104682 261480
rect 134610 261468 134616 261480
rect 134668 261468 134674 261520
rect 141510 261468 141516 261520
rect 141568 261508 141574 261520
rect 167086 261508 167092 261520
rect 141568 261480 167092 261508
rect 141568 261468 141574 261480
rect 167086 261468 167092 261480
rect 167144 261468 167150 261520
rect 255498 261468 255504 261520
rect 255556 261508 255562 261520
rect 276014 261508 276020 261520
rect 255556 261480 276020 261508
rect 255556 261468 255562 261480
rect 276014 261468 276020 261480
rect 276072 261468 276078 261520
rect 255406 261332 255412 261384
rect 255464 261372 255470 261384
rect 259362 261372 259368 261384
rect 255464 261344 259368 261372
rect 255464 261332 255470 261344
rect 259362 261332 259368 261344
rect 259420 261332 259426 261384
rect 168374 260856 168380 260908
rect 168432 260896 168438 260908
rect 191650 260896 191656 260908
rect 168432 260868 191656 260896
rect 168432 260856 168438 260868
rect 191650 260856 191656 260868
rect 191708 260856 191714 260908
rect 255406 260448 255412 260500
rect 255464 260488 255470 260500
rect 260742 260488 260748 260500
rect 255464 260460 260748 260488
rect 255464 260448 255470 260460
rect 260742 260448 260748 260460
rect 260800 260448 260806 260500
rect 169294 260176 169300 260228
rect 169352 260216 169358 260228
rect 191374 260216 191380 260228
rect 169352 260188 191380 260216
rect 169352 260176 169358 260188
rect 191374 260176 191380 260188
rect 191432 260176 191438 260228
rect 55030 260108 55036 260160
rect 55088 260148 55094 260160
rect 66254 260148 66260 260160
rect 55088 260120 66260 260148
rect 55088 260108 55094 260120
rect 66254 260108 66260 260120
rect 66312 260108 66318 260160
rect 129274 260108 129280 260160
rect 129332 260148 129338 260160
rect 170490 260148 170496 260160
rect 129332 260120 170496 260148
rect 129332 260108 129338 260120
rect 170490 260108 170496 260120
rect 170548 260108 170554 260160
rect 259362 260108 259368 260160
rect 259420 260148 259426 260160
rect 278958 260148 278964 260160
rect 259420 260120 278964 260148
rect 259420 260108 259426 260120
rect 278958 260108 278964 260120
rect 279016 260108 279022 260160
rect 48222 259428 48228 259480
rect 48280 259468 48286 259480
rect 67726 259468 67732 259480
rect 48280 259440 67732 259468
rect 48280 259428 48286 259440
rect 67726 259428 67732 259440
rect 67784 259428 67790 259480
rect 100846 259428 100852 259480
rect 100904 259468 100910 259480
rect 149882 259468 149888 259480
rect 100904 259440 149888 259468
rect 100904 259428 100910 259440
rect 149882 259428 149888 259440
rect 149940 259428 149946 259480
rect 176654 259428 176660 259480
rect 176712 259468 176718 259480
rect 191650 259468 191656 259480
rect 176712 259440 191656 259468
rect 176712 259428 176718 259440
rect 191650 259428 191656 259440
rect 191708 259428 191714 259480
rect 285766 259428 285772 259480
rect 285824 259468 285830 259480
rect 287330 259468 287336 259480
rect 285824 259440 287336 259468
rect 285824 259428 285830 259440
rect 287330 259428 287336 259440
rect 287388 259428 287394 259480
rect 64598 259360 64604 259412
rect 64656 259400 64662 259412
rect 66806 259400 66812 259412
rect 64656 259372 66812 259400
rect 64656 259360 64662 259372
rect 66806 259360 66812 259372
rect 66864 259360 66870 259412
rect 255406 259360 255412 259412
rect 255464 259400 255470 259412
rect 265158 259400 265164 259412
rect 255464 259372 265164 259400
rect 255464 259360 255470 259372
rect 265158 259360 265164 259372
rect 265216 259360 265222 259412
rect 273898 259360 273904 259412
rect 273956 259400 273962 259412
rect 274726 259400 274732 259412
rect 273956 259372 274732 259400
rect 273956 259360 273962 259372
rect 274726 259360 274732 259372
rect 274784 259360 274790 259412
rect 186314 259088 186320 259140
rect 186372 259128 186378 259140
rect 187142 259128 187148 259140
rect 186372 259100 187148 259128
rect 186372 259088 186378 259100
rect 187142 259088 187148 259100
rect 187200 259088 187206 259140
rect 52178 258680 52184 258732
rect 52236 258720 52242 258732
rect 61746 258720 61752 258732
rect 52236 258692 61752 258720
rect 52236 258680 52242 258692
rect 61746 258680 61752 258692
rect 61804 258720 61810 258732
rect 66254 258720 66260 258732
rect 61804 258692 66260 258720
rect 61804 258680 61810 258692
rect 66254 258680 66260 258692
rect 66312 258680 66318 258732
rect 98362 258136 98368 258188
rect 98420 258176 98426 258188
rect 113910 258176 113916 258188
rect 98420 258148 113916 258176
rect 98420 258136 98426 258148
rect 113910 258136 113916 258148
rect 113968 258136 113974 258188
rect 171134 258136 171140 258188
rect 171192 258176 171198 258188
rect 190454 258176 190460 258188
rect 171192 258148 190460 258176
rect 171192 258136 171198 258148
rect 190454 258136 190460 258148
rect 190512 258136 190518 258188
rect 108482 258068 108488 258120
rect 108540 258108 108546 258120
rect 187142 258108 187148 258120
rect 108540 258080 187148 258108
rect 108540 258068 108546 258080
rect 187142 258068 187148 258080
rect 187200 258068 187206 258120
rect 66254 258000 66260 258052
rect 66312 258040 66318 258052
rect 68186 258040 68192 258052
rect 66312 258012 68192 258040
rect 66312 258000 66318 258012
rect 68186 258000 68192 258012
rect 68244 258000 68250 258052
rect 255406 258000 255412 258052
rect 255464 258040 255470 258052
rect 261478 258040 261484 258052
rect 255464 258012 261484 258040
rect 255464 258000 255470 258012
rect 261478 258000 261484 258012
rect 261536 258000 261542 258052
rect 39850 257320 39856 257372
rect 39908 257360 39914 257372
rect 52454 257360 52460 257372
rect 39908 257332 52460 257360
rect 39908 257320 39914 257332
rect 52454 257320 52460 257332
rect 52512 257320 52518 257372
rect 101950 257320 101956 257372
rect 102008 257360 102014 257372
rect 112714 257360 112720 257372
rect 102008 257332 112720 257360
rect 102008 257320 102014 257332
rect 112714 257320 112720 257332
rect 112772 257320 112778 257372
rect 169018 257320 169024 257372
rect 169076 257360 169082 257372
rect 185486 257360 185492 257372
rect 169076 257332 185492 257360
rect 169076 257320 169082 257332
rect 185486 257320 185492 257332
rect 185544 257320 185550 257372
rect 255314 257320 255320 257372
rect 255372 257360 255378 257372
rect 256970 257360 256976 257372
rect 255372 257332 256976 257360
rect 255372 257320 255378 257332
rect 256970 257320 256976 257332
rect 257028 257320 257034 257372
rect 259546 257320 259552 257372
rect 259604 257360 259610 257372
rect 580902 257360 580908 257372
rect 259604 257332 580908 257360
rect 259604 257320 259610 257332
rect 580902 257320 580908 257332
rect 580960 257320 580966 257372
rect 185578 257184 185584 257236
rect 185636 257224 185642 257236
rect 190638 257224 190644 257236
rect 185636 257196 190644 257224
rect 185636 257184 185642 257196
rect 190638 257184 190644 257196
rect 190696 257184 190702 257236
rect 52454 256708 52460 256760
rect 52512 256748 52518 256760
rect 53466 256748 53472 256760
rect 52512 256720 53472 256748
rect 52512 256708 52518 256720
rect 53466 256708 53472 256720
rect 53524 256748 53530 256760
rect 66254 256748 66260 256760
rect 53524 256720 66260 256748
rect 53524 256708 53530 256720
rect 66254 256708 66260 256720
rect 66312 256708 66318 256760
rect 125042 256708 125048 256760
rect 125100 256748 125106 256760
rect 187050 256748 187056 256760
rect 125100 256720 187056 256748
rect 125100 256708 125106 256720
rect 187050 256708 187056 256720
rect 187108 256708 187114 256760
rect 100846 256640 100852 256692
rect 100904 256680 100910 256692
rect 143074 256680 143080 256692
rect 100904 256652 143080 256680
rect 100904 256640 100910 256652
rect 143074 256640 143080 256652
rect 143132 256640 143138 256692
rect 180242 256164 180248 256216
rect 180300 256204 180306 256216
rect 182818 256204 182824 256216
rect 180300 256176 182824 256204
rect 180300 256164 180306 256176
rect 182818 256164 182824 256176
rect 182876 256164 182882 256216
rect 166902 256028 166908 256080
rect 166960 256068 166966 256080
rect 173894 256068 173900 256080
rect 166960 256040 173900 256068
rect 166960 256028 166966 256040
rect 173894 256028 173900 256040
rect 173952 256028 173958 256080
rect 50890 255960 50896 256012
rect 50948 256000 50954 256012
rect 56502 256000 56508 256012
rect 50948 255972 56508 256000
rect 50948 255960 50954 255972
rect 56502 255960 56508 255972
rect 56560 255960 56566 256012
rect 147030 255960 147036 256012
rect 147088 256000 147094 256012
rect 170398 256000 170404 256012
rect 147088 255972 170404 256000
rect 147088 255960 147094 255972
rect 170398 255960 170404 255972
rect 170456 255960 170462 256012
rect 175182 255960 175188 256012
rect 175240 256000 175246 256012
rect 191650 256000 191656 256012
rect 175240 255972 191656 256000
rect 175240 255960 175246 255972
rect 191650 255960 191656 255972
rect 191708 255960 191714 256012
rect 255498 255348 255504 255400
rect 255556 255388 255562 255400
rect 265066 255388 265072 255400
rect 255556 255360 265072 255388
rect 255556 255348 255562 255360
rect 265066 255348 265072 255360
rect 265124 255348 265130 255400
rect 100938 255280 100944 255332
rect 100996 255320 101002 255332
rect 148502 255320 148508 255332
rect 100996 255292 148508 255320
rect 100996 255280 101002 255292
rect 148502 255280 148508 255292
rect 148560 255280 148566 255332
rect 255406 255280 255412 255332
rect 255464 255320 255470 255332
rect 274910 255320 274916 255332
rect 255464 255292 274916 255320
rect 255464 255280 255470 255292
rect 274910 255280 274916 255292
rect 274968 255280 274974 255332
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 43438 255252 43444 255264
rect 3476 255224 43444 255252
rect 3476 255212 3482 255224
rect 43438 255212 43444 255224
rect 43496 255212 43502 255264
rect 100846 255212 100852 255264
rect 100904 255252 100910 255264
rect 108942 255252 108948 255264
rect 100904 255224 108948 255252
rect 100904 255212 100910 255224
rect 108942 255212 108948 255224
rect 109000 255252 109006 255264
rect 109000 255224 113174 255252
rect 109000 255212 109006 255224
rect 113146 255184 113174 255224
rect 177758 255212 177764 255264
rect 177816 255252 177822 255264
rect 191006 255252 191012 255264
rect 177816 255224 191012 255252
rect 177816 255212 177822 255224
rect 191006 255212 191012 255224
rect 191064 255212 191070 255264
rect 114646 255184 114652 255196
rect 113146 255156 114652 255184
rect 114646 255144 114652 255156
rect 114704 255144 114710 255196
rect 272334 254600 272340 254652
rect 272392 254640 272398 254652
rect 283190 254640 283196 254652
rect 272392 254612 283196 254640
rect 272392 254600 272398 254612
rect 283190 254600 283196 254612
rect 283248 254600 283254 254652
rect 48130 254532 48136 254584
rect 48188 254572 48194 254584
rect 66806 254572 66812 254584
rect 48188 254544 66812 254572
rect 48188 254532 48194 254544
rect 66806 254532 66812 254544
rect 66864 254532 66870 254584
rect 120718 254532 120724 254584
rect 120776 254572 120782 254584
rect 184382 254572 184388 254584
rect 120776 254544 184388 254572
rect 120776 254532 120782 254544
rect 184382 254532 184388 254544
rect 184440 254532 184446 254584
rect 255406 254532 255412 254584
rect 255464 254572 255470 254584
rect 285766 254572 285772 254584
rect 255464 254544 285772 254572
rect 255464 254532 255470 254544
rect 285766 254532 285772 254544
rect 285824 254532 285830 254584
rect 108390 253920 108396 253972
rect 108448 253960 108454 253972
rect 109678 253960 109684 253972
rect 108448 253932 109684 253960
rect 108448 253920 108454 253932
rect 109678 253920 109684 253932
rect 109736 253920 109742 253972
rect 109862 253920 109868 253972
rect 109920 253960 109926 253972
rect 112438 253960 112444 253972
rect 109920 253932 112444 253960
rect 109920 253920 109926 253932
rect 112438 253920 112444 253932
rect 112496 253920 112502 253972
rect 255498 253920 255504 253972
rect 255556 253960 255562 253972
rect 272058 253960 272064 253972
rect 255556 253932 272064 253960
rect 255556 253920 255562 253932
rect 272058 253920 272064 253932
rect 272116 253960 272122 253972
rect 272334 253960 272340 253972
rect 272116 253932 272340 253960
rect 272116 253920 272122 253932
rect 272334 253920 272340 253932
rect 272392 253920 272398 253972
rect 111794 253240 111800 253292
rect 111852 253280 111858 253292
rect 147122 253280 147128 253292
rect 111852 253252 147128 253280
rect 111852 253240 111858 253252
rect 147122 253240 147128 253252
rect 147180 253240 147186 253292
rect 35158 253172 35164 253224
rect 35216 253212 35222 253224
rect 66990 253212 66996 253224
rect 35216 253184 66996 253212
rect 35216 253172 35222 253184
rect 66990 253172 66996 253184
rect 67048 253212 67054 253224
rect 67266 253212 67272 253224
rect 67048 253184 67272 253212
rect 67048 253172 67054 253184
rect 67266 253172 67272 253184
rect 67324 253172 67330 253224
rect 116670 253172 116676 253224
rect 116728 253212 116734 253224
rect 176010 253212 176016 253224
rect 116728 253184 176016 253212
rect 116728 253172 116734 253184
rect 176010 253172 176016 253184
rect 176068 253172 176074 253224
rect 188890 252968 188896 253020
rect 188948 253008 188954 253020
rect 189718 253008 189724 253020
rect 188948 252980 189724 253008
rect 188948 252968 188954 252980
rect 189718 252968 189724 252980
rect 189776 252968 189782 253020
rect 279326 252764 279332 252816
rect 279384 252804 279390 252816
rect 284386 252804 284392 252816
rect 279384 252776 284392 252804
rect 279384 252764 279390 252776
rect 284386 252764 284392 252776
rect 284444 252764 284450 252816
rect 255406 252696 255412 252748
rect 255464 252736 255470 252748
rect 258258 252736 258264 252748
rect 255464 252708 258264 252736
rect 255464 252696 255470 252708
rect 258258 252696 258264 252708
rect 258316 252696 258322 252748
rect 100846 252560 100852 252612
rect 100904 252600 100910 252612
rect 109678 252600 109684 252612
rect 100904 252572 109684 252600
rect 100904 252560 100910 252572
rect 109678 252560 109684 252572
rect 109736 252560 109742 252612
rect 163498 252560 163504 252612
rect 163556 252600 163562 252612
rect 188890 252600 188896 252612
rect 163556 252572 188896 252600
rect 163556 252560 163562 252572
rect 188890 252560 188896 252572
rect 188948 252560 188954 252612
rect 255498 252560 255504 252612
rect 255556 252600 255562 252612
rect 283098 252600 283104 252612
rect 255556 252572 283104 252600
rect 255556 252560 255562 252572
rect 283098 252560 283104 252572
rect 283156 252560 283162 252612
rect 186038 252492 186044 252544
rect 186096 252532 186102 252544
rect 191098 252532 191104 252544
rect 186096 252504 191104 252532
rect 186096 252492 186102 252504
rect 191098 252492 191104 252504
rect 191156 252492 191162 252544
rect 166258 251880 166264 251932
rect 166316 251920 166322 251932
rect 191006 251920 191012 251932
rect 166316 251892 191012 251920
rect 166316 251880 166322 251892
rect 191006 251880 191012 251892
rect 191064 251880 191070 251932
rect 54754 251812 54760 251864
rect 54812 251852 54818 251864
rect 63494 251852 63500 251864
rect 54812 251824 63500 251852
rect 54812 251812 54818 251824
rect 63494 251812 63500 251824
rect 63552 251812 63558 251864
rect 132034 251812 132040 251864
rect 132092 251852 132098 251864
rect 166350 251852 166356 251864
rect 132092 251824 166356 251852
rect 132092 251812 132098 251824
rect 166350 251812 166356 251824
rect 166408 251812 166414 251864
rect 255406 251812 255412 251864
rect 255464 251852 255470 251864
rect 278866 251852 278872 251864
rect 255464 251824 278872 251852
rect 255464 251812 255470 251824
rect 278866 251812 278872 251824
rect 278924 251852 278930 251864
rect 279326 251852 279332 251864
rect 278924 251824 279332 251852
rect 278924 251812 278930 251824
rect 279326 251812 279332 251824
rect 279384 251812 279390 251864
rect 291102 251812 291108 251864
rect 291160 251852 291166 251864
rect 299566 251852 299572 251864
rect 291160 251824 299572 251852
rect 291160 251812 291166 251824
rect 299566 251812 299572 251824
rect 299624 251812 299630 251864
rect 104250 251744 104256 251796
rect 104308 251784 104314 251796
rect 104802 251784 104808 251796
rect 104308 251756 104808 251784
rect 104308 251744 104314 251756
rect 104802 251744 104808 251756
rect 104860 251744 104866 251796
rect 63494 251268 63500 251320
rect 63552 251308 63558 251320
rect 64690 251308 64696 251320
rect 63552 251280 64696 251308
rect 63552 251268 63558 251280
rect 64690 251268 64696 251280
rect 64748 251308 64754 251320
rect 66806 251308 66812 251320
rect 64748 251280 66812 251308
rect 64748 251268 64754 251280
rect 66806 251268 66812 251280
rect 66864 251268 66870 251320
rect 257982 251268 257988 251320
rect 258040 251308 258046 251320
rect 259546 251308 259552 251320
rect 258040 251280 259552 251308
rect 258040 251268 258046 251280
rect 259546 251268 259552 251280
rect 259604 251268 259610 251320
rect 104802 251200 104808 251252
rect 104860 251240 104866 251252
rect 131114 251240 131120 251252
rect 104860 251212 131120 251240
rect 104860 251200 104866 251212
rect 131114 251200 131120 251212
rect 131172 251240 131178 251252
rect 132034 251240 132040 251252
rect 131172 251212 132040 251240
rect 131172 251200 131178 251212
rect 132034 251200 132040 251212
rect 132092 251200 132098 251252
rect 255314 251200 255320 251252
rect 255372 251240 255378 251252
rect 291102 251240 291108 251252
rect 255372 251212 291108 251240
rect 255372 251200 255378 251212
rect 291102 251200 291108 251212
rect 291160 251200 291166 251252
rect 98730 251132 98736 251184
rect 98788 251172 98794 251184
rect 103422 251172 103428 251184
rect 98788 251144 103428 251172
rect 98788 251132 98794 251144
rect 103422 251132 103428 251144
rect 103480 251172 103486 251184
rect 128354 251172 128360 251184
rect 103480 251144 128360 251172
rect 103480 251132 103486 251144
rect 128354 251132 128360 251144
rect 128412 251172 128418 251184
rect 129274 251172 129280 251184
rect 128412 251144 129280 251172
rect 128412 251132 128418 251144
rect 129274 251132 129280 251144
rect 129332 251132 129338 251184
rect 262490 251132 262496 251184
rect 262548 251172 262554 251184
rect 262858 251172 262864 251184
rect 262548 251144 262864 251172
rect 262548 251132 262554 251144
rect 262858 251132 262864 251144
rect 262916 251132 262922 251184
rect 269022 251132 269028 251184
rect 269080 251172 269086 251184
rect 582650 251172 582656 251184
rect 269080 251144 582656 251172
rect 269080 251132 269086 251144
rect 582650 251132 582656 251144
rect 582708 251132 582714 251184
rect 100846 251064 100852 251116
rect 100904 251104 100910 251116
rect 107562 251104 107568 251116
rect 100904 251076 107568 251104
rect 100904 251064 100910 251076
rect 107562 251064 107568 251076
rect 107620 251104 107626 251116
rect 111058 251104 111064 251116
rect 107620 251076 111064 251104
rect 107620 251064 107626 251076
rect 111058 251064 111064 251076
rect 111116 251064 111122 251116
rect 58986 250520 58992 250572
rect 59044 250560 59050 250572
rect 66806 250560 66812 250572
rect 59044 250532 66812 250560
rect 59044 250520 59050 250532
rect 66806 250520 66812 250532
rect 66864 250520 66870 250572
rect 146110 250520 146116 250572
rect 146168 250560 146174 250572
rect 158714 250560 158720 250572
rect 146168 250532 158720 250560
rect 146168 250520 146174 250532
rect 158714 250520 158720 250532
rect 158772 250520 158778 250572
rect 186314 250520 186320 250572
rect 186372 250560 186378 250572
rect 191650 250560 191656 250572
rect 186372 250532 191656 250560
rect 186372 250520 186378 250532
rect 191650 250520 191656 250532
rect 191708 250520 191714 250572
rect 255406 250520 255412 250572
rect 255464 250560 255470 250572
rect 262490 250560 262496 250572
rect 255464 250532 262496 250560
rect 255464 250520 255470 250532
rect 262490 250520 262496 250532
rect 262548 250520 262554 250572
rect 115290 250452 115296 250504
rect 115348 250492 115354 250504
rect 174722 250492 174728 250504
rect 115348 250464 174728 250492
rect 115348 250452 115354 250464
rect 174722 250452 174728 250464
rect 174780 250452 174786 250504
rect 255498 250452 255504 250504
rect 255556 250492 255562 250504
rect 267918 250492 267924 250504
rect 255556 250464 267924 250492
rect 255556 250452 255562 250464
rect 267918 250452 267924 250464
rect 267976 250492 267982 250504
rect 269022 250492 269028 250504
rect 267976 250464 269028 250492
rect 267976 250452 267982 250464
rect 269022 250452 269028 250464
rect 269080 250452 269086 250504
rect 187142 249908 187148 249960
rect 187200 249948 187206 249960
rect 192662 249948 192668 249960
rect 187200 249920 192668 249948
rect 187200 249908 187206 249920
rect 192662 249908 192668 249920
rect 192720 249908 192726 249960
rect 100846 249704 100852 249756
rect 100904 249744 100910 249756
rect 109862 249744 109868 249756
rect 100904 249716 109868 249744
rect 100904 249704 100910 249716
rect 109862 249704 109868 249716
rect 109920 249704 109926 249756
rect 254210 249364 254216 249416
rect 254268 249404 254274 249416
rect 257982 249404 257988 249416
rect 254268 249376 257988 249404
rect 254268 249364 254274 249376
rect 257982 249364 257988 249376
rect 258040 249404 258046 249416
rect 259546 249404 259552 249416
rect 258040 249376 259552 249404
rect 258040 249364 258046 249376
rect 259546 249364 259552 249376
rect 259604 249364 259610 249416
rect 53650 249024 53656 249076
rect 53708 249064 53714 249076
rect 60642 249064 60648 249076
rect 53708 249036 60648 249064
rect 53708 249024 53714 249036
rect 60642 249024 60648 249036
rect 60700 249064 60706 249076
rect 66438 249064 66444 249076
rect 60700 249036 66444 249064
rect 60700 249024 60706 249036
rect 66438 249024 66444 249036
rect 66496 249024 66502 249076
rect 109862 249024 109868 249076
rect 109920 249064 109926 249076
rect 130562 249064 130568 249076
rect 109920 249036 130568 249064
rect 109920 249024 109926 249036
rect 130562 249024 130568 249036
rect 130620 249064 130626 249076
rect 155494 249064 155500 249076
rect 130620 249036 155500 249064
rect 130620 249024 130626 249036
rect 155494 249024 155500 249036
rect 155552 249024 155558 249076
rect 166350 249024 166356 249076
rect 166408 249064 166414 249076
rect 176102 249064 176108 249076
rect 166408 249036 176108 249064
rect 166408 249024 166414 249036
rect 176102 249024 176108 249036
rect 176160 249024 176166 249076
rect 187142 248412 187148 248464
rect 187200 248452 187206 248464
rect 191006 248452 191012 248464
rect 187200 248424 191012 248452
rect 187200 248412 187206 248424
rect 191006 248412 191012 248424
rect 191064 248412 191070 248464
rect 255406 248412 255412 248464
rect 255464 248452 255470 248464
rect 278038 248452 278044 248464
rect 255464 248424 278044 248452
rect 255464 248412 255470 248424
rect 278038 248412 278044 248424
rect 278096 248412 278102 248464
rect 112530 247732 112536 247784
rect 112588 247772 112594 247784
rect 171778 247772 171784 247784
rect 112588 247744 171784 247772
rect 112588 247732 112594 247744
rect 171778 247732 171784 247744
rect 171836 247732 171842 247784
rect 107010 247664 107016 247716
rect 107068 247704 107074 247716
rect 179506 247704 179512 247716
rect 107068 247676 179512 247704
rect 107068 247664 107074 247676
rect 179506 247664 179512 247676
rect 179564 247664 179570 247716
rect 255406 247664 255412 247716
rect 255464 247704 255470 247716
rect 265066 247704 265072 247716
rect 255464 247676 265072 247704
rect 255464 247664 255470 247676
rect 265066 247664 265072 247676
rect 265124 247664 265130 247716
rect 187602 247460 187608 247512
rect 187660 247500 187666 247512
rect 190454 247500 190460 247512
rect 187660 247472 190460 247500
rect 187660 247460 187666 247472
rect 190454 247460 190460 247472
rect 190512 247460 190518 247512
rect 62022 247052 62028 247104
rect 62080 247092 62086 247104
rect 66806 247092 66812 247104
rect 62080 247064 66812 247092
rect 62080 247052 62086 247064
rect 66806 247052 66812 247064
rect 66864 247052 66870 247104
rect 179506 247052 179512 247104
rect 179564 247092 179570 247104
rect 182910 247092 182916 247104
rect 179564 247064 182916 247092
rect 179564 247052 179570 247064
rect 182910 247052 182916 247064
rect 182968 247052 182974 247104
rect 186958 247052 186964 247104
rect 187016 247092 187022 247104
rect 191742 247092 191748 247104
rect 187016 247064 191748 247092
rect 187016 247052 187022 247064
rect 191742 247052 191748 247064
rect 191800 247052 191806 247104
rect 255498 247052 255504 247104
rect 255556 247092 255562 247104
rect 265710 247092 265716 247104
rect 255556 247064 265716 247092
rect 255556 247052 255562 247064
rect 265710 247052 265716 247064
rect 265768 247092 265774 247104
rect 269206 247092 269212 247104
rect 265768 247064 269212 247092
rect 265768 247052 265774 247064
rect 269206 247052 269212 247064
rect 269264 247052 269270 247104
rect 100662 246984 100668 247036
rect 100720 247024 100726 247036
rect 124950 247024 124956 247036
rect 100720 246996 124956 247024
rect 100720 246984 100726 246996
rect 124950 246984 124956 246996
rect 125008 246984 125014 247036
rect 190362 246372 190368 246424
rect 190420 246412 190426 246424
rect 193398 246412 193404 246424
rect 190420 246384 193404 246412
rect 190420 246372 190426 246384
rect 193398 246372 193404 246384
rect 193456 246372 193462 246424
rect 99374 246304 99380 246356
rect 99432 246344 99438 246356
rect 191190 246344 191196 246356
rect 99432 246316 191196 246344
rect 99432 246304 99438 246316
rect 191190 246304 191196 246316
rect 191248 246304 191254 246356
rect 281442 246304 281448 246356
rect 281500 246344 281506 246356
rect 298278 246344 298284 246356
rect 281500 246316 298284 246344
rect 281500 246304 281506 246316
rect 298278 246304 298284 246316
rect 298336 246304 298342 246356
rect 98638 245624 98644 245676
rect 98696 245664 98702 245676
rect 99374 245664 99380 245676
rect 98696 245636 99380 245664
rect 98696 245624 98702 245636
rect 99374 245624 99380 245636
rect 99432 245624 99438 245676
rect 125134 245624 125140 245676
rect 125192 245664 125198 245676
rect 161474 245664 161480 245676
rect 125192 245636 161480 245664
rect 125192 245624 125198 245636
rect 161474 245624 161480 245636
rect 161532 245664 161538 245676
rect 162670 245664 162676 245676
rect 161532 245636 162676 245664
rect 161532 245624 161538 245636
rect 162670 245624 162676 245636
rect 162728 245624 162734 245676
rect 255498 245624 255504 245676
rect 255556 245664 255562 245676
rect 280798 245664 280804 245676
rect 255556 245636 280804 245664
rect 255556 245624 255562 245636
rect 280798 245624 280804 245636
rect 280856 245664 280862 245676
rect 281442 245664 281448 245676
rect 280856 245636 281448 245664
rect 280856 245624 280862 245636
rect 281442 245624 281448 245636
rect 281500 245624 281506 245676
rect 101030 245556 101036 245608
rect 101088 245596 101094 245608
rect 155954 245596 155960 245608
rect 101088 245568 155960 245596
rect 101088 245556 101094 245568
rect 155954 245556 155960 245568
rect 156012 245556 156018 245608
rect 255406 245556 255412 245608
rect 255464 245596 255470 245608
rect 289814 245596 289820 245608
rect 255464 245568 289820 245596
rect 255464 245556 255470 245568
rect 289814 245556 289820 245568
rect 289872 245556 289878 245608
rect 100846 245488 100852 245540
rect 100904 245528 100910 245540
rect 108390 245528 108396 245540
rect 100904 245500 108396 245528
rect 100904 245488 100910 245500
rect 108390 245488 108396 245500
rect 108448 245488 108454 245540
rect 138842 245488 138848 245540
rect 138900 245528 138906 245540
rect 187694 245528 187700 245540
rect 138900 245500 187700 245528
rect 138900 245488 138906 245500
rect 187694 245488 187700 245500
rect 187752 245488 187758 245540
rect 155954 244876 155960 244928
rect 156012 244916 156018 244928
rect 193490 244916 193496 244928
rect 156012 244888 193496 244916
rect 156012 244876 156018 244888
rect 193490 244876 193496 244888
rect 193548 244876 193554 244928
rect 255406 244264 255412 244316
rect 255464 244304 255470 244316
rect 270402 244304 270408 244316
rect 255464 244276 270408 244304
rect 255464 244264 255470 244276
rect 270402 244264 270408 244276
rect 270460 244264 270466 244316
rect 289814 244264 289820 244316
rect 289872 244304 289878 244316
rect 293954 244304 293960 244316
rect 289872 244276 293960 244304
rect 289872 244264 289878 244276
rect 293954 244264 293960 244276
rect 294012 244264 294018 244316
rect 255866 244196 255872 244248
rect 255924 244236 255930 244248
rect 285674 244236 285680 244248
rect 255924 244208 285680 244236
rect 255924 244196 255930 244208
rect 285674 244196 285680 244208
rect 285732 244196 285738 244248
rect 111150 243516 111156 243568
rect 111208 243556 111214 243568
rect 151170 243556 151176 243568
rect 111208 243528 151176 243556
rect 111208 243516 111214 243528
rect 151170 243516 151176 243528
rect 151228 243516 151234 243568
rect 183462 243516 183468 243568
rect 183520 243556 183526 243568
rect 192478 243556 192484 243568
rect 183520 243528 192484 243556
rect 183520 243516 183526 243528
rect 192478 243516 192484 243528
rect 192536 243516 192542 243568
rect 255498 243516 255504 243568
rect 255556 243556 255562 243568
rect 277486 243556 277492 243568
rect 255556 243528 277492 243556
rect 255556 243516 255562 243528
rect 277486 243516 277492 243528
rect 277544 243516 277550 243568
rect 157334 243312 157340 243364
rect 157392 243352 157398 243364
rect 158162 243352 158168 243364
rect 157392 243324 158168 243352
rect 157392 243312 157398 243324
rect 158162 243312 158168 243324
rect 158220 243312 158226 243364
rect 100846 242972 100852 243024
rect 100904 243012 100910 243024
rect 102778 243012 102784 243024
rect 100904 242984 102784 243012
rect 100904 242972 100910 242984
rect 102778 242972 102784 242984
rect 102836 242972 102842 243024
rect 52362 242904 52368 242956
rect 52420 242944 52426 242956
rect 66714 242944 66720 242956
rect 52420 242916 66720 242944
rect 52420 242904 52426 242916
rect 66714 242904 66720 242916
rect 66772 242904 66778 242956
rect 67634 242904 67640 242956
rect 67692 242944 67698 242956
rect 68462 242944 68468 242956
rect 67692 242916 68468 242944
rect 67692 242904 67698 242916
rect 68462 242904 68468 242916
rect 68520 242904 68526 242956
rect 102870 242904 102876 242956
rect 102928 242944 102934 242956
rect 157334 242944 157340 242956
rect 102928 242916 157340 242944
rect 102928 242904 102934 242916
rect 157334 242904 157340 242916
rect 157392 242904 157398 242956
rect 182082 242904 182088 242956
rect 182140 242944 182146 242956
rect 184290 242944 184296 242956
rect 182140 242916 184296 242944
rect 182140 242904 182146 242916
rect 184290 242904 184296 242916
rect 184348 242904 184354 242956
rect 3418 242156 3424 242208
rect 3476 242196 3482 242208
rect 22738 242196 22744 242208
rect 3476 242168 22744 242196
rect 3476 242156 3482 242168
rect 22738 242156 22744 242168
rect 22796 242156 22802 242208
rect 109770 242156 109776 242208
rect 109828 242196 109834 242208
rect 178862 242196 178868 242208
rect 109828 242168 178868 242196
rect 109828 242156 109834 242168
rect 178862 242156 178868 242168
rect 178920 242156 178926 242208
rect 261018 242196 261024 242208
rect 249168 242168 261024 242196
rect 100846 242088 100852 242140
rect 100904 242128 100910 242140
rect 103606 242128 103612 242140
rect 100904 242100 103612 242128
rect 100904 242088 100910 242100
rect 103606 242088 103612 242100
rect 103664 242088 103670 242140
rect 249168 242072 249196 242168
rect 261018 242156 261024 242168
rect 261076 242156 261082 242208
rect 249150 242020 249156 242072
rect 249208 242020 249214 242072
rect 249794 242020 249800 242072
rect 249852 242060 249858 242072
rect 253014 242060 253020 242072
rect 249852 242032 253020 242060
rect 249852 242020 249858 242032
rect 253014 242020 253020 242032
rect 253072 242020 253078 242072
rect 162302 241952 162308 242004
rect 162360 241992 162366 242004
rect 162762 241992 162768 242004
rect 162360 241964 162768 241992
rect 162360 241952 162366 241964
rect 162762 241952 162768 241964
rect 162820 241952 162826 242004
rect 186314 241544 186320 241596
rect 186372 241584 186378 241596
rect 191742 241584 191748 241596
rect 186372 241556 191748 241584
rect 186372 241544 186378 241556
rect 191742 241544 191748 241556
rect 191800 241544 191806 241596
rect 191834 241544 191840 241596
rect 191892 241584 191898 241596
rect 213270 241584 213276 241596
rect 191892 241556 213276 241584
rect 191892 241544 191898 241556
rect 213270 241544 213276 241556
rect 213328 241544 213334 241596
rect 53742 241476 53748 241528
rect 53800 241516 53806 241528
rect 66806 241516 66812 241528
rect 53800 241488 66812 241516
rect 53800 241476 53806 241488
rect 66806 241476 66812 241488
rect 66864 241476 66870 241528
rect 98408 241476 98414 241528
rect 98466 241516 98472 241528
rect 103422 241516 103428 241528
rect 98466 241488 103428 241516
rect 98466 241476 98472 241488
rect 103422 241476 103428 241488
rect 103480 241516 103486 241528
rect 106274 241516 106280 241528
rect 103480 241488 106280 241516
rect 103480 241476 103486 241488
rect 106274 241476 106280 241488
rect 106332 241476 106338 241528
rect 162302 241476 162308 241528
rect 162360 241516 162366 241528
rect 197170 241516 197176 241528
rect 162360 241488 197176 241516
rect 162360 241476 162366 241488
rect 197170 241476 197176 241488
rect 197228 241476 197234 241528
rect 14458 241408 14464 241460
rect 14516 241448 14522 241460
rect 93118 241448 93124 241460
rect 14516 241420 93124 241448
rect 14516 241408 14522 241420
rect 93118 241408 93124 241420
rect 93176 241448 93182 241460
rect 93440 241448 93446 241460
rect 93176 241420 93446 241448
rect 93176 241408 93182 241420
rect 93440 241408 93446 241420
rect 93498 241408 93504 241460
rect 95648 241408 95654 241460
rect 95706 241448 95712 241460
rect 110414 241448 110420 241460
rect 95706 241420 110420 241448
rect 95706 241408 95712 241420
rect 110414 241408 110420 241420
rect 110472 241408 110478 241460
rect 174722 241408 174728 241460
rect 174780 241448 174786 241460
rect 259454 241448 259460 241460
rect 174780 241420 259460 241448
rect 174780 241408 174786 241420
rect 259454 241408 259460 241420
rect 259512 241408 259518 241460
rect 73522 241340 73528 241392
rect 73580 241380 73586 241392
rect 105630 241380 105636 241392
rect 73580 241352 105636 241380
rect 73580 241340 73586 241352
rect 105630 241340 105636 241352
rect 105688 241340 105694 241392
rect 269758 241000 269764 241052
rect 269816 241040 269822 241052
rect 273438 241040 273444 241052
rect 269816 241012 273444 241040
rect 269816 241000 269822 241012
rect 273438 241000 273444 241012
rect 273496 241000 273502 241052
rect 152826 240728 152832 240780
rect 152884 240768 152890 240780
rect 180242 240768 180248 240780
rect 152884 240740 180248 240768
rect 152884 240728 152890 240740
rect 180242 240728 180248 240740
rect 180300 240728 180306 240780
rect 192662 240728 192668 240780
rect 192720 240768 192726 240780
rect 209038 240768 209044 240780
rect 192720 240740 209044 240768
rect 192720 240728 192726 240740
rect 209038 240728 209044 240740
rect 209096 240728 209102 240780
rect 244918 240728 244924 240780
rect 244976 240768 244982 240780
rect 263778 240768 263784 240780
rect 244976 240740 263784 240768
rect 244976 240728 244982 240740
rect 263778 240728 263784 240740
rect 263836 240728 263842 240780
rect 69474 240252 69480 240304
rect 69532 240252 69538 240304
rect 69492 240088 69520 240252
rect 74534 240116 74540 240168
rect 74592 240156 74598 240168
rect 74902 240156 74908 240168
rect 74592 240128 74908 240156
rect 74592 240116 74598 240128
rect 74902 240116 74908 240128
rect 74960 240116 74966 240168
rect 82814 240116 82820 240168
rect 82872 240156 82878 240168
rect 83734 240156 83740 240168
rect 82872 240128 83740 240156
rect 82872 240116 82878 240128
rect 83734 240116 83740 240128
rect 83792 240116 83798 240168
rect 84194 240116 84200 240168
rect 84252 240156 84258 240168
rect 84838 240156 84844 240168
rect 84252 240128 84844 240156
rect 84252 240116 84258 240128
rect 84838 240116 84844 240128
rect 84896 240116 84902 240168
rect 86954 240116 86960 240168
rect 87012 240156 87018 240168
rect 87598 240156 87604 240168
rect 87012 240128 87604 240156
rect 87012 240116 87018 240128
rect 87598 240116 87604 240128
rect 87656 240116 87662 240168
rect 165706 240088 165712 240100
rect 69492 240060 165712 240088
rect 165706 240048 165712 240060
rect 165764 240088 165770 240100
rect 169018 240088 169024 240100
rect 165764 240060 169024 240088
rect 165764 240048 165770 240060
rect 169018 240048 169024 240060
rect 169076 240048 169082 240100
rect 183370 240088 183376 240100
rect 180766 240060 183376 240088
rect 69014 239980 69020 240032
rect 69072 240020 69078 240032
rect 69934 240020 69940 240032
rect 69072 239992 69940 240020
rect 69072 239980 69078 239992
rect 69934 239980 69940 239992
rect 69992 239980 69998 240032
rect 70486 239980 70492 240032
rect 70544 240020 70550 240032
rect 71314 240020 71320 240032
rect 70544 239992 71320 240020
rect 70544 239980 70550 239992
rect 71314 239980 71320 239992
rect 71372 239980 71378 240032
rect 95142 239980 95148 240032
rect 95200 240020 95206 240032
rect 98730 240020 98736 240032
rect 95200 239992 98736 240020
rect 95200 239980 95206 239992
rect 98730 239980 98736 239992
rect 98788 239980 98794 240032
rect 103422 239980 103428 240032
rect 103480 240020 103486 240032
rect 180766 240020 180794 240060
rect 183370 240048 183376 240060
rect 183428 240088 183434 240100
rect 195238 240088 195244 240100
rect 183428 240060 195244 240088
rect 183428 240048 183434 240060
rect 195238 240048 195244 240060
rect 195296 240048 195302 240100
rect 213270 240048 213276 240100
rect 213328 240088 213334 240100
rect 230750 240088 230756 240100
rect 213328 240060 230756 240088
rect 213328 240048 213334 240060
rect 230750 240048 230756 240060
rect 230808 240088 230814 240100
rect 237650 240088 237656 240100
rect 230808 240060 237656 240088
rect 230808 240048 230814 240060
rect 237650 240048 237656 240060
rect 237708 240048 237714 240100
rect 251818 240048 251824 240100
rect 251876 240088 251882 240100
rect 252278 240088 252284 240100
rect 251876 240060 252284 240088
rect 251876 240048 251882 240060
rect 252278 240048 252284 240060
rect 252336 240088 252342 240100
rect 283006 240088 283012 240100
rect 252336 240060 283012 240088
rect 252336 240048 252342 240060
rect 283006 240048 283012 240060
rect 283064 240048 283070 240100
rect 103480 239992 180794 240020
rect 103480 239980 103486 239992
rect 222194 239980 222200 240032
rect 222252 240020 222258 240032
rect 223482 240020 223488 240032
rect 222252 239992 223488 240020
rect 222252 239980 222258 239992
rect 223482 239980 223488 239992
rect 223540 239980 223546 240032
rect 80054 239776 80060 239828
rect 80112 239816 80118 239828
rect 80974 239816 80980 239828
rect 80112 239788 80980 239816
rect 80112 239776 80118 239788
rect 80974 239776 80980 239788
rect 81032 239776 81038 239828
rect 224862 239572 224868 239624
rect 224920 239612 224926 239624
rect 225966 239612 225972 239624
rect 224920 239584 225972 239612
rect 224920 239572 224926 239584
rect 225966 239572 225972 239584
rect 226024 239572 226030 239624
rect 89346 239436 89352 239488
rect 89404 239476 89410 239488
rect 91922 239476 91928 239488
rect 89404 239448 91928 239476
rect 89404 239436 89410 239448
rect 91922 239436 91928 239448
rect 91980 239436 91986 239488
rect 56410 239368 56416 239420
rect 56468 239408 56474 239420
rect 71038 239408 71044 239420
rect 56468 239380 71044 239408
rect 56468 239368 56474 239380
rect 71038 239368 71044 239380
rect 71096 239368 71102 239420
rect 169018 239368 169024 239420
rect 169076 239408 169082 239420
rect 209130 239408 209136 239420
rect 169076 239380 209136 239408
rect 169076 239368 169082 239380
rect 209130 239368 209136 239380
rect 209188 239368 209194 239420
rect 237374 239368 237380 239420
rect 237432 239408 237438 239420
rect 256878 239408 256884 239420
rect 237432 239380 256884 239408
rect 237432 239368 237438 239380
rect 256878 239368 256884 239380
rect 256936 239368 256942 239420
rect 258810 239368 258816 239420
rect 258868 239408 258874 239420
rect 270770 239408 270776 239420
rect 258868 239380 270776 239408
rect 258868 239368 258874 239380
rect 270770 239368 270776 239380
rect 270828 239368 270834 239420
rect 247034 238756 247040 238808
rect 247092 238796 247098 238808
rect 252462 238796 252468 238808
rect 247092 238768 252468 238796
rect 247092 238756 247098 238768
rect 252462 238756 252468 238768
rect 252520 238756 252526 238808
rect 67818 238688 67824 238740
rect 67876 238728 67882 238740
rect 102870 238728 102876 238740
rect 67876 238700 102876 238728
rect 67876 238688 67882 238700
rect 102870 238688 102876 238700
rect 102928 238688 102934 238740
rect 180058 238688 180064 238740
rect 180116 238728 180122 238740
rect 213914 238728 213920 238740
rect 180116 238700 213920 238728
rect 180116 238688 180122 238700
rect 213914 238688 213920 238700
rect 213972 238688 213978 238740
rect 221090 238688 221096 238740
rect 221148 238728 221154 238740
rect 273898 238728 273904 238740
rect 221148 238700 273904 238728
rect 221148 238688 221154 238700
rect 273898 238688 273904 238700
rect 273956 238688 273962 238740
rect 193582 238620 193588 238672
rect 193640 238660 193646 238672
rect 215294 238660 215300 238672
rect 193640 238632 215300 238660
rect 193640 238620 193646 238632
rect 215294 238620 215300 238632
rect 215352 238620 215358 238672
rect 242710 238620 242716 238672
rect 242768 238660 242774 238672
rect 274634 238660 274640 238672
rect 242768 238632 274640 238660
rect 242768 238620 242774 238632
rect 274634 238620 274640 238632
rect 274692 238620 274698 238672
rect 215294 238348 215300 238400
rect 215352 238388 215358 238400
rect 216306 238388 216312 238400
rect 215352 238360 216312 238388
rect 215352 238348 215358 238360
rect 216306 238348 216312 238360
rect 216364 238348 216370 238400
rect 106274 238076 106280 238128
rect 106332 238116 106338 238128
rect 173250 238116 173256 238128
rect 106332 238088 173256 238116
rect 106332 238076 106338 238088
rect 173250 238076 173256 238088
rect 173308 238076 173314 238128
rect 96890 238008 96896 238060
rect 96948 238048 96954 238060
rect 108390 238048 108396 238060
rect 96948 238020 108396 238048
rect 96948 238008 96954 238020
rect 108390 238008 108396 238020
rect 108448 238008 108454 238060
rect 110414 238008 110420 238060
rect 110472 238048 110478 238060
rect 180794 238048 180800 238060
rect 110472 238020 180800 238048
rect 110472 238008 110478 238020
rect 180794 238008 180800 238020
rect 180852 238008 180858 238060
rect 213914 237396 213920 237448
rect 213972 237436 213978 237448
rect 214650 237436 214656 237448
rect 213972 237408 214656 237436
rect 213972 237396 213978 237408
rect 214650 237396 214656 237408
rect 214708 237396 214714 237448
rect 242250 237396 242256 237448
rect 242308 237436 242314 237448
rect 242710 237436 242716 237448
rect 242308 237408 242716 237436
rect 242308 237396 242314 237408
rect 242710 237396 242716 237408
rect 242768 237396 242774 237448
rect 92566 237328 92572 237380
rect 92624 237368 92630 237380
rect 125042 237368 125048 237380
rect 92624 237340 125048 237368
rect 92624 237328 92630 237340
rect 125042 237328 125048 237340
rect 125100 237328 125106 237380
rect 169754 237328 169760 237380
rect 169812 237368 169818 237380
rect 189718 237368 189724 237380
rect 169812 237340 189724 237368
rect 169812 237328 169818 237340
rect 189718 237328 189724 237340
rect 189776 237328 189782 237380
rect 193674 237328 193680 237380
rect 193732 237368 193738 237380
rect 237926 237368 237932 237380
rect 193732 237340 237932 237368
rect 193732 237328 193738 237340
rect 237926 237328 237932 237340
rect 237984 237328 237990 237380
rect 177390 237260 177396 237312
rect 177448 237300 177454 237312
rect 201494 237300 201500 237312
rect 177448 237272 201500 237300
rect 177448 237260 177454 237272
rect 201494 237260 201500 237272
rect 201552 237300 201558 237312
rect 201954 237300 201960 237312
rect 201552 237272 201960 237300
rect 201552 237260 201558 237272
rect 201954 237260 201960 237272
rect 202012 237260 202018 237312
rect 74442 236648 74448 236700
rect 74500 236688 74506 236700
rect 77294 236688 77300 236700
rect 74500 236660 77300 236688
rect 74500 236648 74506 236660
rect 77294 236648 77300 236660
rect 77352 236648 77358 236700
rect 207658 236648 207664 236700
rect 207716 236688 207722 236700
rect 221090 236688 221096 236700
rect 207716 236660 221096 236688
rect 207716 236648 207722 236660
rect 221090 236648 221096 236660
rect 221148 236648 221154 236700
rect 242158 236648 242164 236700
rect 242216 236688 242222 236700
rect 266446 236688 266452 236700
rect 242216 236660 266452 236688
rect 242216 236648 242222 236660
rect 266446 236648 266452 236660
rect 266504 236648 266510 236700
rect 89622 236444 89628 236496
rect 89680 236484 89686 236496
rect 91094 236484 91100 236496
rect 89680 236456 91100 236484
rect 89680 236444 89686 236456
rect 91094 236444 91100 236456
rect 91152 236444 91158 236496
rect 91094 236308 91100 236360
rect 91152 236348 91158 236360
rect 94774 236348 94780 236360
rect 91152 236320 94780 236348
rect 91152 236308 91158 236320
rect 94774 236308 94780 236320
rect 94832 236308 94838 236360
rect 77662 236172 77668 236224
rect 77720 236212 77726 236224
rect 83550 236212 83556 236224
rect 77720 236184 83556 236212
rect 77720 236172 77726 236184
rect 83550 236172 83556 236184
rect 83608 236172 83614 236224
rect 91186 235968 91192 236020
rect 91244 235968 91250 236020
rect 94682 235968 94688 236020
rect 94740 236008 94746 236020
rect 95234 236008 95240 236020
rect 94740 235980 95240 236008
rect 94740 235968 94746 235980
rect 95234 235968 95240 235980
rect 95292 235968 95298 236020
rect 237466 235968 237472 236020
rect 237524 236008 237530 236020
rect 237926 236008 237932 236020
rect 237524 235980 237932 236008
rect 237524 235968 237530 235980
rect 237926 235968 237932 235980
rect 237984 235968 237990 236020
rect 91204 235940 91232 235968
rect 124306 235940 124312 235952
rect 91204 235912 124312 235940
rect 124306 235900 124312 235912
rect 124364 235900 124370 235952
rect 192570 235900 192576 235952
rect 192628 235940 192634 235952
rect 205726 235940 205732 235952
rect 192628 235912 205732 235940
rect 192628 235900 192634 235912
rect 205726 235900 205732 235912
rect 205784 235900 205790 235952
rect 205726 235424 205732 235476
rect 205784 235464 205790 235476
rect 206738 235464 206744 235476
rect 205784 235436 206744 235464
rect 205784 235424 205790 235436
rect 206738 235424 206744 235436
rect 206796 235424 206802 235476
rect 193122 235288 193128 235340
rect 193180 235328 193186 235340
rect 220814 235328 220820 235340
rect 193180 235300 220820 235328
rect 193180 235288 193186 235300
rect 220814 235288 220820 235300
rect 220872 235288 220878 235340
rect 222838 235288 222844 235340
rect 222896 235328 222902 235340
rect 252738 235328 252744 235340
rect 222896 235300 252744 235328
rect 222896 235288 222902 235300
rect 252738 235288 252744 235300
rect 252796 235288 252802 235340
rect 213178 235220 213184 235272
rect 213236 235260 213242 235272
rect 255498 235260 255504 235272
rect 213236 235232 255504 235260
rect 213236 235220 213242 235232
rect 255498 235220 255504 235232
rect 255556 235260 255562 235272
rect 582650 235260 582656 235272
rect 255556 235232 582656 235260
rect 255556 235220 255562 235232
rect 582650 235220 582656 235232
rect 582708 235220 582714 235272
rect 82078 234540 82084 234592
rect 82136 234580 82142 234592
rect 108482 234580 108488 234592
rect 82136 234552 108488 234580
rect 82136 234540 82142 234552
rect 108482 234540 108488 234552
rect 108540 234540 108546 234592
rect 185578 234540 185584 234592
rect 185636 234580 185642 234592
rect 256970 234580 256976 234592
rect 185636 234552 256976 234580
rect 185636 234540 185642 234552
rect 256970 234540 256976 234552
rect 257028 234540 257034 234592
rect 67726 233996 67732 234048
rect 67784 234036 67790 234048
rect 71774 234036 71780 234048
rect 67784 234008 71780 234036
rect 67784 233996 67790 234008
rect 71774 233996 71780 234008
rect 71832 233996 71838 234048
rect 97902 233860 97908 233912
rect 97960 233900 97966 233912
rect 99466 233900 99472 233912
rect 97960 233872 99472 233900
rect 97960 233860 97966 233872
rect 99466 233860 99472 233872
rect 99524 233860 99530 233912
rect 177390 233860 177396 233912
rect 177448 233900 177454 233912
rect 259730 233900 259736 233912
rect 177448 233872 259736 233900
rect 177448 233860 177454 233872
rect 259730 233860 259736 233872
rect 259788 233860 259794 233912
rect 290458 233656 290464 233708
rect 290516 233696 290522 233708
rect 291102 233696 291108 233708
rect 290516 233668 291108 233696
rect 290516 233656 290522 233668
rect 291102 233656 291108 233668
rect 291160 233656 291166 233708
rect 291102 233248 291108 233300
rect 291160 233288 291166 233300
rect 580258 233288 580264 233300
rect 291160 233260 580264 233288
rect 291160 233248 291166 233260
rect 580258 233248 580264 233260
rect 580316 233248 580322 233300
rect 80330 233180 80336 233232
rect 80388 233220 80394 233232
rect 161474 233220 161480 233232
rect 80388 233192 161480 233220
rect 80388 233180 80394 233192
rect 161474 233180 161480 233192
rect 161532 233220 161538 233232
rect 162302 233220 162308 233232
rect 161532 233192 162308 233220
rect 161532 233180 161538 233192
rect 162302 233180 162308 233192
rect 162360 233180 162366 233232
rect 174630 233180 174636 233232
rect 174688 233220 174694 233232
rect 175182 233220 175188 233232
rect 174688 233192 175188 233220
rect 174688 233180 174694 233192
rect 175182 233180 175188 233192
rect 175240 233220 175246 233232
rect 259638 233220 259644 233232
rect 175240 233192 259644 233220
rect 175240 233180 175246 233192
rect 259638 233180 259644 233192
rect 259696 233180 259702 233232
rect 278038 233180 278044 233232
rect 278096 233220 278102 233232
rect 281810 233220 281816 233232
rect 278096 233192 281816 233220
rect 278096 233180 278102 233192
rect 281810 233180 281816 233192
rect 281868 233180 281874 233232
rect 117958 233112 117964 233164
rect 118016 233152 118022 233164
rect 121638 233152 121644 233164
rect 118016 233124 121644 233152
rect 118016 233112 118022 233124
rect 121638 233112 121644 233124
rect 121696 233112 121702 233164
rect 266998 232568 267004 232620
rect 267056 232608 267062 232620
rect 276290 232608 276296 232620
rect 267056 232580 276296 232608
rect 267056 232568 267062 232580
rect 276290 232568 276296 232580
rect 276348 232568 276354 232620
rect 88334 232500 88340 232552
rect 88392 232540 88398 232552
rect 117958 232540 117964 232552
rect 88392 232512 117964 232540
rect 88392 232500 88398 232512
rect 117958 232500 117964 232512
rect 118016 232500 118022 232552
rect 133230 232500 133236 232552
rect 133288 232540 133294 232552
rect 210418 232540 210424 232552
rect 133288 232512 210424 232540
rect 133288 232500 133294 232512
rect 210418 232500 210424 232512
rect 210476 232500 210482 232552
rect 239398 232500 239404 232552
rect 239456 232540 239462 232552
rect 274910 232540 274916 232552
rect 239456 232512 274916 232540
rect 239456 232500 239462 232512
rect 274910 232500 274916 232512
rect 274968 232500 274974 232552
rect 281810 231820 281816 231872
rect 281868 231860 281874 231872
rect 580166 231860 580172 231872
rect 281868 231832 580172 231860
rect 281868 231820 281874 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 79962 231140 79968 231192
rect 80020 231180 80026 231192
rect 87598 231180 87604 231192
rect 80020 231152 87604 231180
rect 80020 231140 80026 231152
rect 87598 231140 87604 231152
rect 87656 231140 87662 231192
rect 89714 231140 89720 231192
rect 89772 231180 89778 231192
rect 124122 231180 124128 231192
rect 89772 231152 124128 231180
rect 89772 231140 89778 231152
rect 124122 231140 124128 231152
rect 124180 231180 124186 231192
rect 130654 231180 130660 231192
rect 124180 231152 130660 231180
rect 124180 231140 124186 231152
rect 130654 231140 130660 231152
rect 130712 231140 130718 231192
rect 153930 231140 153936 231192
rect 153988 231180 153994 231192
rect 215938 231180 215944 231192
rect 153988 231152 215944 231180
rect 153988 231140 153994 231152
rect 215938 231140 215944 231152
rect 215996 231140 216002 231192
rect 60366 231072 60372 231124
rect 60424 231112 60430 231124
rect 79318 231112 79324 231124
rect 60424 231084 79324 231112
rect 60424 231072 60430 231084
rect 79318 231072 79324 231084
rect 79376 231072 79382 231124
rect 84194 231072 84200 231124
rect 84252 231112 84258 231124
rect 114738 231112 114744 231124
rect 84252 231084 114744 231112
rect 84252 231072 84258 231084
rect 114738 231072 114744 231084
rect 114796 231112 114802 231124
rect 182542 231112 182548 231124
rect 114796 231084 182548 231112
rect 114796 231072 114802 231084
rect 182542 231072 182548 231084
rect 182600 231072 182606 231124
rect 235258 231072 235264 231124
rect 235316 231112 235322 231124
rect 255682 231112 255688 231124
rect 235316 231084 255688 231112
rect 235316 231072 235322 231084
rect 255682 231072 255688 231084
rect 255740 231072 255746 231124
rect 257338 231072 257344 231124
rect 257396 231112 257402 231124
rect 278958 231112 278964 231124
rect 257396 231084 278964 231112
rect 257396 231072 257402 231084
rect 278958 231072 278964 231084
rect 279016 231072 279022 231124
rect 179230 230392 179236 230444
rect 179288 230432 179294 230444
rect 215386 230432 215392 230444
rect 179288 230404 215392 230432
rect 179288 230392 179294 230404
rect 215386 230392 215392 230404
rect 215444 230392 215450 230444
rect 63218 229712 63224 229764
rect 63276 229752 63282 229764
rect 75914 229752 75920 229764
rect 63276 229724 75920 229752
rect 63276 229712 63282 229724
rect 75914 229712 75920 229724
rect 75972 229712 75978 229764
rect 184750 229712 184756 229764
rect 184808 229752 184814 229764
rect 203518 229752 203524 229764
rect 184808 229724 203524 229752
rect 184808 229712 184814 229724
rect 203518 229712 203524 229724
rect 203576 229712 203582 229764
rect 3418 229168 3424 229220
rect 3476 229208 3482 229220
rect 96982 229208 96988 229220
rect 3476 229180 96988 229208
rect 3476 229168 3482 229180
rect 96982 229168 96988 229180
rect 97040 229168 97046 229220
rect 75914 229100 75920 229152
rect 75972 229140 75978 229152
rect 175918 229140 175924 229152
rect 75972 229112 175924 229140
rect 75972 229100 75978 229112
rect 175918 229100 175924 229112
rect 175976 229100 175982 229152
rect 107562 229032 107568 229084
rect 107620 229072 107626 229084
rect 280338 229072 280344 229084
rect 107620 229044 280344 229072
rect 107620 229032 107626 229044
rect 280338 229032 280344 229044
rect 280396 229032 280402 229084
rect 191190 228964 191196 229016
rect 191248 229004 191254 229016
rect 253198 229004 253204 229016
rect 191248 228976 253204 229004
rect 191248 228964 191254 228976
rect 253198 228964 253204 228976
rect 253256 228964 253262 229016
rect 106918 228692 106924 228744
rect 106976 228732 106982 228744
rect 107562 228732 107568 228744
rect 106976 228704 107568 228732
rect 106976 228692 106982 228704
rect 107562 228692 107568 228704
rect 107620 228692 107626 228744
rect 80054 228352 80060 228404
rect 80112 228392 80118 228404
rect 106366 228392 106372 228404
rect 80112 228364 106372 228392
rect 80112 228352 80118 228364
rect 106366 228352 106372 228364
rect 106424 228392 106430 228404
rect 111150 228392 111156 228404
rect 106424 228364 111156 228392
rect 106424 228352 106430 228364
rect 111150 228352 111156 228364
rect 111208 228352 111214 228404
rect 96522 227740 96528 227792
rect 96580 227780 96586 227792
rect 100846 227780 100852 227792
rect 96580 227752 100852 227780
rect 96580 227740 96586 227752
rect 100846 227740 100852 227752
rect 100904 227740 100910 227792
rect 252738 227740 252744 227792
rect 252796 227780 252802 227792
rect 253198 227780 253204 227792
rect 252796 227752 253204 227780
rect 252796 227740 252802 227752
rect 253198 227740 253204 227752
rect 253256 227740 253262 227792
rect 149882 227672 149888 227724
rect 149940 227712 149946 227724
rect 262398 227712 262404 227724
rect 149940 227684 262404 227712
rect 149940 227672 149946 227684
rect 262398 227672 262404 227684
rect 262456 227672 262462 227724
rect 158162 227604 158168 227656
rect 158220 227644 158226 227656
rect 204346 227644 204352 227656
rect 158220 227616 204352 227644
rect 158220 227604 158226 227616
rect 204346 227604 204352 227616
rect 204404 227604 204410 227656
rect 78582 226992 78588 227044
rect 78640 227032 78646 227044
rect 111150 227032 111156 227044
rect 78640 227004 111156 227032
rect 78640 226992 78646 227004
rect 111150 226992 111156 227004
rect 111208 227032 111214 227044
rect 118050 227032 118056 227044
rect 111208 227004 118056 227032
rect 111208 226992 111214 227004
rect 118050 226992 118056 227004
rect 118108 226992 118114 227044
rect 158162 226312 158168 226364
rect 158220 226352 158226 226364
rect 158622 226352 158628 226364
rect 158220 226324 158628 226352
rect 158220 226312 158226 226324
rect 158622 226312 158628 226324
rect 158680 226312 158686 226364
rect 108298 225632 108304 225684
rect 108356 225672 108362 225684
rect 122098 225672 122104 225684
rect 108356 225644 122104 225672
rect 108356 225632 108362 225644
rect 122098 225632 122104 225644
rect 122156 225632 122162 225684
rect 184382 225632 184388 225684
rect 184440 225672 184446 225684
rect 244274 225672 244280 225684
rect 184440 225644 244280 225672
rect 184440 225632 184446 225644
rect 244274 225632 244280 225644
rect 244332 225632 244338 225684
rect 109678 225564 109684 225616
rect 109736 225604 109742 225616
rect 245654 225604 245660 225616
rect 109736 225576 245660 225604
rect 109736 225564 109742 225576
rect 245654 225564 245660 225576
rect 245712 225604 245718 225616
rect 265066 225604 265072 225616
rect 245712 225576 265072 225604
rect 245712 225564 245718 225576
rect 265066 225564 265072 225576
rect 265124 225564 265130 225616
rect 244274 224884 244280 224936
rect 244332 224924 244338 224936
rect 245010 224924 245016 224936
rect 244332 224896 245016 224924
rect 244332 224884 244338 224896
rect 245010 224884 245016 224896
rect 245068 224924 245074 224936
rect 272058 224924 272064 224936
rect 245068 224896 272064 224924
rect 245068 224884 245074 224896
rect 272058 224884 272064 224896
rect 272116 224884 272122 224936
rect 91370 224272 91376 224324
rect 91428 224312 91434 224324
rect 182910 224312 182916 224324
rect 91428 224284 182916 224312
rect 91428 224272 91434 224284
rect 182910 224272 182916 224284
rect 182968 224272 182974 224324
rect 178862 224204 178868 224256
rect 178920 224244 178926 224256
rect 219434 224244 219440 224256
rect 178920 224216 219440 224244
rect 178920 224204 178926 224216
rect 219434 224204 219440 224216
rect 219492 224244 219498 224256
rect 281718 224244 281724 224256
rect 219492 224216 281724 224244
rect 219492 224204 219498 224216
rect 281718 224204 281724 224216
rect 281776 224204 281782 224256
rect 196710 223524 196716 223576
rect 196768 223564 196774 223576
rect 197262 223564 197268 223576
rect 196768 223536 197268 223564
rect 196768 223524 196774 223536
rect 197262 223524 197268 223536
rect 197320 223564 197326 223576
rect 269298 223564 269304 223576
rect 197320 223536 269304 223564
rect 197320 223524 197326 223536
rect 269298 223524 269304 223536
rect 269356 223524 269362 223576
rect 102778 222844 102784 222896
rect 102836 222884 102842 222896
rect 204898 222884 204904 222896
rect 102836 222856 204904 222884
rect 102836 222844 102842 222856
rect 204898 222844 204904 222856
rect 204956 222844 204962 222896
rect 214558 222844 214564 222896
rect 214616 222884 214622 222896
rect 255590 222884 255596 222896
rect 214616 222856 255596 222884
rect 214616 222844 214622 222856
rect 255590 222844 255596 222856
rect 255648 222844 255654 222896
rect 87046 222096 87052 222148
rect 87104 222136 87110 222148
rect 116026 222136 116032 222148
rect 87104 222108 116032 222136
rect 87104 222096 87110 222108
rect 116026 222096 116032 222108
rect 116084 222136 116090 222148
rect 116578 222136 116584 222148
rect 116084 222108 116584 222136
rect 116084 222096 116090 222108
rect 116578 222096 116584 222108
rect 116636 222096 116642 222148
rect 112622 221416 112628 221468
rect 112680 221456 112686 221468
rect 270586 221456 270592 221468
rect 112680 221428 270592 221456
rect 112680 221416 112686 221428
rect 270586 221416 270592 221428
rect 270644 221416 270650 221468
rect 97994 220736 98000 220788
rect 98052 220776 98058 220788
rect 98914 220776 98920 220788
rect 98052 220748 98920 220776
rect 98052 220736 98058 220748
rect 98914 220736 98920 220748
rect 98972 220736 98978 220788
rect 215938 220736 215944 220788
rect 215996 220776 216002 220788
rect 292666 220776 292672 220788
rect 215996 220748 292672 220776
rect 215996 220736 216002 220748
rect 292666 220736 292672 220748
rect 292724 220736 292730 220788
rect 59170 220124 59176 220176
rect 59228 220164 59234 220176
rect 159542 220164 159548 220176
rect 59228 220136 159548 220164
rect 59228 220124 59234 220136
rect 159542 220124 159548 220136
rect 159600 220124 159606 220176
rect 266354 220096 266360 220108
rect 103486 220068 266360 220096
rect 98914 219988 98920 220040
rect 98972 220028 98978 220040
rect 103486 220028 103514 220068
rect 266354 220056 266360 220068
rect 266412 220056 266418 220108
rect 98972 220000 103514 220028
rect 98972 219988 98978 220000
rect 159542 219376 159548 219428
rect 159600 219416 159606 219428
rect 258810 219416 258816 219428
rect 159600 219388 258816 219416
rect 159600 219376 159606 219388
rect 258810 219376 258816 219388
rect 258868 219376 258874 219428
rect 213270 219308 213276 219360
rect 213328 219348 213334 219360
rect 285950 219348 285956 219360
rect 213328 219320 285956 219348
rect 213328 219308 213334 219320
rect 285950 219308 285956 219320
rect 286008 219308 286014 219360
rect 285674 218764 285680 218816
rect 285732 218804 285738 218816
rect 285950 218804 285956 218816
rect 285732 218776 285956 218804
rect 285732 218764 285738 218776
rect 285950 218764 285956 218776
rect 286008 218764 286014 218816
rect 82814 218696 82820 218748
rect 82872 218736 82878 218748
rect 180058 218736 180064 218748
rect 82872 218708 180064 218736
rect 82872 218696 82878 218708
rect 180058 218696 180064 218708
rect 180116 218736 180122 218748
rect 213178 218736 213184 218748
rect 180116 218708 213184 218736
rect 180116 218696 180122 218708
rect 213178 218696 213184 218708
rect 213236 218696 213242 218748
rect 182910 217948 182916 218000
rect 182968 217988 182974 218000
rect 246298 217988 246304 218000
rect 182968 217960 246304 217988
rect 182968 217948 182974 217960
rect 246298 217948 246304 217960
rect 246356 217948 246362 218000
rect 155402 217268 155408 217320
rect 155460 217308 155466 217320
rect 247034 217308 247040 217320
rect 155460 217280 247040 217308
rect 155460 217268 155466 217280
rect 247034 217268 247040 217280
rect 247092 217268 247098 217320
rect 285122 217268 285128 217320
rect 285180 217308 285186 217320
rect 295518 217308 295524 217320
rect 285180 217280 295524 217308
rect 285180 217268 285186 217280
rect 295518 217268 295524 217280
rect 295576 217268 295582 217320
rect 74534 217132 74540 217184
rect 74592 217172 74598 217184
rect 75638 217172 75644 217184
rect 74592 217144 75644 217172
rect 74592 217132 74598 217144
rect 75638 217132 75644 217144
rect 75696 217132 75702 217184
rect 75638 216656 75644 216708
rect 75696 216696 75702 216708
rect 172330 216696 172336 216708
rect 75696 216668 172336 216696
rect 75696 216656 75702 216668
rect 172330 216656 172336 216668
rect 172388 216656 172394 216708
rect 137554 215976 137560 216028
rect 137612 216016 137618 216028
rect 220078 216016 220084 216028
rect 137612 215988 220084 216016
rect 137612 215976 137618 215988
rect 220078 215976 220084 215988
rect 220136 215976 220142 216028
rect 256050 215976 256056 216028
rect 256108 216016 256114 216028
rect 268010 216016 268016 216028
rect 256108 215988 268016 216016
rect 256108 215976 256114 215988
rect 268010 215976 268016 215988
rect 268068 215976 268074 216028
rect 86954 215908 86960 215960
rect 87012 215948 87018 215960
rect 88242 215948 88248 215960
rect 87012 215920 88248 215948
rect 87012 215908 87018 215920
rect 88242 215908 88248 215920
rect 88300 215948 88306 215960
rect 262214 215948 262220 215960
rect 88300 215920 262220 215948
rect 88300 215908 88306 215920
rect 262214 215908 262220 215920
rect 262272 215908 262278 215960
rect 156690 215228 156696 215280
rect 156748 215268 156754 215280
rect 281810 215268 281816 215280
rect 156748 215240 281816 215268
rect 156748 215228 156754 215240
rect 281810 215228 281816 215240
rect 281868 215228 281874 215280
rect 3510 214888 3516 214940
rect 3568 214928 3574 214940
rect 7558 214928 7564 214940
rect 3568 214900 7564 214928
rect 3568 214888 3574 214900
rect 7558 214888 7564 214900
rect 7616 214888 7622 214940
rect 169754 214548 169760 214600
rect 169812 214588 169818 214600
rect 257338 214588 257344 214600
rect 169812 214560 257344 214588
rect 169812 214548 169818 214560
rect 257338 214548 257344 214560
rect 257396 214548 257402 214600
rect 93118 213868 93124 213920
rect 93176 213908 93182 213920
rect 95694 213908 95700 213920
rect 93176 213880 95700 213908
rect 93176 213868 93182 213880
rect 95694 213868 95700 213880
rect 95752 213868 95758 213920
rect 149790 213868 149796 213920
rect 149848 213908 149854 213920
rect 169754 213908 169760 213920
rect 149848 213880 169760 213908
rect 149848 213868 149854 213880
rect 169754 213868 169760 213880
rect 169812 213868 169818 213920
rect 182818 213868 182824 213920
rect 182876 213908 182882 213920
rect 183462 213908 183468 213920
rect 182876 213880 183468 213908
rect 182876 213868 182882 213880
rect 183462 213868 183468 213880
rect 183520 213908 183526 213920
rect 239398 213908 239404 213920
rect 183520 213880 239404 213908
rect 183520 213868 183526 213880
rect 239398 213868 239404 213880
rect 239456 213868 239462 213920
rect 95234 212508 95240 212560
rect 95292 212548 95298 212560
rect 95694 212548 95700 212560
rect 95292 212520 95700 212548
rect 95292 212508 95298 212520
rect 95694 212508 95700 212520
rect 95752 212548 95758 212560
rect 273346 212548 273352 212560
rect 95752 212520 273352 212548
rect 95752 212508 95758 212520
rect 273346 212508 273352 212520
rect 273404 212508 273410 212560
rect 103606 212440 103612 212492
rect 103664 212480 103670 212492
rect 264974 212480 264980 212492
rect 103664 212452 264980 212480
rect 103664 212440 103670 212452
rect 264974 212440 264980 212452
rect 265032 212440 265038 212492
rect 108390 211760 108396 211812
rect 108448 211800 108454 211812
rect 270494 211800 270500 211812
rect 108448 211772 270500 211800
rect 108448 211760 108454 211772
rect 270494 211760 270500 211772
rect 270552 211760 270558 211812
rect 98822 211148 98828 211200
rect 98880 211188 98886 211200
rect 103606 211188 103612 211200
rect 98880 211160 103612 211188
rect 98880 211148 98886 211160
rect 103606 211148 103612 211160
rect 103664 211148 103670 211200
rect 50890 211080 50896 211132
rect 50948 211120 50954 211132
rect 166994 211120 167000 211132
rect 50948 211092 167000 211120
rect 50948 211080 50954 211092
rect 166994 211080 167000 211092
rect 167052 211120 167058 211132
rect 249794 211120 249800 211132
rect 167052 211092 249800 211120
rect 167052 211080 167058 211092
rect 249794 211080 249800 211092
rect 249852 211080 249858 211132
rect 138014 211012 138020 211064
rect 138072 211052 138078 211064
rect 138750 211052 138756 211064
rect 138072 211024 138756 211052
rect 138072 211012 138078 211024
rect 138750 211012 138756 211024
rect 138808 211052 138814 211064
rect 177390 211052 177396 211064
rect 138808 211024 177396 211052
rect 138808 211012 138814 211024
rect 177390 211012 177396 211024
rect 177448 211012 177454 211064
rect 59170 209040 59176 209092
rect 59228 209080 59234 209092
rect 69014 209080 69020 209092
rect 59228 209052 69020 209080
rect 59228 209040 59234 209052
rect 69014 209040 69020 209052
rect 69072 209040 69078 209092
rect 176562 208292 176568 208344
rect 176620 208332 176626 208344
rect 290458 208332 290464 208344
rect 176620 208304 290464 208332
rect 176620 208292 176626 208304
rect 290458 208292 290464 208304
rect 290516 208292 290522 208344
rect 176010 207816 176016 207868
rect 176068 207856 176074 207868
rect 176562 207856 176568 207868
rect 176068 207828 176568 207856
rect 176068 207816 176074 207828
rect 176562 207816 176568 207828
rect 176620 207816 176626 207868
rect 97258 207000 97264 207052
rect 97316 207040 97322 207052
rect 102226 207040 102232 207052
rect 97316 207012 102232 207040
rect 97316 207000 97322 207012
rect 102226 207000 102232 207012
rect 102284 207040 102290 207052
rect 263686 207040 263692 207052
rect 102284 207012 263692 207040
rect 102284 207000 102290 207012
rect 263686 207000 263692 207012
rect 263744 207000 263750 207052
rect 265066 206932 265072 206984
rect 265124 206972 265130 206984
rect 265710 206972 265716 206984
rect 265124 206944 265716 206972
rect 265124 206932 265130 206944
rect 265710 206932 265716 206944
rect 265768 206972 265774 206984
rect 579798 206972 579804 206984
rect 265768 206944 579804 206972
rect 265768 206932 265774 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 93854 206320 93860 206372
rect 93912 206360 93918 206372
rect 104986 206360 104992 206372
rect 93912 206332 104992 206360
rect 93912 206320 93918 206332
rect 104986 206320 104992 206332
rect 105044 206360 105050 206372
rect 105722 206360 105728 206372
rect 105044 206332 105728 206360
rect 105044 206320 105050 206332
rect 105722 206320 105728 206332
rect 105780 206320 105786 206372
rect 95878 206252 95884 206304
rect 95936 206292 95942 206304
rect 256694 206292 256700 206304
rect 95936 206264 256700 206292
rect 95936 206252 95942 206264
rect 256694 206252 256700 206264
rect 256752 206252 256758 206304
rect 95326 205980 95332 206032
rect 95384 206020 95390 206032
rect 95878 206020 95884 206032
rect 95384 205992 95884 206020
rect 95384 205980 95390 205992
rect 95878 205980 95884 205992
rect 95936 205980 95942 206032
rect 105722 205640 105728 205692
rect 105780 205680 105786 205692
rect 258074 205680 258080 205692
rect 105780 205652 258080 205680
rect 105780 205640 105786 205652
rect 258074 205640 258080 205652
rect 258132 205680 258138 205692
rect 258350 205680 258356 205692
rect 258132 205652 258356 205680
rect 258132 205640 258138 205652
rect 258350 205640 258356 205652
rect 258408 205640 258414 205692
rect 96614 204892 96620 204944
rect 96672 204932 96678 204944
rect 111886 204932 111892 204944
rect 96672 204904 111892 204932
rect 96672 204892 96678 204904
rect 111886 204892 111892 204904
rect 111944 204892 111950 204944
rect 274634 204688 274640 204740
rect 274692 204728 274698 204740
rect 274818 204728 274824 204740
rect 274692 204700 274824 204728
rect 274692 204688 274698 204700
rect 274818 204688 274824 204700
rect 274876 204688 274882 204740
rect 111886 204280 111892 204332
rect 111944 204320 111950 204332
rect 274634 204320 274640 204332
rect 111944 204292 274640 204320
rect 111944 204280 111950 204292
rect 274634 204280 274640 204292
rect 274692 204280 274698 204332
rect 191098 204212 191104 204264
rect 191156 204252 191162 204264
rect 193306 204252 193312 204264
rect 191156 204224 193312 204252
rect 191156 204212 191162 204224
rect 193306 204212 193312 204224
rect 193364 204212 193370 204264
rect 188982 203532 188988 203584
rect 189040 203572 189046 203584
rect 195974 203572 195980 203584
rect 189040 203544 195980 203572
rect 189040 203532 189046 203544
rect 195974 203532 195980 203544
rect 196032 203532 196038 203584
rect 97994 202784 98000 202836
rect 98052 202824 98058 202836
rect 98914 202824 98920 202836
rect 98052 202796 98920 202824
rect 98052 202784 98058 202796
rect 98914 202784 98920 202796
rect 98972 202784 98978 202836
rect 180150 202172 180156 202224
rect 180208 202212 180214 202224
rect 196618 202212 196624 202224
rect 180208 202184 196624 202212
rect 180208 202172 180214 202184
rect 196618 202172 196624 202184
rect 196676 202172 196682 202224
rect 3510 202104 3516 202156
rect 3568 202144 3574 202156
rect 97994 202144 98000 202156
rect 3568 202116 98000 202144
rect 3568 202104 3574 202116
rect 97994 202104 98000 202116
rect 98052 202104 98058 202156
rect 195882 202104 195888 202156
rect 195940 202144 195946 202156
rect 253934 202144 253940 202156
rect 195940 202116 253940 202144
rect 195940 202104 195946 202116
rect 253934 202104 253940 202116
rect 253992 202104 253998 202156
rect 260190 200812 260196 200864
rect 260248 200852 260254 200864
rect 271966 200852 271972 200864
rect 260248 200824 271972 200852
rect 260248 200812 260254 200824
rect 271966 200812 271972 200824
rect 272024 200812 272030 200864
rect 44082 200744 44088 200796
rect 44140 200784 44146 200796
rect 134702 200784 134708 200796
rect 44140 200756 134708 200784
rect 44140 200744 44146 200756
rect 134702 200744 134708 200756
rect 134760 200744 134766 200796
rect 149790 200744 149796 200796
rect 149848 200784 149854 200796
rect 188338 200784 188344 200796
rect 149848 200756 188344 200784
rect 149848 200744 149854 200756
rect 188338 200744 188344 200756
rect 188396 200744 188402 200796
rect 200022 200744 200028 200796
rect 200080 200784 200086 200796
rect 582466 200784 582472 200796
rect 200080 200756 582472 200784
rect 200080 200744 200086 200756
rect 582466 200744 582472 200756
rect 582524 200744 582530 200796
rect 53466 200064 53472 200116
rect 53524 200104 53530 200116
rect 291378 200104 291384 200116
rect 53524 200076 291384 200104
rect 53524 200064 53530 200076
rect 291378 200064 291384 200076
rect 291436 200064 291442 200116
rect 53466 198704 53472 198756
rect 53524 198744 53530 198756
rect 53650 198744 53656 198756
rect 53524 198716 53656 198744
rect 53524 198704 53530 198716
rect 53650 198704 53656 198716
rect 53708 198704 53714 198756
rect 31754 197956 31760 198008
rect 31812 197996 31818 198008
rect 186958 197996 186964 198008
rect 31812 197968 186964 197996
rect 31812 197956 31818 197968
rect 186958 197956 186964 197968
rect 187016 197956 187022 198008
rect 255222 197956 255228 198008
rect 255280 197996 255286 198008
rect 280246 197996 280252 198008
rect 255280 197968 280252 197996
rect 255280 197956 255286 197968
rect 280246 197956 280252 197968
rect 280304 197956 280310 198008
rect 37274 196596 37280 196648
rect 37332 196636 37338 196648
rect 152642 196636 152648 196648
rect 37332 196608 152648 196636
rect 37332 196596 37338 196608
rect 152642 196596 152648 196608
rect 152700 196596 152706 196648
rect 123478 195304 123484 195356
rect 123536 195344 123542 195356
rect 140038 195344 140044 195356
rect 123536 195316 140044 195344
rect 123536 195304 123542 195316
rect 140038 195304 140044 195316
rect 140096 195304 140102 195356
rect 261478 195304 261484 195356
rect 261536 195344 261542 195356
rect 276198 195344 276204 195356
rect 261536 195316 276204 195344
rect 261536 195304 261542 195316
rect 276198 195304 276204 195316
rect 276256 195304 276262 195356
rect 97810 195236 97816 195288
rect 97868 195276 97874 195288
rect 123570 195276 123576 195288
rect 97868 195248 123576 195276
rect 97868 195236 97874 195248
rect 123570 195236 123576 195248
rect 123628 195236 123634 195288
rect 197354 195236 197360 195288
rect 197412 195276 197418 195288
rect 283098 195276 283104 195288
rect 197412 195248 283104 195276
rect 197412 195236 197418 195248
rect 283098 195236 283104 195248
rect 283156 195236 283162 195288
rect 108298 193808 108304 193860
rect 108356 193848 108362 193860
rect 129182 193848 129188 193860
rect 108356 193820 129188 193848
rect 108356 193808 108362 193820
rect 129182 193808 129188 193820
rect 129240 193808 129246 193860
rect 131758 193808 131764 193860
rect 131816 193848 131822 193860
rect 147030 193848 147036 193860
rect 131816 193820 147036 193848
rect 131816 193808 131822 193820
rect 147030 193808 147036 193820
rect 147088 193808 147094 193860
rect 148502 193808 148508 193860
rect 148560 193848 148566 193860
rect 162210 193848 162216 193860
rect 148560 193820 162216 193848
rect 148560 193808 148566 193820
rect 162210 193808 162216 193820
rect 162268 193808 162274 193860
rect 251910 192516 251916 192568
rect 251968 192556 251974 192568
rect 277578 192556 277584 192568
rect 251968 192528 277584 192556
rect 251968 192516 251974 192528
rect 277578 192516 277584 192528
rect 277636 192516 277642 192568
rect 187602 192448 187608 192500
rect 187660 192488 187666 192500
rect 228358 192488 228364 192500
rect 187660 192460 228364 192488
rect 187660 192448 187666 192460
rect 228358 192448 228364 192460
rect 228416 192448 228422 192500
rect 255958 192448 255964 192500
rect 256016 192488 256022 192500
rect 256602 192488 256608 192500
rect 256016 192460 256608 192488
rect 256016 192448 256022 192460
rect 256602 192448 256608 192460
rect 256660 192488 256666 192500
rect 580166 192488 580172 192500
rect 256660 192460 580172 192488
rect 256660 192448 256666 192460
rect 580166 192448 580172 192460
rect 580224 192448 580230 192500
rect 222930 191088 222936 191140
rect 222988 191128 222994 191140
rect 260926 191128 260932 191140
rect 222988 191100 260932 191128
rect 222988 191088 222994 191100
rect 260926 191088 260932 191100
rect 260984 191088 260990 191140
rect 80698 189728 80704 189780
rect 80756 189768 80762 189780
rect 145558 189768 145564 189780
rect 80756 189740 145564 189768
rect 80756 189728 80762 189740
rect 145558 189728 145564 189740
rect 145616 189728 145622 189780
rect 195238 189728 195244 189780
rect 195296 189768 195302 189780
rect 226610 189768 226616 189780
rect 195296 189740 226616 189768
rect 195296 189728 195302 189740
rect 226610 189728 226616 189740
rect 226668 189728 226674 189780
rect 61746 188300 61752 188352
rect 61804 188340 61810 188352
rect 71774 188340 71780 188352
rect 61804 188312 71780 188340
rect 61804 188300 61810 188312
rect 71774 188300 71780 188312
rect 71832 188300 71838 188352
rect 81342 188300 81348 188352
rect 81400 188340 81406 188352
rect 103514 188340 103520 188352
rect 81400 188312 103520 188340
rect 81400 188300 81406 188312
rect 103514 188300 103520 188312
rect 103572 188300 103578 188352
rect 114554 188300 114560 188352
rect 114612 188340 114618 188352
rect 131850 188340 131856 188352
rect 114612 188312 131856 188340
rect 114612 188300 114618 188312
rect 131850 188300 131856 188312
rect 131908 188300 131914 188352
rect 137370 188300 137376 188352
rect 137428 188340 137434 188352
rect 148410 188340 148416 188352
rect 137428 188312 148416 188340
rect 137428 188300 137434 188312
rect 148410 188300 148416 188312
rect 148468 188300 148474 188352
rect 175918 188300 175924 188352
rect 175976 188340 175982 188352
rect 185670 188340 185676 188352
rect 175976 188312 185676 188340
rect 175976 188300 175982 188312
rect 185670 188300 185676 188312
rect 185728 188300 185734 188352
rect 195790 188300 195796 188352
rect 195848 188340 195854 188352
rect 298094 188340 298100 188352
rect 195848 188312 298100 188340
rect 195848 188300 195854 188312
rect 298094 188300 298100 188312
rect 298152 188300 298158 188352
rect 145558 188096 145564 188148
rect 145616 188136 145622 188148
rect 154022 188136 154028 188148
rect 145616 188108 154028 188136
rect 145616 188096 145622 188108
rect 154022 188096 154028 188108
rect 154080 188096 154086 188148
rect 193122 187008 193128 187060
rect 193180 187048 193186 187060
rect 234614 187048 234620 187060
rect 193180 187020 234620 187048
rect 193180 187008 193186 187020
rect 234614 187008 234620 187020
rect 234672 187008 234678 187060
rect 9674 186940 9680 186992
rect 9732 186980 9738 186992
rect 186314 186980 186320 186992
rect 9732 186952 186320 186980
rect 9732 186940 9738 186952
rect 186314 186940 186320 186952
rect 186372 186940 186378 186992
rect 228358 186940 228364 186992
rect 228416 186980 228422 186992
rect 278866 186980 278872 186992
rect 228416 186952 278872 186980
rect 228416 186940 228422 186952
rect 278866 186940 278872 186952
rect 278924 186940 278930 186992
rect 202138 185580 202144 185632
rect 202196 185620 202202 185632
rect 243538 185620 243544 185632
rect 202196 185592 243544 185620
rect 202196 185580 202202 185592
rect 243538 185580 243544 185592
rect 243596 185580 243602 185632
rect 79318 184900 79324 184952
rect 79376 184940 79382 184952
rect 204254 184940 204260 184952
rect 79376 184912 204260 184940
rect 79376 184900 79382 184912
rect 204254 184900 204260 184912
rect 204312 184900 204318 184952
rect 73154 184220 73160 184272
rect 73212 184260 73218 184272
rect 91738 184260 91744 184272
rect 73212 184232 91744 184260
rect 73212 184220 73218 184232
rect 91738 184220 91744 184232
rect 91796 184220 91802 184272
rect 118786 184220 118792 184272
rect 118844 184260 118850 184272
rect 137462 184260 137468 184272
rect 118844 184232 137468 184260
rect 118844 184220 118850 184232
rect 137462 184220 137468 184232
rect 137520 184220 137526 184272
rect 89622 184152 89628 184204
rect 89680 184192 89686 184204
rect 126514 184192 126520 184204
rect 89680 184164 126520 184192
rect 89680 184152 89686 184164
rect 126514 184152 126520 184164
rect 126572 184152 126578 184204
rect 180150 184152 180156 184204
rect 180208 184192 180214 184204
rect 190454 184192 190460 184204
rect 180208 184164 190460 184192
rect 180208 184152 180214 184164
rect 190454 184152 190460 184164
rect 190512 184152 190518 184204
rect 196710 184152 196716 184204
rect 196768 184192 196774 184204
rect 218698 184192 218704 184204
rect 196768 184164 218704 184192
rect 196768 184152 196774 184164
rect 218698 184152 218704 184164
rect 218756 184152 218762 184204
rect 33778 182792 33784 182844
rect 33836 182832 33842 182844
rect 140130 182832 140136 182844
rect 33836 182804 140136 182832
rect 33836 182792 33842 182804
rect 140130 182792 140136 182804
rect 140188 182792 140194 182844
rect 86862 181500 86868 181552
rect 86920 181540 86926 181552
rect 117314 181540 117320 181552
rect 86920 181512 117320 181540
rect 86920 181500 86926 181512
rect 117314 181500 117320 181512
rect 117372 181500 117378 181552
rect 140038 181500 140044 181552
rect 140096 181540 140102 181552
rect 145650 181540 145656 181552
rect 140096 181512 145656 181540
rect 140096 181500 140102 181512
rect 145650 181500 145656 181512
rect 145708 181500 145714 181552
rect 63126 181432 63132 181484
rect 63184 181472 63190 181484
rect 180150 181472 180156 181484
rect 63184 181444 180156 181472
rect 63184 181432 63190 181444
rect 180150 181432 180156 181444
rect 180208 181432 180214 181484
rect 207750 181432 207756 181484
rect 207808 181472 207814 181484
rect 288526 181472 288532 181484
rect 207808 181444 288532 181472
rect 207808 181432 207814 181444
rect 288526 181432 288532 181444
rect 288584 181432 288590 181484
rect 88426 180072 88432 180124
rect 88484 180112 88490 180124
rect 116118 180112 116124 180124
rect 88484 180084 116124 180112
rect 88484 180072 88490 180084
rect 116118 180072 116124 180084
rect 116176 180072 116182 180124
rect 203518 180072 203524 180124
rect 203576 180112 203582 180124
rect 240226 180112 240232 180124
rect 203576 180084 240232 180112
rect 203576 180072 203582 180084
rect 240226 180072 240232 180084
rect 240284 180072 240290 180124
rect 52178 179392 52184 179444
rect 52236 179432 52242 179444
rect 167730 179432 167736 179444
rect 52236 179404 167736 179432
rect 52236 179392 52242 179404
rect 167730 179392 167736 179404
rect 167788 179392 167794 179444
rect 172422 179392 172428 179444
rect 172480 179432 172486 179444
rect 202874 179432 202880 179444
rect 172480 179404 202880 179432
rect 172480 179392 172486 179404
rect 202874 179392 202880 179404
rect 202932 179392 202938 179444
rect 87598 178644 87604 178696
rect 87656 178684 87662 178696
rect 105078 178684 105084 178696
rect 87656 178656 105084 178684
rect 87656 178644 87662 178656
rect 105078 178644 105084 178656
rect 105136 178644 105142 178696
rect 106918 178644 106924 178696
rect 106976 178684 106982 178696
rect 142982 178684 142988 178696
rect 106976 178656 142988 178684
rect 106976 178644 106982 178656
rect 142982 178644 142988 178656
rect 143040 178644 143046 178696
rect 182818 178644 182824 178696
rect 182876 178684 182882 178696
rect 227714 178684 227720 178696
rect 182876 178656 227720 178684
rect 182876 178644 182882 178656
rect 227714 178644 227720 178656
rect 227772 178644 227778 178696
rect 247678 178644 247684 178696
rect 247736 178684 247742 178696
rect 248322 178684 248328 178696
rect 247736 178656 248328 178684
rect 247736 178644 247742 178656
rect 248322 178644 248328 178656
rect 248380 178684 248386 178696
rect 580166 178684 580172 178696
rect 248380 178656 580172 178684
rect 248380 178644 248386 178656
rect 580166 178644 580172 178656
rect 580224 178644 580230 178696
rect 243538 178304 243544 178356
rect 243596 178344 243602 178356
rect 249886 178344 249892 178356
rect 243596 178316 249892 178344
rect 243596 178304 243602 178316
rect 249886 178304 249892 178316
rect 249944 178304 249950 178356
rect 190362 177284 190368 177336
rect 190420 177324 190426 177336
rect 274726 177324 274732 177336
rect 190420 177296 274732 177324
rect 190420 177284 190426 177296
rect 274726 177284 274732 177296
rect 274784 177284 274790 177336
rect 195974 175312 195980 175364
rect 196032 175352 196038 175364
rect 213178 175352 213184 175364
rect 196032 175324 213184 175352
rect 196032 175312 196038 175324
rect 213178 175312 213184 175324
rect 213236 175312 213242 175364
rect 113818 175244 113824 175296
rect 113876 175284 113882 175296
rect 204898 175284 204904 175296
rect 113876 175256 204904 175284
rect 113876 175244 113882 175256
rect 204898 175244 204904 175256
rect 204956 175244 204962 175296
rect 248966 175244 248972 175296
rect 249024 175284 249030 175296
rect 583018 175284 583024 175296
rect 249024 175256 583024 175284
rect 249024 175244 249030 175256
rect 583018 175244 583024 175256
rect 583076 175244 583082 175296
rect 150526 175176 150532 175228
rect 150584 175216 150590 175228
rect 195974 175216 195980 175228
rect 150584 175188 195980 175216
rect 150584 175176 150590 175188
rect 195974 175176 195980 175188
rect 196032 175176 196038 175228
rect 88334 174496 88340 174548
rect 88392 174536 88398 174548
rect 150526 174536 150532 174548
rect 88392 174508 150532 174536
rect 88392 174496 88398 174508
rect 150526 174496 150532 174508
rect 150584 174496 150590 174548
rect 154022 173884 154028 173936
rect 154080 173924 154086 173936
rect 220814 173924 220820 173936
rect 154080 173896 220820 173924
rect 154080 173884 154086 173896
rect 220814 173884 220820 173896
rect 220872 173924 220878 173936
rect 221458 173924 221464 173936
rect 220872 173896 221464 173924
rect 220872 173884 220878 173896
rect 221458 173884 221464 173896
rect 221516 173884 221522 173936
rect 222286 173816 222292 173868
rect 222344 173856 222350 173868
rect 222930 173856 222936 173868
rect 222344 173828 222936 173856
rect 222344 173816 222350 173828
rect 222930 173816 222936 173828
rect 222988 173816 222994 173868
rect 57698 173136 57704 173188
rect 57756 173176 57762 173188
rect 201586 173176 201592 173188
rect 57756 173148 201592 173176
rect 57756 173136 57762 173148
rect 201586 173136 201592 173148
rect 201644 173176 201650 173188
rect 202138 173176 202144 173188
rect 201644 173148 202144 173176
rect 201644 173136 201650 173148
rect 202138 173136 202144 173148
rect 202196 173136 202202 173188
rect 227990 173136 227996 173188
rect 228048 173176 228054 173188
rect 251818 173176 251824 173188
rect 228048 173148 251824 173176
rect 228048 173136 228054 173148
rect 251818 173136 251824 173148
rect 251876 173176 251882 173188
rect 341518 173176 341524 173188
rect 251876 173148 341524 173176
rect 251876 173136 251882 173148
rect 341518 173136 341524 173148
rect 341576 173136 341582 173188
rect 87138 172524 87144 172576
rect 87196 172564 87202 172576
rect 222286 172564 222292 172576
rect 87196 172536 222292 172564
rect 87196 172524 87202 172536
rect 222286 172524 222292 172536
rect 222344 172524 222350 172576
rect 205818 172456 205824 172508
rect 205876 172496 205882 172508
rect 303614 172496 303620 172508
rect 205876 172468 303620 172496
rect 205876 172456 205882 172468
rect 303614 172456 303620 172468
rect 303672 172496 303678 172508
rect 304074 172496 304080 172508
rect 303672 172468 304080 172496
rect 303672 172456 303678 172468
rect 304074 172456 304080 172468
rect 304132 172456 304138 172508
rect 304074 171776 304080 171828
rect 304132 171816 304138 171828
rect 320174 171816 320180 171828
rect 304132 171788 320180 171816
rect 304132 171776 304138 171788
rect 320174 171776 320180 171788
rect 320232 171776 320238 171828
rect 92658 171096 92664 171148
rect 92716 171136 92722 171148
rect 222838 171136 222844 171148
rect 92716 171108 222844 171136
rect 92716 171096 92722 171108
rect 222838 171096 222844 171108
rect 222896 171096 222902 171148
rect 91186 170348 91192 170400
rect 91244 170388 91250 170400
rect 154022 170388 154028 170400
rect 91244 170360 154028 170388
rect 91244 170348 91250 170360
rect 154022 170348 154028 170360
rect 154080 170348 154086 170400
rect 154390 169804 154396 169856
rect 154448 169844 154454 169856
rect 154448 169816 213960 169844
rect 154448 169804 154454 169816
rect 213932 169788 213960 169816
rect 86218 169736 86224 169788
rect 86276 169776 86282 169788
rect 86276 169748 213868 169776
rect 86276 169736 86282 169748
rect 213840 169708 213868 169748
rect 213914 169736 213920 169788
rect 213972 169776 213978 169788
rect 214558 169776 214564 169788
rect 213972 169748 214564 169776
rect 213972 169736 213978 169748
rect 214558 169736 214564 169748
rect 214616 169736 214622 169788
rect 216858 169776 216864 169788
rect 214668 169748 216864 169776
rect 214668 169708 214696 169748
rect 216858 169736 216864 169748
rect 216916 169776 216922 169788
rect 217962 169776 217968 169788
rect 216916 169748 217968 169776
rect 216916 169736 216922 169748
rect 217962 169736 217968 169748
rect 218020 169776 218026 169788
rect 582742 169776 582748 169788
rect 218020 169748 582748 169776
rect 218020 169736 218026 169748
rect 582742 169736 582748 169748
rect 582800 169736 582806 169788
rect 213840 169680 214696 169708
rect 134702 168444 134708 168496
rect 134760 168484 134766 168496
rect 227990 168484 227996 168496
rect 134760 168456 227996 168484
rect 134760 168444 134766 168456
rect 227990 168444 227996 168456
rect 228048 168444 228054 168496
rect 73338 168376 73344 168428
rect 73396 168416 73402 168428
rect 73396 168388 200114 168416
rect 73396 168376 73402 168388
rect 200086 168348 200114 168388
rect 200298 168348 200304 168360
rect 200086 168320 200304 168348
rect 200298 168308 200304 168320
rect 200356 168348 200362 168360
rect 254026 168348 254032 168360
rect 200356 168320 254032 168348
rect 200356 168308 200362 168320
rect 254026 168308 254032 168320
rect 254084 168308 254090 168360
rect 192570 167124 192576 167136
rect 74506 167096 192576 167124
rect 67726 167016 67732 167068
rect 67784 167056 67790 167068
rect 68922 167056 68928 167068
rect 67784 167028 68928 167056
rect 67784 167016 67790 167028
rect 68922 167016 68928 167028
rect 68980 167056 68986 167068
rect 74506 167056 74534 167096
rect 192570 167084 192576 167096
rect 192628 167084 192634 167136
rect 68980 167028 74534 167056
rect 68980 167016 68986 167028
rect 101398 167016 101404 167068
rect 101456 167056 101462 167068
rect 101582 167056 101588 167068
rect 101456 167028 101588 167056
rect 101456 167016 101462 167028
rect 101582 167016 101588 167028
rect 101640 167056 101646 167068
rect 233234 167056 233240 167068
rect 101640 167028 233240 167056
rect 101640 167016 101646 167028
rect 233234 167016 233240 167028
rect 233292 167016 233298 167068
rect 63218 166268 63224 166320
rect 63276 166308 63282 166320
rect 164050 166308 164056 166320
rect 63276 166280 164056 166308
rect 63276 166268 63282 166280
rect 164050 166268 164056 166280
rect 164108 166308 164114 166320
rect 190454 166308 190460 166320
rect 164108 166280 190460 166308
rect 164108 166268 164114 166280
rect 190454 166268 190460 166280
rect 190512 166268 190518 166320
rect 198734 166268 198740 166320
rect 198792 166308 198798 166320
rect 263594 166308 263600 166320
rect 198792 166280 263600 166308
rect 198792 166268 198798 166280
rect 263594 166268 263600 166280
rect 263652 166268 263658 166320
rect 90358 165588 90364 165640
rect 90416 165628 90422 165640
rect 208394 165628 208400 165640
rect 90416 165600 208400 165628
rect 90416 165588 90422 165600
rect 208394 165588 208400 165600
rect 208452 165588 208458 165640
rect 154482 164908 154488 164960
rect 154540 164948 154546 164960
rect 195790 164948 195796 164960
rect 154540 164920 195796 164948
rect 154540 164908 154546 164920
rect 195790 164908 195796 164920
rect 195848 164948 195854 164960
rect 197538 164948 197544 164960
rect 195848 164920 197544 164948
rect 195848 164908 195854 164920
rect 197538 164908 197544 164920
rect 197596 164908 197602 164960
rect 60458 164840 60464 164892
rect 60516 164880 60522 164892
rect 83458 164880 83464 164892
rect 60516 164852 83464 164880
rect 60516 164840 60522 164852
rect 83458 164840 83464 164852
rect 83516 164840 83522 164892
rect 193858 164840 193864 164892
rect 193916 164880 193922 164892
rect 262582 164880 262588 164892
rect 193916 164852 262588 164880
rect 193916 164840 193922 164852
rect 262582 164840 262588 164852
rect 262640 164840 262646 164892
rect 210418 164160 210424 164212
rect 210476 164200 210482 164212
rect 293954 164200 293960 164212
rect 210476 164172 293960 164200
rect 210476 164160 210482 164172
rect 293954 164160 293960 164172
rect 294012 164200 294018 164212
rect 294414 164200 294420 164212
rect 294012 164172 294420 164200
rect 294012 164160 294018 164172
rect 294414 164160 294420 164172
rect 294472 164160 294478 164212
rect 82906 163548 82912 163600
rect 82964 163588 82970 163600
rect 154390 163588 154396 163600
rect 82964 163560 154396 163588
rect 82964 163548 82970 163560
rect 154390 163548 154396 163560
rect 154448 163548 154454 163600
rect 88978 163480 88984 163532
rect 89036 163520 89042 163532
rect 169754 163520 169760 163532
rect 89036 163492 169760 163520
rect 89036 163480 89042 163492
rect 169754 163480 169760 163492
rect 169812 163520 169818 163532
rect 196802 163520 196808 163532
rect 169812 163492 196808 163520
rect 169812 163480 169818 163492
rect 196802 163480 196808 163492
rect 196860 163480 196866 163532
rect 294414 163480 294420 163532
rect 294472 163520 294478 163532
rect 582926 163520 582932 163532
rect 294472 163492 582932 163520
rect 294472 163480 294478 163492
rect 582926 163480 582932 163492
rect 582984 163480 582990 163532
rect 208394 162800 208400 162852
rect 208452 162840 208458 162852
rect 270678 162840 270684 162852
rect 208452 162812 270684 162840
rect 208452 162800 208458 162812
rect 270678 162800 270684 162812
rect 270736 162800 270742 162852
rect 222194 161848 222200 161900
rect 222252 161888 222258 161900
rect 222930 161888 222936 161900
rect 222252 161860 222936 161888
rect 222252 161848 222258 161860
rect 222930 161848 222936 161860
rect 222988 161848 222994 161900
rect 152642 161508 152648 161560
rect 152700 161548 152706 161560
rect 222194 161548 222200 161560
rect 152700 161520 222200 161548
rect 152700 161508 152706 161520
rect 222194 161508 222200 161520
rect 222252 161508 222258 161560
rect 73062 161440 73068 161492
rect 73120 161480 73126 161492
rect 198734 161480 198740 161492
rect 73120 161452 198740 161480
rect 73120 161440 73126 161452
rect 198734 161440 198740 161452
rect 198792 161440 198798 161492
rect 234614 160692 234620 160744
rect 234672 160732 234678 160744
rect 259546 160732 259552 160744
rect 234672 160704 259552 160732
rect 234672 160692 234678 160704
rect 259546 160692 259552 160704
rect 259604 160692 259610 160744
rect 156782 160148 156788 160200
rect 156840 160188 156846 160200
rect 157242 160188 157248 160200
rect 156840 160160 157248 160188
rect 156840 160148 156846 160160
rect 157242 160148 157248 160160
rect 157300 160188 157306 160200
rect 224218 160188 224224 160200
rect 157300 160160 224224 160188
rect 157300 160148 157306 160160
rect 224218 160148 224224 160160
rect 224276 160148 224282 160200
rect 64598 160080 64604 160132
rect 64656 160120 64662 160132
rect 165062 160120 165068 160132
rect 64656 160092 165068 160120
rect 64656 160080 64662 160092
rect 165062 160080 165068 160092
rect 165120 160080 165126 160132
rect 194594 160080 194600 160132
rect 194652 160120 194658 160132
rect 195882 160120 195888 160132
rect 194652 160092 195888 160120
rect 194652 160080 194658 160092
rect 195882 160080 195888 160092
rect 195940 160120 195946 160132
rect 276658 160120 276664 160132
rect 195940 160092 276664 160120
rect 195940 160080 195946 160092
rect 276658 160080 276664 160092
rect 276716 160080 276722 160132
rect 242894 159468 242900 159520
rect 242952 159508 242958 159520
rect 243538 159508 243544 159520
rect 242952 159480 243544 159508
rect 242952 159468 242958 159480
rect 243538 159468 243544 159480
rect 243596 159468 243602 159520
rect 119338 159332 119344 159384
rect 119396 159372 119402 159384
rect 242894 159372 242900 159384
rect 119396 159344 242900 159372
rect 119396 159332 119402 159344
rect 242894 159332 242900 159344
rect 242952 159332 242958 159384
rect 249058 159332 249064 159384
rect 249116 159372 249122 159384
rect 261202 159372 261208 159384
rect 249116 159344 261208 159372
rect 249116 159332 249122 159344
rect 261202 159332 261208 159344
rect 261260 159332 261266 159384
rect 91830 158720 91836 158772
rect 91888 158760 91894 158772
rect 92382 158760 92388 158772
rect 91888 158732 92388 158760
rect 91888 158720 91894 158732
rect 92382 158720 92388 158732
rect 92440 158760 92446 158772
rect 220814 158760 220820 158772
rect 92440 158732 220820 158760
rect 92440 158720 92446 158732
rect 220814 158720 220820 158732
rect 220872 158720 220878 158772
rect 65978 157972 65984 158024
rect 66036 158012 66042 158024
rect 182818 158012 182824 158024
rect 66036 157984 182824 158012
rect 66036 157972 66042 157984
rect 182818 157972 182824 157984
rect 182876 157972 182882 158024
rect 202782 157972 202788 158024
rect 202840 158012 202846 158024
rect 267734 158012 267740 158024
rect 202840 157984 267740 158012
rect 202840 157972 202846 157984
rect 267734 157972 267740 157984
rect 267792 157972 267798 158024
rect 105538 157360 105544 157412
rect 105596 157400 105602 157412
rect 225046 157400 225052 157412
rect 105596 157372 225052 157400
rect 105596 157360 105602 157372
rect 225046 157360 225052 157372
rect 225104 157360 225110 157412
rect 53558 156612 53564 156664
rect 53616 156652 53622 156664
rect 67818 156652 67824 156664
rect 53616 156624 67824 156652
rect 53616 156612 53622 156624
rect 67818 156612 67824 156624
rect 67876 156652 67882 156664
rect 68646 156652 68652 156664
rect 67876 156624 68652 156652
rect 67876 156612 67882 156624
rect 68646 156612 68652 156624
rect 68704 156612 68710 156664
rect 196618 156612 196624 156664
rect 196676 156652 196682 156664
rect 205726 156652 205732 156664
rect 196676 156624 205732 156652
rect 196676 156612 196682 156624
rect 205726 156612 205732 156624
rect 205784 156612 205790 156664
rect 97258 156408 97264 156460
rect 97316 156448 97322 156460
rect 97902 156448 97908 156460
rect 97316 156420 97908 156448
rect 97316 156408 97322 156420
rect 97902 156408 97908 156420
rect 97960 156408 97966 156460
rect 247034 156408 247040 156460
rect 247092 156448 247098 156460
rect 247678 156448 247684 156460
rect 247092 156420 247684 156448
rect 247092 156408 247098 156420
rect 247678 156408 247684 156420
rect 247736 156408 247742 156460
rect 68646 156000 68652 156052
rect 68704 156040 68710 156052
rect 189902 156040 189908 156052
rect 68704 156012 189908 156040
rect 68704 156000 68710 156012
rect 189902 156000 189908 156012
rect 189960 156000 189966 156052
rect 207106 156000 207112 156052
rect 207164 156040 207170 156052
rect 247034 156040 247040 156052
rect 207164 156012 247040 156040
rect 207164 156000 207170 156012
rect 247034 156000 247040 156012
rect 247092 156000 247098 156052
rect 97902 155932 97908 155984
rect 97960 155972 97966 155984
rect 226426 155972 226432 155984
rect 97960 155944 226432 155972
rect 97960 155932 97966 155944
rect 226426 155932 226432 155944
rect 226484 155932 226490 155984
rect 56226 155864 56232 155916
rect 56284 155904 56290 155916
rect 56502 155904 56508 155916
rect 56284 155876 56508 155904
rect 56284 155864 56290 155876
rect 56502 155864 56508 155876
rect 56560 155864 56566 155916
rect 215386 155184 215392 155236
rect 215444 155224 215450 155236
rect 222286 155224 222292 155236
rect 215444 155196 222292 155224
rect 215444 155184 215450 155196
rect 222286 155184 222292 155196
rect 222344 155184 222350 155236
rect 263594 155184 263600 155236
rect 263652 155224 263658 155236
rect 299474 155224 299480 155236
rect 263652 155196 299480 155224
rect 263652 155184 263658 155196
rect 299474 155184 299480 155196
rect 299532 155184 299538 155236
rect 204346 154912 204352 154964
rect 204404 154952 204410 154964
rect 204898 154952 204904 154964
rect 204404 154924 204904 154952
rect 204404 154912 204410 154924
rect 204898 154912 204904 154924
rect 204956 154912 204962 154964
rect 56502 154640 56508 154692
rect 56560 154680 56566 154692
rect 137462 154680 137468 154692
rect 56560 154652 137468 154680
rect 56560 154640 56566 154652
rect 137462 154640 137468 154652
rect 137520 154640 137526 154692
rect 91922 154572 91928 154624
rect 91980 154612 91986 154624
rect 201678 154612 201684 154624
rect 91980 154584 201684 154612
rect 91980 154572 91986 154584
rect 201678 154572 201684 154584
rect 201736 154612 201742 154624
rect 202782 154612 202788 154624
rect 201736 154584 202788 154612
rect 201736 154572 201742 154584
rect 202782 154572 202788 154584
rect 202840 154572 202846 154624
rect 204898 154572 204904 154624
rect 204956 154612 204962 154624
rect 263594 154612 263600 154624
rect 204956 154584 263600 154612
rect 204956 154572 204962 154584
rect 263594 154572 263600 154584
rect 263652 154572 263658 154624
rect 222194 154504 222200 154556
rect 222252 154544 222258 154556
rect 282914 154544 282920 154556
rect 222252 154516 282920 154544
rect 222252 154504 222258 154516
rect 282914 154504 282920 154516
rect 282972 154504 282978 154556
rect 189166 153824 189172 153876
rect 189224 153864 189230 153876
rect 201494 153864 201500 153876
rect 189224 153836 201500 153864
rect 189224 153824 189230 153836
rect 201494 153824 201500 153836
rect 201552 153824 201558 153876
rect 237374 153824 237380 153876
rect 237432 153864 237438 153876
rect 265618 153864 265624 153876
rect 237432 153836 265624 153864
rect 237432 153824 237438 153836
rect 265618 153824 265624 153836
rect 265676 153864 265682 153876
rect 342254 153864 342260 153876
rect 265676 153836 342260 153864
rect 265676 153824 265682 153836
rect 342254 153824 342260 153836
rect 342312 153824 342318 153876
rect 67266 153280 67272 153332
rect 67324 153320 67330 153332
rect 112438 153320 112444 153332
rect 67324 153292 112444 153320
rect 67324 153280 67330 153292
rect 112438 153280 112444 153292
rect 112496 153280 112502 153332
rect 129090 153280 129096 153332
rect 129148 153320 129154 153332
rect 223574 153320 223580 153332
rect 129148 153292 223580 153320
rect 129148 153280 129154 153292
rect 223574 153280 223580 153292
rect 223632 153280 223638 153332
rect 49510 153212 49516 153264
rect 49568 153252 49574 153264
rect 186222 153252 186228 153264
rect 49568 153224 186228 153252
rect 49568 153212 49574 153224
rect 186222 153212 186228 153224
rect 186280 153212 186286 153264
rect 211154 153144 211160 153196
rect 211212 153184 211218 153196
rect 271874 153184 271880 153196
rect 211212 153156 271880 153184
rect 211212 153144 211218 153156
rect 271874 153144 271880 153156
rect 271932 153144 271938 153196
rect 192570 153076 192576 153128
rect 192628 153116 192634 153128
rect 237374 153116 237380 153128
rect 192628 153088 237380 153116
rect 192628 153076 192634 153088
rect 237374 153076 237380 153088
rect 237432 153076 237438 153128
rect 92750 152532 92756 152584
rect 92808 152572 92814 152584
rect 154482 152572 154488 152584
rect 92808 152544 154488 152572
rect 92808 152532 92814 152544
rect 154482 152532 154488 152544
rect 154540 152532 154546 152584
rect 133230 152464 133236 152516
rect 133288 152504 133294 152516
rect 207106 152504 207112 152516
rect 133288 152476 207112 152504
rect 133288 152464 133294 152476
rect 207106 152464 207112 152476
rect 207164 152464 207170 152516
rect 54938 151784 54944 151836
rect 54996 151824 55002 151836
rect 127710 151824 127716 151836
rect 54996 151796 127716 151824
rect 54996 151784 55002 151796
rect 127710 151784 127716 151796
rect 127768 151784 127774 151836
rect 80054 151104 80060 151156
rect 80112 151144 80118 151156
rect 90358 151144 90364 151156
rect 80112 151116 90364 151144
rect 80112 151104 80118 151116
rect 90358 151104 90364 151116
rect 90416 151104 90422 151156
rect 57790 151036 57796 151088
rect 57848 151076 57854 151088
rect 189166 151076 189172 151088
rect 57848 151048 189172 151076
rect 57848 151036 57854 151048
rect 189166 151036 189172 151048
rect 189224 151036 189230 151088
rect 170490 150492 170496 150544
rect 170548 150532 170554 150544
rect 224954 150532 224960 150544
rect 170548 150504 224960 150532
rect 170548 150492 170554 150504
rect 224954 150492 224960 150504
rect 225012 150492 225018 150544
rect 189166 150424 189172 150476
rect 189224 150464 189230 150476
rect 189810 150464 189816 150476
rect 189224 150436 189816 150464
rect 189224 150424 189230 150436
rect 189810 150424 189816 150436
rect 189868 150424 189874 150476
rect 218238 150424 218244 150476
rect 218296 150464 218302 150476
rect 323578 150464 323584 150476
rect 218296 150436 323584 150464
rect 218296 150424 218302 150436
rect 323578 150424 323584 150436
rect 323636 150424 323642 150476
rect 197354 149948 197360 150000
rect 197412 149988 197418 150000
rect 197630 149988 197636 150000
rect 197412 149960 197636 149988
rect 197412 149948 197418 149960
rect 197630 149948 197636 149960
rect 197688 149948 197694 150000
rect 191098 149812 191104 149864
rect 191156 149852 191162 149864
rect 224862 149852 224868 149864
rect 191156 149824 224868 149852
rect 191156 149812 191162 149824
rect 224862 149812 224868 149824
rect 224920 149812 224926 149864
rect 81986 149744 81992 149796
rect 82044 149784 82050 149796
rect 102134 149784 102140 149796
rect 82044 149756 102140 149784
rect 82044 149744 82050 149756
rect 102134 149744 102140 149756
rect 102192 149744 102198 149796
rect 218330 149744 218336 149796
rect 218388 149784 218394 149796
rect 268102 149784 268108 149796
rect 218388 149756 268108 149784
rect 218388 149744 218394 149756
rect 268102 149744 268108 149756
rect 268160 149744 268166 149796
rect 70302 149676 70308 149728
rect 70360 149716 70366 149728
rect 77938 149716 77944 149728
rect 70360 149688 77944 149716
rect 70360 149676 70366 149688
rect 77938 149676 77944 149688
rect 77996 149676 78002 149728
rect 86862 149676 86868 149728
rect 86920 149716 86926 149728
rect 126330 149716 126336 149728
rect 86920 149688 126336 149716
rect 86920 149676 86926 149688
rect 126330 149676 126336 149688
rect 126388 149716 126394 149728
rect 216674 149716 216680 149728
rect 126388 149688 216680 149716
rect 126388 149676 126394 149688
rect 216674 149676 216680 149688
rect 216732 149676 216738 149728
rect 224862 149676 224868 149728
rect 224920 149716 224926 149728
rect 305638 149716 305644 149728
rect 224920 149688 305644 149716
rect 224920 149676 224926 149688
rect 305638 149676 305644 149688
rect 305696 149676 305702 149728
rect 82814 149472 82820 149524
rect 82872 149512 82878 149524
rect 86310 149512 86316 149524
rect 82872 149484 86316 149512
rect 82872 149472 82878 149484
rect 86310 149472 86316 149484
rect 86368 149472 86374 149524
rect 230014 148996 230020 149048
rect 230072 149036 230078 149048
rect 276014 149036 276020 149048
rect 230072 149008 276020 149036
rect 230072 148996 230078 149008
rect 276014 148996 276020 149008
rect 276072 148996 276078 149048
rect 220906 148424 220912 148436
rect 132466 148396 220912 148424
rect 52454 148316 52460 148368
rect 52512 148356 52518 148368
rect 80698 148356 80704 148368
rect 52512 148328 80704 148356
rect 52512 148316 52518 148328
rect 80698 148316 80704 148328
rect 80756 148316 80762 148368
rect 91002 148316 91008 148368
rect 91060 148356 91066 148368
rect 127618 148356 127624 148368
rect 91060 148328 127624 148356
rect 91060 148316 91066 148328
rect 127618 148316 127624 148328
rect 127676 148356 127682 148368
rect 132466 148356 132494 148396
rect 220906 148384 220912 148396
rect 220964 148384 220970 148436
rect 127676 148328 132494 148356
rect 127676 148316 127682 148328
rect 186222 148316 186228 148368
rect 186280 148356 186286 148368
rect 188798 148356 188804 148368
rect 186280 148328 188804 148356
rect 186280 148316 186286 148328
rect 188798 148316 188804 148328
rect 188856 148356 188862 148368
rect 196710 148356 196716 148368
rect 188856 148328 196716 148356
rect 188856 148316 188862 148328
rect 196710 148316 196716 148328
rect 196768 148316 196774 148368
rect 213914 148316 213920 148368
rect 213972 148356 213978 148368
rect 317414 148356 317420 148368
rect 213972 148328 317420 148356
rect 213972 148316 213978 148328
rect 317414 148316 317420 148328
rect 317472 148316 317478 148368
rect 57882 147636 57888 147688
rect 57940 147676 57946 147688
rect 184290 147676 184296 147688
rect 57940 147648 184296 147676
rect 57940 147636 57946 147648
rect 184290 147636 184296 147648
rect 184348 147636 184354 147688
rect 211890 147636 211896 147688
rect 211948 147676 211954 147688
rect 213914 147676 213920 147688
rect 211948 147648 213920 147676
rect 211948 147636 211954 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 97810 147092 97816 147144
rect 97868 147132 97874 147144
rect 101398 147132 101404 147144
rect 97868 147104 101404 147132
rect 97868 147092 97874 147104
rect 101398 147092 101404 147104
rect 101456 147092 101462 147144
rect 215386 146956 215392 147008
rect 215444 146996 215450 147008
rect 216214 146996 216220 147008
rect 215444 146968 216220 146996
rect 215444 146956 215450 146968
rect 216214 146956 216220 146968
rect 216272 146956 216278 147008
rect 4246 146888 4252 146940
rect 4304 146928 4310 146940
rect 97442 146928 97448 146940
rect 4304 146900 97448 146928
rect 4304 146888 4310 146900
rect 97442 146888 97448 146900
rect 97500 146888 97506 146940
rect 255314 146752 255320 146804
rect 255372 146792 255378 146804
rect 256050 146792 256056 146804
rect 255372 146764 256056 146792
rect 255372 146752 255378 146764
rect 256050 146752 256056 146764
rect 256108 146752 256114 146804
rect 113910 146344 113916 146396
rect 113968 146384 113974 146396
rect 227806 146384 227812 146396
rect 113968 146356 227812 146384
rect 113968 146344 113974 146356
rect 227806 146344 227812 146356
rect 227864 146344 227870 146396
rect 80514 146276 80520 146328
rect 80572 146316 80578 146328
rect 208486 146316 208492 146328
rect 80572 146288 208492 146316
rect 80572 146276 80578 146288
rect 208486 146276 208492 146288
rect 208544 146276 208550 146328
rect 214558 146276 214564 146328
rect 214616 146316 214622 146328
rect 255314 146316 255320 146328
rect 214616 146288 255320 146316
rect 214616 146276 214622 146288
rect 255314 146276 255320 146288
rect 255372 146276 255378 146328
rect 3418 146208 3424 146260
rect 3476 146248 3482 146260
rect 86862 146248 86868 146260
rect 3476 146220 86868 146248
rect 3476 146208 3482 146220
rect 86862 146208 86868 146220
rect 86920 146208 86926 146260
rect 213178 146208 213184 146260
rect 213236 146248 213242 146260
rect 216766 146248 216772 146260
rect 213236 146220 216772 146248
rect 213236 146208 213242 146220
rect 216766 146208 216772 146220
rect 216824 146208 216830 146260
rect 94314 145596 94320 145648
rect 94372 145636 94378 145648
rect 129090 145636 129096 145648
rect 94372 145608 129096 145636
rect 94372 145596 94378 145608
rect 129090 145596 129096 145608
rect 129148 145596 129154 145648
rect 252830 145596 252836 145648
rect 252888 145636 252894 145648
rect 327074 145636 327080 145648
rect 252888 145608 327080 145636
rect 252888 145596 252894 145608
rect 327074 145596 327080 145608
rect 327132 145596 327138 145648
rect 71774 145528 71780 145580
rect 71832 145568 71838 145580
rect 107562 145568 107568 145580
rect 71832 145540 107568 145568
rect 71832 145528 71838 145540
rect 107562 145528 107568 145540
rect 107620 145568 107626 145580
rect 197998 145568 198004 145580
rect 107620 145540 198004 145568
rect 107620 145528 107626 145540
rect 197998 145528 198004 145540
rect 198056 145528 198062 145580
rect 198826 145528 198832 145580
rect 198884 145568 198890 145580
rect 287238 145568 287244 145580
rect 198884 145540 287244 145568
rect 198884 145528 198890 145540
rect 287238 145528 287244 145540
rect 287296 145528 287302 145580
rect 86862 144916 86868 144968
rect 86920 144956 86926 144968
rect 87690 144956 87696 144968
rect 86920 144928 87696 144956
rect 86920 144916 86926 144928
rect 87690 144916 87696 144928
rect 87748 144916 87754 144968
rect 177298 144916 177304 144968
rect 177356 144956 177362 144968
rect 209866 144956 209872 144968
rect 177356 144928 209872 144956
rect 177356 144916 177362 144928
rect 209866 144916 209872 144928
rect 209924 144916 209930 144968
rect 222930 144848 222936 144900
rect 222988 144888 222994 144900
rect 226518 144888 226524 144900
rect 222988 144860 226524 144888
rect 222988 144848 222994 144860
rect 226518 144848 226524 144860
rect 226576 144848 226582 144900
rect 200206 144440 200212 144492
rect 200264 144480 200270 144492
rect 207750 144480 207756 144492
rect 200264 144452 207756 144480
rect 200264 144440 200270 144452
rect 207750 144440 207756 144452
rect 207808 144440 207814 144492
rect 78674 144372 78680 144424
rect 78732 144412 78738 144424
rect 82170 144412 82176 144424
rect 78732 144384 82176 144412
rect 78732 144372 78738 144384
rect 82170 144372 82176 144384
rect 82228 144372 82234 144424
rect 102318 144168 102324 144220
rect 102376 144208 102382 144220
rect 184198 144208 184204 144220
rect 102376 144180 184204 144208
rect 102376 144168 102382 144180
rect 184198 144168 184204 144180
rect 184256 144168 184262 144220
rect 188430 144168 188436 144220
rect 188488 144208 188494 144220
rect 196526 144208 196532 144220
rect 188488 144180 196532 144208
rect 188488 144168 188494 144180
rect 196526 144168 196532 144180
rect 196584 144168 196590 144220
rect 206830 144168 206836 144220
rect 206888 144208 206894 144220
rect 284938 144208 284944 144220
rect 206888 144180 284944 144208
rect 206888 144168 206894 144180
rect 284938 144168 284944 144180
rect 284996 144208 285002 144220
rect 298738 144208 298744 144220
rect 284996 144180 298744 144208
rect 284996 144168 285002 144180
rect 298738 144168 298744 144180
rect 298796 144168 298802 144220
rect 202046 143664 202052 143676
rect 180766 143636 202052 143664
rect 53650 143556 53656 143608
rect 53708 143596 53714 143608
rect 153930 143596 153936 143608
rect 53708 143568 153936 143596
rect 53708 143556 53714 143568
rect 153930 143556 153936 143568
rect 153988 143556 153994 143608
rect 169662 143556 169668 143608
rect 169720 143596 169726 143608
rect 180766 143596 180794 143636
rect 202046 143624 202052 143636
rect 202104 143624 202110 143676
rect 169720 143568 180794 143596
rect 169720 143556 169726 143568
rect 196802 143556 196808 143608
rect 196860 143596 196866 143608
rect 201310 143596 201316 143608
rect 196860 143568 201316 143596
rect 196860 143556 196866 143568
rect 201310 143556 201316 143568
rect 201368 143556 201374 143608
rect 214006 143488 214012 143540
rect 214064 143528 214070 143540
rect 216858 143528 216864 143540
rect 214064 143500 216864 143528
rect 214064 143488 214070 143500
rect 216858 143488 216864 143500
rect 216916 143488 216922 143540
rect 219526 143488 219532 143540
rect 219584 143528 219590 143540
rect 220078 143528 220084 143540
rect 219584 143500 220084 143528
rect 219584 143488 219590 143500
rect 220078 143488 220084 143500
rect 220136 143488 220142 143540
rect 82906 142808 82912 142860
rect 82964 142848 82970 142860
rect 83550 142848 83556 142860
rect 82964 142820 83556 142848
rect 82964 142808 82970 142820
rect 83550 142808 83556 142820
rect 83608 142808 83614 142860
rect 88426 142264 88432 142316
rect 88484 142304 88490 142316
rect 213270 142304 213276 142316
rect 88484 142276 213276 142304
rect 88484 142264 88490 142276
rect 213270 142264 213276 142276
rect 213328 142264 213334 142316
rect 189074 142196 189080 142248
rect 189132 142236 189138 142248
rect 206830 142236 206836 142248
rect 189132 142208 206836 142236
rect 189132 142196 189138 142208
rect 206830 142196 206836 142208
rect 206888 142196 206894 142248
rect 215294 142196 215300 142248
rect 215352 142236 215358 142248
rect 221458 142236 221464 142248
rect 215352 142208 221464 142236
rect 215352 142196 215358 142208
rect 221458 142196 221464 142208
rect 221516 142196 221522 142248
rect 223206 142196 223212 142248
rect 223264 142236 223270 142248
rect 223264 142208 229094 142236
rect 223264 142196 223270 142208
rect 211798 142128 211804 142180
rect 211856 142168 211862 142180
rect 212810 142168 212816 142180
rect 211856 142140 212816 142168
rect 211856 142128 211862 142140
rect 212810 142128 212816 142140
rect 212868 142128 212874 142180
rect 219986 142128 219992 142180
rect 220044 142168 220050 142180
rect 225598 142168 225604 142180
rect 220044 142140 225604 142168
rect 220044 142128 220050 142140
rect 225598 142128 225604 142140
rect 225656 142128 225662 142180
rect 229066 142168 229094 142208
rect 240778 142168 240784 142180
rect 229066 142140 240784 142168
rect 240778 142128 240784 142140
rect 240836 142128 240842 142180
rect 76282 141380 76288 141432
rect 76340 141420 76346 141432
rect 159450 141420 159456 141432
rect 76340 141392 159456 141420
rect 76340 141380 76346 141392
rect 159450 141380 159456 141392
rect 159508 141420 159514 141432
rect 203150 141420 203156 141432
rect 159508 141392 203156 141420
rect 159508 141380 159514 141392
rect 203150 141380 203156 141392
rect 203208 141380 203214 141432
rect 218790 141380 218796 141432
rect 218848 141420 218854 141432
rect 227898 141420 227904 141432
rect 218848 141392 227904 141420
rect 218848 141380 218854 141392
rect 227898 141380 227904 141392
rect 227956 141380 227962 141432
rect 223574 141176 223580 141228
rect 223632 141216 223638 141228
rect 224494 141216 224500 141228
rect 223632 141188 224500 141216
rect 223632 141176 223638 141188
rect 224494 141176 224500 141188
rect 224552 141176 224558 141228
rect 65886 140836 65892 140888
rect 65944 140876 65950 140888
rect 70486 140876 70492 140888
rect 65944 140848 70492 140876
rect 65944 140836 65950 140848
rect 70486 140836 70492 140848
rect 70544 140836 70550 140888
rect 214374 140876 214380 140888
rect 193324 140848 214380 140876
rect 58986 140768 58992 140820
rect 59044 140808 59050 140820
rect 59262 140808 59268 140820
rect 59044 140780 59268 140808
rect 59044 140768 59050 140780
rect 59262 140768 59268 140780
rect 59320 140808 59326 140820
rect 105630 140808 105636 140820
rect 59320 140780 105636 140808
rect 59320 140768 59326 140780
rect 105630 140768 105636 140780
rect 105688 140768 105694 140820
rect 186314 140768 186320 140820
rect 186372 140808 186378 140820
rect 193214 140808 193220 140820
rect 186372 140780 193220 140808
rect 186372 140768 186378 140780
rect 193214 140768 193220 140780
rect 193272 140768 193278 140820
rect 193324 140752 193352 140848
rect 214374 140836 214380 140848
rect 214432 140836 214438 140888
rect 280890 140836 280896 140888
rect 280948 140876 280954 140888
rect 288618 140876 288624 140888
rect 280948 140848 288624 140876
rect 280948 140836 280954 140848
rect 288618 140836 288624 140848
rect 288676 140836 288682 140888
rect 203426 140768 203432 140820
rect 203484 140808 203490 140820
rect 287698 140808 287704 140820
rect 203484 140780 287704 140808
rect 203484 140768 203490 140780
rect 287698 140768 287704 140780
rect 287756 140768 287762 140820
rect 80422 140700 80428 140752
rect 80480 140740 80486 140752
rect 83458 140740 83464 140752
rect 80480 140712 83464 140740
rect 80480 140700 80486 140712
rect 83458 140700 83464 140712
rect 83516 140700 83522 140752
rect 193306 140700 193312 140752
rect 193364 140700 193370 140752
rect 221458 140700 221464 140752
rect 221516 140740 221522 140752
rect 251910 140740 251916 140752
rect 221516 140712 251916 140740
rect 221516 140700 221522 140712
rect 251910 140700 251916 140712
rect 251968 140700 251974 140752
rect 210050 140496 210056 140548
rect 210108 140536 210114 140548
rect 210108 140508 219434 140536
rect 210108 140496 210114 140508
rect 193030 140428 193036 140480
rect 193088 140468 193094 140480
rect 197354 140468 197360 140480
rect 193088 140440 197360 140468
rect 193088 140428 193094 140440
rect 197354 140428 197360 140440
rect 197412 140428 197418 140480
rect 215386 140468 215392 140480
rect 200086 140440 215392 140468
rect 63126 140088 63132 140140
rect 63184 140128 63190 140140
rect 76006 140128 76012 140140
rect 63184 140100 76012 140128
rect 63184 140088 63190 140100
rect 76006 140088 76012 140100
rect 76064 140088 76070 140140
rect 46842 140020 46848 140072
rect 46900 140060 46906 140072
rect 71406 140060 71412 140072
rect 46900 140032 71412 140060
rect 46900 140020 46906 140032
rect 71406 140020 71412 140032
rect 71464 140020 71470 140072
rect 75822 140020 75828 140072
rect 75880 140060 75886 140072
rect 91922 140060 91928 140072
rect 75880 140032 91928 140060
rect 75880 140020 75886 140032
rect 91922 140020 91928 140032
rect 91980 140020 91986 140072
rect 86862 139408 86868 139460
rect 86920 139448 86926 139460
rect 200086 139448 200114 140440
rect 215386 140428 215392 140440
rect 215444 140428 215450 140480
rect 219406 140060 219434 140508
rect 224586 140428 224592 140480
rect 224644 140468 224650 140480
rect 225690 140468 225696 140480
rect 224644 140440 225696 140468
rect 224644 140428 224650 140440
rect 225690 140428 225696 140440
rect 225748 140428 225754 140480
rect 289078 140060 289084 140072
rect 219406 140032 289084 140060
rect 289078 140020 289084 140032
rect 289136 140020 289142 140072
rect 86920 139420 200114 139448
rect 86920 139408 86926 139420
rect 251174 139408 251180 139460
rect 251232 139448 251238 139460
rect 251910 139448 251916 139460
rect 251232 139420 251916 139448
rect 251232 139408 251238 139420
rect 251910 139408 251916 139420
rect 251968 139408 251974 139460
rect 134610 139340 134616 139392
rect 134668 139380 134674 139392
rect 188522 139380 188528 139392
rect 134668 139352 188528 139380
rect 134668 139340 134674 139352
rect 188522 139340 188528 139352
rect 188580 139340 188586 139392
rect 226334 139340 226340 139392
rect 226392 139380 226398 139392
rect 236086 139380 236092 139392
rect 226392 139352 236092 139380
rect 226392 139340 226398 139352
rect 236086 139340 236092 139352
rect 236144 139340 236150 139392
rect 78030 138728 78036 138780
rect 78088 138768 78094 138780
rect 113818 138768 113824 138780
rect 78088 138740 113824 138768
rect 78088 138728 78094 138740
rect 113818 138728 113824 138740
rect 113876 138728 113882 138780
rect 52086 138660 52092 138712
rect 52144 138700 52150 138712
rect 72326 138700 72332 138712
rect 52144 138672 72332 138700
rect 52144 138660 52150 138672
rect 72326 138660 72332 138672
rect 72384 138660 72390 138712
rect 81894 138660 81900 138712
rect 81952 138700 81958 138712
rect 177298 138700 177304 138712
rect 81952 138672 177304 138700
rect 81952 138660 81958 138672
rect 177298 138660 177304 138672
rect 177356 138660 177362 138712
rect 75914 138048 75920 138100
rect 75972 138088 75978 138100
rect 76374 138088 76380 138100
rect 75972 138060 76380 138088
rect 75972 138048 75978 138060
rect 76374 138048 76380 138060
rect 76432 138048 76438 138100
rect 2866 137912 2872 137964
rect 2924 137952 2930 137964
rect 73062 137952 73068 137964
rect 2924 137924 73068 137952
rect 2924 137912 2930 137924
rect 73062 137912 73068 137924
rect 73120 137912 73126 137964
rect 86126 137912 86132 137964
rect 86184 137952 86190 137964
rect 193306 137952 193312 137964
rect 86184 137924 193312 137952
rect 86184 137912 86190 137924
rect 193306 137912 193312 137924
rect 193364 137912 193370 137964
rect 226702 137912 226708 137964
rect 226760 137952 226766 137964
rect 240134 137952 240140 137964
rect 226760 137924 240140 137952
rect 226760 137912 226766 137924
rect 240134 137912 240140 137924
rect 240192 137952 240198 137964
rect 241422 137952 241428 137964
rect 240192 137924 241428 137952
rect 240192 137912 240198 137924
rect 241422 137912 241428 137924
rect 241480 137912 241486 137964
rect 67174 137300 67180 137352
rect 67232 137340 67238 137352
rect 67542 137340 67548 137352
rect 67232 137312 67548 137340
rect 67232 137300 67238 137312
rect 67542 137300 67548 137312
rect 67600 137300 67606 137352
rect 64782 137232 64788 137284
rect 64840 137272 64846 137284
rect 69198 137272 69204 137284
rect 64840 137244 69204 137272
rect 64840 137232 64846 137244
rect 69198 137232 69204 137244
rect 69256 137232 69262 137284
rect 79594 137232 79600 137284
rect 79652 137272 79658 137284
rect 189074 137272 189080 137284
rect 79652 137244 189080 137272
rect 79652 137232 79658 137244
rect 189074 137232 189080 137244
rect 189132 137232 189138 137284
rect 241422 137232 241428 137284
rect 241480 137272 241486 137284
rect 282178 137272 282184 137284
rect 241480 137244 282184 137272
rect 241480 137232 241486 137244
rect 282178 137232 282184 137244
rect 282236 137232 282242 137284
rect 75546 136688 75552 136740
rect 75604 136728 75610 136740
rect 78766 136728 78772 136740
rect 75604 136700 78772 136728
rect 75604 136688 75610 136700
rect 78766 136688 78772 136700
rect 78824 136688 78830 136740
rect 78490 136620 78496 136672
rect 78548 136660 78554 136672
rect 79318 136660 79324 136672
rect 78548 136632 79324 136660
rect 78548 136620 78554 136632
rect 79318 136620 79324 136632
rect 79376 136620 79382 136672
rect 85482 136620 85488 136672
rect 85540 136660 85546 136672
rect 86218 136660 86224 136672
rect 85540 136632 86224 136660
rect 85540 136620 85546 136632
rect 86218 136620 86224 136632
rect 86276 136620 86282 136672
rect 173802 136552 173808 136604
rect 173860 136592 173866 136604
rect 191742 136592 191748 136604
rect 173860 136564 191748 136592
rect 173860 136552 173866 136564
rect 191742 136552 191748 136564
rect 191800 136552 191806 136604
rect 226702 136280 226708 136332
rect 226760 136320 226766 136332
rect 229830 136320 229836 136332
rect 226760 136292 229836 136320
rect 226760 136280 226766 136292
rect 229830 136280 229836 136292
rect 229888 136280 229894 136332
rect 91738 136144 91744 136196
rect 91796 136184 91802 136196
rect 95970 136184 95976 136196
rect 91796 136156 95976 136184
rect 91796 136144 91802 136156
rect 95970 136144 95976 136156
rect 96028 136144 96034 136196
rect 91002 135872 91008 135924
rect 91060 135912 91066 135924
rect 126606 135912 126612 135924
rect 91060 135884 126612 135912
rect 91060 135872 91066 135884
rect 126606 135872 126612 135884
rect 126664 135872 126670 135924
rect 240042 135872 240048 135924
rect 240100 135912 240106 135924
rect 333974 135912 333980 135924
rect 240100 135884 333980 135912
rect 240100 135872 240106 135884
rect 333974 135872 333980 135884
rect 334032 135872 334038 135924
rect 91186 135532 91192 135584
rect 91244 135572 91250 135584
rect 91830 135572 91836 135584
rect 91244 135544 91836 135572
rect 91244 135532 91250 135544
rect 91830 135532 91836 135544
rect 91888 135532 91894 135584
rect 4798 135260 4804 135312
rect 4856 135300 4862 135312
rect 91186 135300 91192 135312
rect 4856 135272 91192 135300
rect 4856 135260 4862 135272
rect 91186 135260 91192 135272
rect 91244 135260 91250 135312
rect 184198 135260 184204 135312
rect 184256 135300 184262 135312
rect 191742 135300 191748 135312
rect 184256 135272 191748 135300
rect 184256 135260 184262 135272
rect 191742 135260 191748 135272
rect 191800 135260 191806 135312
rect 97442 135192 97448 135244
rect 97500 135232 97506 135244
rect 182910 135232 182916 135244
rect 97500 135204 182916 135232
rect 97500 135192 97506 135204
rect 182910 135192 182916 135204
rect 182968 135192 182974 135244
rect 188982 135192 188988 135244
rect 189040 135232 189046 135244
rect 189718 135232 189724 135244
rect 189040 135204 189724 135232
rect 189040 135192 189046 135204
rect 189718 135192 189724 135204
rect 189776 135192 189782 135244
rect 226334 135192 226340 135244
rect 226392 135232 226398 135244
rect 258718 135232 258724 135244
rect 226392 135204 258724 135232
rect 226392 135192 226398 135204
rect 258718 135192 258724 135204
rect 258776 135192 258782 135244
rect 70302 134988 70308 135040
rect 70360 135028 70366 135040
rect 72418 135028 72424 135040
rect 70360 135000 72424 135028
rect 70360 134988 70366 135000
rect 72418 134988 72424 135000
rect 72476 134988 72482 135040
rect 75914 134620 75920 134632
rect 64846 134592 75920 134620
rect 3418 134512 3424 134564
rect 3476 134552 3482 134564
rect 64846 134552 64874 134592
rect 75914 134580 75920 134592
rect 75972 134580 75978 134632
rect 94406 134580 94412 134632
rect 94464 134620 94470 134632
rect 95142 134620 95148 134632
rect 94464 134592 95148 134620
rect 94464 134580 94470 134592
rect 95142 134580 95148 134592
rect 95200 134580 95206 134632
rect 3476 134524 64874 134552
rect 3476 134512 3482 134524
rect 95142 133968 95148 134020
rect 95200 134008 95206 134020
rect 156782 134008 156788 134020
rect 95200 133980 156788 134008
rect 95200 133968 95206 133980
rect 156782 133968 156788 133980
rect 156840 133968 156846 134020
rect 188890 133968 188896 134020
rect 188948 134008 188954 134020
rect 190454 134008 190460 134020
rect 188948 133980 190460 134008
rect 188948 133968 188954 133980
rect 190454 133968 190460 133980
rect 190512 133968 190518 134020
rect 226702 133900 226708 133952
rect 226760 133940 226766 133952
rect 302878 133940 302884 133952
rect 226760 133912 302884 133940
rect 226760 133900 226766 133912
rect 302878 133900 302884 133912
rect 302936 133900 302942 133952
rect 64598 133832 64604 133884
rect 64656 133872 64662 133884
rect 66806 133872 66812 133884
rect 64656 133844 66812 133872
rect 64656 133832 64662 133844
rect 66806 133832 66812 133844
rect 66864 133832 66870 133884
rect 96706 133832 96712 133884
rect 96764 133872 96770 133884
rect 114002 133872 114008 133884
rect 96764 133844 114008 133872
rect 96764 133832 96770 133844
rect 114002 133832 114008 133844
rect 114060 133832 114066 133884
rect 165062 133832 165068 133884
rect 165120 133872 165126 133884
rect 186314 133872 186320 133884
rect 165120 133844 186320 133872
rect 165120 133832 165126 133844
rect 186314 133832 186320 133844
rect 186372 133832 186378 133884
rect 226334 133832 226340 133884
rect 226392 133872 226398 133884
rect 269114 133872 269120 133884
rect 226392 133844 269120 133872
rect 226392 133832 226398 133844
rect 269114 133832 269120 133844
rect 269172 133832 269178 133884
rect 226702 133764 226708 133816
rect 226760 133804 226766 133816
rect 233878 133804 233884 133816
rect 226760 133776 233884 133804
rect 226760 133764 226766 133776
rect 233878 133764 233884 133776
rect 233936 133764 233942 133816
rect 226426 133492 226432 133544
rect 226484 133532 226490 133544
rect 226702 133532 226708 133544
rect 226484 133504 226708 133532
rect 226484 133492 226490 133504
rect 226702 133492 226708 133504
rect 226760 133492 226766 133544
rect 113818 133152 113824 133204
rect 113876 133192 113882 133204
rect 126422 133192 126428 133204
rect 113876 133164 126428 133192
rect 113876 133152 113882 133164
rect 126422 133152 126428 133164
rect 126480 133152 126486 133204
rect 134610 133152 134616 133204
rect 134668 133192 134674 133204
rect 148502 133192 148508 133204
rect 134668 133164 148508 133192
rect 134668 133152 134674 133164
rect 148502 133152 148508 133164
rect 148560 133152 148566 133204
rect 148686 133152 148692 133204
rect 148744 133192 148750 133204
rect 184382 133192 184388 133204
rect 148744 133164 184388 133192
rect 148744 133152 148750 133164
rect 184382 133152 184388 133164
rect 184440 133152 184446 133204
rect 50982 132404 50988 132456
rect 51040 132444 51046 132456
rect 66806 132444 66812 132456
rect 51040 132416 66812 132444
rect 51040 132404 51046 132416
rect 66806 132404 66812 132416
rect 66864 132404 66870 132456
rect 105630 132404 105636 132456
rect 105688 132444 105694 132456
rect 105688 132416 180794 132444
rect 105688 132404 105694 132416
rect 57698 132336 57704 132388
rect 57756 132376 57762 132388
rect 66254 132376 66260 132388
rect 57756 132348 66260 132376
rect 57756 132336 57762 132348
rect 66254 132336 66260 132348
rect 66312 132336 66318 132388
rect 96706 132336 96712 132388
rect 96764 132376 96770 132388
rect 148594 132376 148600 132388
rect 96764 132348 148600 132376
rect 96764 132336 96770 132348
rect 148594 132336 148600 132348
rect 148652 132336 148658 132388
rect 180766 132376 180794 132416
rect 188338 132404 188344 132456
rect 188396 132444 188402 132456
rect 191650 132444 191656 132456
rect 188396 132416 191656 132444
rect 188396 132404 188402 132416
rect 191650 132404 191656 132416
rect 191708 132404 191714 132456
rect 226334 132404 226340 132456
rect 226392 132444 226398 132456
rect 231946 132444 231952 132456
rect 226392 132416 231952 132444
rect 226392 132404 226398 132416
rect 231946 132404 231952 132416
rect 232004 132404 232010 132456
rect 191098 132376 191104 132388
rect 180766 132348 191104 132376
rect 191098 132336 191104 132348
rect 191156 132336 191162 132388
rect 41322 131724 41328 131776
rect 41380 131764 41386 131776
rect 48314 131764 48320 131776
rect 41380 131736 48320 131764
rect 41380 131724 41386 131736
rect 48314 131724 48320 131736
rect 48372 131724 48378 131776
rect 231210 131724 231216 131776
rect 231268 131764 231274 131776
rect 276014 131764 276020 131776
rect 231268 131736 276020 131764
rect 231268 131724 231274 131736
rect 276014 131724 276020 131736
rect 276072 131724 276078 131776
rect 148410 131112 148416 131164
rect 148468 131152 148474 131164
rect 153838 131152 153844 131164
rect 148468 131124 153844 131152
rect 148468 131112 148474 131124
rect 153838 131112 153844 131124
rect 153896 131112 153902 131164
rect 176010 131044 176016 131096
rect 176068 131084 176074 131096
rect 189994 131084 190000 131096
rect 176068 131056 190000 131084
rect 176068 131044 176074 131056
rect 189994 131044 190000 131056
rect 190052 131044 190058 131096
rect 226702 131044 226708 131096
rect 226760 131084 226766 131096
rect 230474 131084 230480 131096
rect 226760 131056 230480 131084
rect 226760 131044 226766 131056
rect 230474 131044 230480 131056
rect 230532 131084 230538 131096
rect 273254 131084 273260 131096
rect 230532 131056 273260 131084
rect 230532 131044 230538 131056
rect 273254 131044 273260 131056
rect 273312 131044 273318 131096
rect 226794 130976 226800 131028
rect 226852 131016 226858 131028
rect 240318 131016 240324 131028
rect 226852 130988 240324 131016
rect 226852 130976 226858 130988
rect 240318 130976 240324 130988
rect 240376 130976 240382 131028
rect 96798 130364 96804 130416
rect 96856 130404 96862 130416
rect 170490 130404 170496 130416
rect 96856 130376 170496 130404
rect 96856 130364 96862 130376
rect 170490 130364 170496 130376
rect 170548 130364 170554 130416
rect 176010 130364 176016 130416
rect 176068 130404 176074 130416
rect 176562 130404 176568 130416
rect 176068 130376 176568 130404
rect 176068 130364 176074 130376
rect 176562 130364 176568 130376
rect 176620 130364 176626 130416
rect 96706 130160 96712 130212
rect 96764 130200 96770 130212
rect 102962 130200 102968 130212
rect 96764 130172 102968 130200
rect 96764 130160 96770 130172
rect 102962 130160 102968 130172
rect 103020 130160 103026 130212
rect 94774 129684 94780 129736
rect 94832 129724 94838 129736
rect 95878 129724 95884 129736
rect 94832 129696 95884 129724
rect 94832 129684 94838 129696
rect 95878 129684 95884 129696
rect 95936 129684 95942 129736
rect 187510 129724 187516 129736
rect 99346 129696 187516 129724
rect 94958 129616 94964 129668
rect 95016 129656 95022 129668
rect 99346 129656 99374 129696
rect 187510 129684 187516 129696
rect 187568 129724 187574 129736
rect 191742 129724 191748 129736
rect 187568 129696 191748 129724
rect 187568 129684 187574 129696
rect 191742 129684 191748 129696
rect 191800 129684 191806 129736
rect 229738 129684 229744 129736
rect 229796 129724 229802 129736
rect 259454 129724 259460 129736
rect 229796 129696 259460 129724
rect 229796 129684 229802 129696
rect 259454 129684 259460 129696
rect 259512 129684 259518 129736
rect 95016 129628 99374 129656
rect 95016 129616 95022 129628
rect 226518 129004 226524 129056
rect 226576 129044 226582 129056
rect 226702 129044 226708 129056
rect 226576 129016 226708 129044
rect 226576 129004 226582 129016
rect 226702 129004 226708 129016
rect 226760 129044 226766 129056
rect 299474 129044 299480 129056
rect 226760 129016 299480 129044
rect 226760 129004 226766 129016
rect 299474 129004 299480 129016
rect 299532 129004 299538 129056
rect 63218 128256 63224 128308
rect 63276 128296 63282 128308
rect 66806 128296 66812 128308
rect 63276 128268 66812 128296
rect 63276 128256 63282 128268
rect 66806 128256 66812 128268
rect 66864 128256 66870 128308
rect 97626 128256 97632 128308
rect 97684 128296 97690 128308
rect 142982 128296 142988 128308
rect 97684 128268 142988 128296
rect 97684 128256 97690 128268
rect 142982 128256 142988 128268
rect 143040 128256 143046 128308
rect 226702 127644 226708 127696
rect 226760 127684 226766 127696
rect 226886 127684 226892 127696
rect 226760 127656 226892 127684
rect 226760 127644 226766 127656
rect 226886 127644 226892 127656
rect 226944 127684 226950 127696
rect 260098 127684 260104 127696
rect 226944 127656 260104 127684
rect 226944 127644 226950 127656
rect 260098 127644 260104 127656
rect 260156 127644 260162 127696
rect 126330 127576 126336 127628
rect 126388 127616 126394 127628
rect 135990 127616 135996 127628
rect 126388 127588 135996 127616
rect 126388 127576 126394 127588
rect 135990 127576 135996 127588
rect 136048 127576 136054 127628
rect 227990 127576 227996 127628
rect 228048 127616 228054 127628
rect 267918 127616 267924 127628
rect 228048 127588 267924 127616
rect 228048 127576 228054 127588
rect 267918 127576 267924 127588
rect 267976 127576 267982 127628
rect 268378 127576 268384 127628
rect 268436 127616 268442 127628
rect 295334 127616 295340 127628
rect 268436 127588 295340 127616
rect 268436 127576 268442 127588
rect 295334 127576 295340 127588
rect 295392 127576 295398 127628
rect 192294 127004 192300 127016
rect 158732 126976 192300 127004
rect 97258 126896 97264 126948
rect 97316 126936 97322 126948
rect 111242 126936 111248 126948
rect 97316 126908 111248 126936
rect 97316 126896 97322 126908
rect 111242 126896 111248 126908
rect 111300 126896 111306 126948
rect 158070 126896 158076 126948
rect 158128 126936 158134 126948
rect 158732 126936 158760 126976
rect 192294 126964 192300 126976
rect 192352 127004 192358 127016
rect 192846 127004 192852 127016
rect 192352 126976 192852 127004
rect 192352 126964 192358 126976
rect 192846 126964 192852 126976
rect 192904 126964 192910 127016
rect 158128 126908 158760 126936
rect 158128 126896 158134 126908
rect 226334 126896 226340 126948
rect 226392 126936 226398 126948
rect 242894 126936 242900 126948
rect 226392 126908 242900 126936
rect 226392 126896 226398 126908
rect 242894 126896 242900 126908
rect 242952 126936 242958 126948
rect 243354 126936 243360 126948
rect 242952 126908 243360 126936
rect 242952 126896 242958 126908
rect 243354 126896 243360 126908
rect 243412 126896 243418 126948
rect 295334 126896 295340 126948
rect 295392 126936 295398 126948
rect 302326 126936 302332 126948
rect 295392 126908 302332 126936
rect 295392 126896 295398 126908
rect 302326 126896 302332 126908
rect 302384 126896 302390 126948
rect 182818 126828 182824 126880
rect 182876 126868 182882 126880
rect 192386 126868 192392 126880
rect 182876 126840 192392 126868
rect 182876 126828 182882 126840
rect 192386 126828 192392 126840
rect 192444 126828 192450 126880
rect 108482 126216 108488 126268
rect 108540 126256 108546 126268
rect 187510 126256 187516 126268
rect 108540 126228 187516 126256
rect 108540 126216 108546 126228
rect 187510 126216 187516 126228
rect 187568 126216 187574 126268
rect 243354 126216 243360 126268
rect 243412 126256 243418 126268
rect 351914 126256 351920 126268
rect 243412 126228 351920 126256
rect 243412 126216 243418 126228
rect 351914 126216 351920 126228
rect 351972 126216 351978 126268
rect 187510 125672 187516 125724
rect 187568 125712 187574 125724
rect 190362 125712 190368 125724
rect 187568 125684 190368 125712
rect 187568 125672 187574 125684
rect 190362 125672 190368 125684
rect 190420 125672 190426 125724
rect 52178 125536 52184 125588
rect 52236 125576 52242 125588
rect 66898 125576 66904 125588
rect 52236 125548 66904 125576
rect 52236 125536 52242 125548
rect 66898 125536 66904 125548
rect 66956 125536 66962 125588
rect 97534 125536 97540 125588
rect 97592 125576 97598 125588
rect 148686 125576 148692 125588
rect 97592 125548 148692 125576
rect 97592 125536 97598 125548
rect 148686 125536 148692 125548
rect 148744 125536 148750 125588
rect 167730 125536 167736 125588
rect 167788 125576 167794 125588
rect 190270 125576 190276 125588
rect 167788 125548 190276 125576
rect 167788 125536 167794 125548
rect 190270 125536 190276 125548
rect 190328 125536 190334 125588
rect 56502 124856 56508 124908
rect 56560 124896 56566 124908
rect 66806 124896 66812 124908
rect 56560 124868 66812 124896
rect 56560 124856 56566 124868
rect 66806 124856 66812 124868
rect 66864 124856 66870 124908
rect 96614 124856 96620 124908
rect 96672 124896 96678 124908
rect 175918 124896 175924 124908
rect 96672 124868 175924 124896
rect 96672 124856 96678 124868
rect 175918 124856 175924 124868
rect 175976 124856 175982 124908
rect 232498 124856 232504 124908
rect 232556 124896 232562 124908
rect 295426 124896 295432 124908
rect 232556 124868 295432 124896
rect 232556 124856 232562 124868
rect 295426 124856 295432 124868
rect 295484 124856 295490 124908
rect 188798 124788 188804 124840
rect 188856 124828 188862 124840
rect 192938 124828 192944 124840
rect 188856 124800 192944 124828
rect 188856 124788 188862 124800
rect 192938 124788 192944 124800
rect 192996 124788 193002 124840
rect 226518 124720 226524 124772
rect 226576 124760 226582 124772
rect 229738 124760 229744 124772
rect 226576 124732 229744 124760
rect 226576 124720 226582 124732
rect 229738 124720 229744 124732
rect 229796 124720 229802 124772
rect 61930 124108 61936 124160
rect 61988 124148 61994 124160
rect 66254 124148 66260 124160
rect 61988 124120 66260 124148
rect 61988 124108 61994 124120
rect 66254 124108 66260 124120
rect 66312 124108 66318 124160
rect 97902 124108 97908 124160
rect 97960 124148 97966 124160
rect 152642 124148 152648 124160
rect 97960 124120 152648 124148
rect 97960 124108 97966 124120
rect 152642 124108 152648 124120
rect 152700 124108 152706 124160
rect 226334 124108 226340 124160
rect 226392 124148 226398 124160
rect 229094 124148 229100 124160
rect 226392 124120 229100 124148
rect 226392 124108 226398 124120
rect 229094 124108 229100 124120
rect 229152 124148 229158 124160
rect 280798 124148 280804 124160
rect 229152 124120 280804 124148
rect 229152 124108 229158 124120
rect 280798 124108 280804 124120
rect 280856 124148 280862 124160
rect 582834 124148 582840 124160
rect 280856 124120 582840 124148
rect 280856 124108 280862 124120
rect 582834 124108 582840 124120
rect 582892 124108 582898 124160
rect 228358 123428 228364 123480
rect 228416 123468 228422 123480
rect 255958 123468 255964 123480
rect 228416 123440 255964 123468
rect 228416 123428 228422 123440
rect 255958 123428 255964 123440
rect 256016 123428 256022 123480
rect 191742 122856 191748 122868
rect 188264 122828 191748 122856
rect 59078 122748 59084 122800
rect 59136 122788 59142 122800
rect 66346 122788 66352 122800
rect 59136 122760 66352 122788
rect 59136 122748 59142 122760
rect 66346 122748 66352 122760
rect 66404 122748 66410 122800
rect 97534 122748 97540 122800
rect 97592 122788 97598 122800
rect 119338 122788 119344 122800
rect 97592 122760 119344 122788
rect 97592 122748 97598 122760
rect 119338 122748 119344 122760
rect 119396 122748 119402 122800
rect 155862 122748 155868 122800
rect 155920 122788 155926 122800
rect 188264 122788 188292 122828
rect 191742 122816 191748 122828
rect 191800 122816 191806 122868
rect 155920 122760 188292 122788
rect 155920 122748 155926 122760
rect 226334 122748 226340 122800
rect 226392 122788 226398 122800
rect 247034 122788 247040 122800
rect 226392 122760 247040 122788
rect 226392 122748 226398 122760
rect 247034 122748 247040 122760
rect 247092 122748 247098 122800
rect 189810 122340 189816 122392
rect 189868 122380 189874 122392
rect 190362 122380 190368 122392
rect 189868 122352 190368 122380
rect 189868 122340 189874 122352
rect 190362 122340 190368 122352
rect 190420 122340 190426 122392
rect 112438 122068 112444 122120
rect 112496 122108 112502 122120
rect 188338 122108 188344 122120
rect 112496 122080 188344 122108
rect 112496 122068 112502 122080
rect 188338 122068 188344 122080
rect 188396 122068 188402 122120
rect 225690 122068 225696 122120
rect 225748 122108 225754 122120
rect 313274 122108 313280 122120
rect 225748 122080 313280 122108
rect 225748 122068 225754 122080
rect 313274 122068 313280 122080
rect 313332 122068 313338 122120
rect 61838 121388 61844 121440
rect 61896 121428 61902 121440
rect 66806 121428 66812 121440
rect 61896 121400 66812 121428
rect 61896 121388 61902 121400
rect 66806 121388 66812 121400
rect 66864 121388 66870 121440
rect 97718 121388 97724 121440
rect 97776 121428 97782 121440
rect 151170 121428 151176 121440
rect 97776 121400 151176 121428
rect 97776 121388 97782 121400
rect 151170 121388 151176 121400
rect 151228 121388 151234 121440
rect 159542 121388 159548 121440
rect 159600 121428 159606 121440
rect 191190 121428 191196 121440
rect 159600 121400 191196 121428
rect 159600 121388 159606 121400
rect 191190 121388 191196 121400
rect 191248 121388 191254 121440
rect 226426 121388 226432 121440
rect 226484 121428 226490 121440
rect 244366 121428 244372 121440
rect 226484 121400 244372 121428
rect 226484 121388 226490 121400
rect 244366 121388 244372 121400
rect 244424 121388 244430 121440
rect 240870 120708 240876 120760
rect 240928 120748 240934 120760
rect 274634 120748 274640 120760
rect 240928 120720 274640 120748
rect 240928 120708 240934 120720
rect 274634 120708 274640 120720
rect 274692 120708 274698 120760
rect 184750 120640 184756 120692
rect 184808 120680 184814 120692
rect 191742 120680 191748 120692
rect 184808 120652 191748 120680
rect 184808 120640 184814 120652
rect 191742 120640 191748 120652
rect 191800 120640 191806 120692
rect 97534 120096 97540 120148
rect 97592 120136 97598 120148
rect 105538 120136 105544 120148
rect 97592 120108 105544 120136
rect 97592 120096 97598 120108
rect 105538 120096 105544 120108
rect 105596 120096 105602 120148
rect 49510 120028 49516 120080
rect 49568 120068 49574 120080
rect 66806 120068 66812 120080
rect 49568 120040 66812 120068
rect 49568 120028 49574 120040
rect 66806 120028 66812 120040
rect 66864 120028 66870 120080
rect 97718 120028 97724 120080
rect 97776 120068 97782 120080
rect 122098 120068 122104 120080
rect 97776 120040 122104 120068
rect 97776 120028 97782 120040
rect 122098 120028 122104 120040
rect 122156 120028 122162 120080
rect 184290 120028 184296 120080
rect 184348 120068 184354 120080
rect 191742 120068 191748 120080
rect 184348 120040 191748 120068
rect 184348 120028 184354 120040
rect 191742 120028 191748 120040
rect 191800 120028 191806 120080
rect 284938 119348 284944 119400
rect 284996 119388 285002 119400
rect 289906 119388 289912 119400
rect 284996 119360 289912 119388
rect 284996 119348 285002 119360
rect 289906 119348 289912 119360
rect 289964 119348 289970 119400
rect 57790 118600 57796 118652
rect 57848 118640 57854 118652
rect 66898 118640 66904 118652
rect 57848 118612 66904 118640
rect 57848 118600 57854 118612
rect 66898 118600 66904 118612
rect 66956 118600 66962 118652
rect 97902 118600 97908 118652
rect 97960 118640 97966 118652
rect 133230 118640 133236 118652
rect 97960 118612 133236 118640
rect 97960 118600 97966 118612
rect 133230 118600 133236 118612
rect 133288 118600 133294 118652
rect 64506 118532 64512 118584
rect 64564 118572 64570 118584
rect 66806 118572 66812 118584
rect 64564 118544 66812 118572
rect 64564 118532 64570 118544
rect 66806 118532 66812 118544
rect 66864 118532 66870 118584
rect 97810 117920 97816 117972
rect 97868 117960 97874 117972
rect 100018 117960 100024 117972
rect 97868 117932 100024 117960
rect 97868 117920 97874 117932
rect 100018 117920 100024 117932
rect 100076 117960 100082 117972
rect 173250 117960 173256 117972
rect 100076 117932 173256 117960
rect 100076 117920 100082 117932
rect 173250 117920 173256 117932
rect 173308 117920 173314 117972
rect 180150 117920 180156 117972
rect 180208 117960 180214 117972
rect 187694 117960 187700 117972
rect 180208 117932 187700 117960
rect 180208 117920 180214 117932
rect 187694 117920 187700 117932
rect 187752 117920 187758 117972
rect 187694 117376 187700 117428
rect 187752 117416 187758 117428
rect 188982 117416 188988 117428
rect 187752 117388 188988 117416
rect 187752 117376 187758 117388
rect 188982 117376 188988 117388
rect 189040 117416 189046 117428
rect 191742 117416 191748 117428
rect 189040 117388 191748 117416
rect 189040 117376 189046 117388
rect 191742 117376 191748 117388
rect 191800 117376 191806 117428
rect 226518 117376 226524 117428
rect 226576 117416 226582 117428
rect 233878 117416 233884 117428
rect 226576 117388 233884 117416
rect 226576 117376 226582 117388
rect 233878 117376 233884 117388
rect 233936 117376 233942 117428
rect 226702 117308 226708 117360
rect 226760 117348 226766 117360
rect 244274 117348 244280 117360
rect 226760 117320 244280 117348
rect 226760 117308 226766 117320
rect 244274 117308 244280 117320
rect 244332 117308 244338 117360
rect 97350 117240 97356 117292
rect 97408 117280 97414 117292
rect 145650 117280 145656 117292
rect 97408 117252 145656 117280
rect 97408 117240 97414 117252
rect 145650 117240 145656 117252
rect 145708 117240 145714 117292
rect 185670 117240 185676 117292
rect 185728 117280 185734 117292
rect 191742 117280 191748 117292
rect 185728 117252 191748 117280
rect 185728 117240 185734 117252
rect 191742 117240 191748 117252
rect 191800 117240 191806 117292
rect 54938 117172 54944 117224
rect 54996 117212 55002 117224
rect 66806 117212 66812 117224
rect 54996 117184 66812 117212
rect 54996 117172 55002 117184
rect 66806 117172 66812 117184
rect 66864 117172 66870 117224
rect 97902 117172 97908 117224
rect 97960 117212 97966 117224
rect 136082 117212 136088 117224
rect 97960 117184 136088 117212
rect 97960 117172 97966 117184
rect 136082 117172 136088 117184
rect 136140 117172 136146 117224
rect 231762 116560 231768 116612
rect 231820 116600 231826 116612
rect 262398 116600 262404 116612
rect 231820 116572 262404 116600
rect 231820 116560 231826 116572
rect 262398 116560 262404 116572
rect 262456 116560 262462 116612
rect 291654 116560 291660 116612
rect 291712 116600 291718 116612
rect 304258 116600 304264 116612
rect 291712 116572 304264 116600
rect 291712 116560 291718 116572
rect 304258 116560 304264 116572
rect 304316 116560 304322 116612
rect 185762 116016 185768 116068
rect 185820 116056 185826 116068
rect 191282 116056 191288 116068
rect 185820 116028 191288 116056
rect 185820 116016 185826 116028
rect 191282 116016 191288 116028
rect 191340 116016 191346 116068
rect 226702 115948 226708 116000
rect 226760 115988 226766 116000
rect 230474 115988 230480 116000
rect 226760 115960 230480 115988
rect 226760 115948 226766 115960
rect 230474 115948 230480 115960
rect 230532 115988 230538 116000
rect 231762 115988 231768 116000
rect 230532 115960 231768 115988
rect 230532 115948 230538 115960
rect 231762 115948 231768 115960
rect 231820 115948 231826 116000
rect 57882 115880 57888 115932
rect 57940 115920 57946 115932
rect 66806 115920 66812 115932
rect 57940 115892 66812 115920
rect 57940 115880 57946 115892
rect 66806 115880 66812 115892
rect 66864 115880 66870 115932
rect 175182 115880 175188 115932
rect 175240 115920 175246 115932
rect 191006 115920 191012 115932
rect 175240 115892 191012 115920
rect 175240 115880 175246 115892
rect 191006 115880 191012 115892
rect 191064 115880 191070 115932
rect 63310 115268 63316 115320
rect 63368 115308 63374 115320
rect 66806 115308 66812 115320
rect 63368 115280 66812 115308
rect 63368 115268 63374 115280
rect 66806 115268 66812 115280
rect 66864 115268 66870 115320
rect 233326 115200 233332 115252
rect 233384 115240 233390 115252
rect 280154 115240 280160 115252
rect 233384 115212 280160 115240
rect 233384 115200 233390 115212
rect 280154 115200 280160 115212
rect 280212 115200 280218 115252
rect 97534 114588 97540 114640
rect 97592 114628 97598 114640
rect 112438 114628 112444 114640
rect 97592 114600 112444 114628
rect 97592 114588 97598 114600
rect 112438 114588 112444 114600
rect 112496 114588 112502 114640
rect 97902 114520 97908 114572
rect 97960 114560 97966 114572
rect 170490 114560 170496 114572
rect 97960 114532 170496 114560
rect 97960 114520 97966 114532
rect 170490 114520 170496 114532
rect 170548 114520 170554 114572
rect 226334 114520 226340 114572
rect 226392 114560 226398 114572
rect 233326 114560 233332 114572
rect 226392 114532 233332 114560
rect 226392 114520 226398 114532
rect 233326 114520 233332 114532
rect 233384 114520 233390 114572
rect 58986 114452 58992 114504
rect 59044 114492 59050 114504
rect 66806 114492 66812 114504
rect 59044 114464 66812 114492
rect 59044 114452 59050 114464
rect 66806 114452 66812 114464
rect 66864 114452 66870 114504
rect 7558 113772 7564 113824
rect 7616 113812 7622 113824
rect 65978 113812 65984 113824
rect 7616 113784 65984 113812
rect 7616 113772 7622 113784
rect 65978 113772 65984 113784
rect 66036 113772 66042 113824
rect 96706 113772 96712 113824
rect 96764 113812 96770 113824
rect 134794 113812 134800 113824
rect 96764 113784 134800 113812
rect 96764 113772 96770 113784
rect 134794 113772 134800 113784
rect 134852 113772 134858 113824
rect 160922 113772 160928 113824
rect 160980 113812 160986 113824
rect 183370 113812 183376 113824
rect 160980 113784 183376 113812
rect 160980 113772 160986 113784
rect 183370 113772 183376 113784
rect 183428 113772 183434 113824
rect 188246 113228 188252 113280
rect 188304 113268 188310 113280
rect 191190 113268 191196 113280
rect 188304 113240 191196 113268
rect 188304 113228 188310 113240
rect 191190 113228 191196 113240
rect 191248 113228 191254 113280
rect 183370 113160 183376 113212
rect 183428 113200 183434 113212
rect 191742 113200 191748 113212
rect 183428 113172 191748 113200
rect 183428 113160 183434 113172
rect 191742 113160 191748 113172
rect 191800 113160 191806 113212
rect 63126 113092 63132 113144
rect 63184 113132 63190 113144
rect 66806 113132 66812 113144
rect 63184 113104 66812 113132
rect 63184 113092 63190 113104
rect 66806 113092 66812 113104
rect 66864 113092 66870 113144
rect 226702 113092 226708 113144
rect 226760 113132 226766 113144
rect 233234 113132 233240 113144
rect 226760 113104 233240 113132
rect 226760 113092 226766 113104
rect 233234 113092 233240 113104
rect 233292 113092 233298 113144
rect 60550 113024 60556 113076
rect 60608 113064 60614 113076
rect 66898 113064 66904 113076
rect 60608 113036 66904 113064
rect 60608 113024 60614 113036
rect 66898 113024 66904 113036
rect 66956 113024 66962 113076
rect 225598 112480 225604 112532
rect 225656 112520 225662 112532
rect 253014 112520 253020 112532
rect 225656 112492 253020 112520
rect 225656 112480 225662 112492
rect 253014 112480 253020 112492
rect 253072 112480 253078 112532
rect 104250 112412 104256 112464
rect 104308 112452 104314 112464
rect 191558 112452 191564 112464
rect 104308 112424 191564 112452
rect 104308 112412 104314 112424
rect 191558 112412 191564 112424
rect 191616 112412 191622 112464
rect 233234 112412 233240 112464
rect 233292 112452 233298 112464
rect 324406 112452 324412 112464
rect 233292 112424 324412 112452
rect 233292 112412 233298 112424
rect 324406 112412 324412 112424
rect 324464 112412 324470 112464
rect 98086 111936 98092 111988
rect 98144 111976 98150 111988
rect 101582 111976 101588 111988
rect 98144 111948 101588 111976
rect 98144 111936 98150 111948
rect 101582 111936 101588 111948
rect 101640 111936 101646 111988
rect 96890 111868 96896 111920
rect 96948 111908 96954 111920
rect 98638 111908 98644 111920
rect 96948 111880 98644 111908
rect 96948 111868 96954 111880
rect 98638 111868 98644 111880
rect 98696 111868 98702 111920
rect 97902 111800 97908 111852
rect 97960 111840 97966 111852
rect 160738 111840 160744 111852
rect 97960 111812 160744 111840
rect 97960 111800 97966 111812
rect 160738 111800 160744 111812
rect 160796 111800 160802 111852
rect 55122 111732 55128 111784
rect 55180 111772 55186 111784
rect 66806 111772 66812 111784
rect 55180 111744 66812 111772
rect 55180 111732 55186 111744
rect 66806 111732 66812 111744
rect 66864 111732 66870 111784
rect 97350 111732 97356 111784
rect 97408 111772 97414 111784
rect 113910 111772 113916 111784
rect 97408 111744 113916 111772
rect 97408 111732 97414 111744
rect 113910 111732 113916 111744
rect 113968 111732 113974 111784
rect 153930 111732 153936 111784
rect 153988 111772 153994 111784
rect 191374 111772 191380 111784
rect 153988 111744 191380 111772
rect 153988 111732 153994 111744
rect 191374 111732 191380 111744
rect 191432 111732 191438 111784
rect 252646 111732 252652 111784
rect 252704 111772 252710 111784
rect 253014 111772 253020 111784
rect 252704 111744 253020 111772
rect 252704 111732 252710 111744
rect 253014 111732 253020 111744
rect 253072 111772 253078 111784
rect 260190 111772 260196 111784
rect 253072 111744 260196 111772
rect 253072 111732 253078 111744
rect 260190 111732 260196 111744
rect 260248 111732 260254 111784
rect 226334 111120 226340 111172
rect 226392 111160 226398 111172
rect 229094 111160 229100 111172
rect 226392 111132 229100 111160
rect 226392 111120 226398 111132
rect 229094 111120 229100 111132
rect 229152 111160 229158 111172
rect 235994 111160 236000 111172
rect 229152 111132 236000 111160
rect 229152 111120 229158 111132
rect 235994 111120 236000 111132
rect 236052 111120 236058 111172
rect 159358 111052 159364 111104
rect 159416 111092 159422 111104
rect 185762 111092 185768 111104
rect 159416 111064 185768 111092
rect 159416 111052 159422 111064
rect 185762 111052 185768 111064
rect 185820 111052 185826 111104
rect 226518 111052 226524 111104
rect 226576 111092 226582 111104
rect 291194 111092 291200 111104
rect 226576 111064 291200 111092
rect 226576 111052 226582 111064
rect 291194 111052 291200 111064
rect 291252 111052 291258 111104
rect 2866 110780 2872 110832
rect 2924 110820 2930 110832
rect 4798 110820 4804 110832
rect 2924 110792 4804 110820
rect 2924 110780 2930 110792
rect 4798 110780 4804 110792
rect 4856 110780 4862 110832
rect 291194 110440 291200 110492
rect 291252 110480 291258 110492
rect 291838 110480 291844 110492
rect 291252 110452 291844 110480
rect 291252 110440 291258 110452
rect 291838 110440 291844 110452
rect 291896 110440 291902 110492
rect 59262 110372 59268 110424
rect 59320 110412 59326 110424
rect 66806 110412 66812 110424
rect 59320 110384 66812 110412
rect 59320 110372 59326 110384
rect 66806 110372 66812 110384
rect 66864 110372 66870 110424
rect 226978 109760 226984 109812
rect 227036 109800 227042 109812
rect 267826 109800 267832 109812
rect 227036 109772 267832 109800
rect 227036 109760 227042 109772
rect 267826 109760 267832 109772
rect 267884 109760 267890 109812
rect 104250 109692 104256 109744
rect 104308 109732 104314 109744
rect 149790 109732 149796 109744
rect 104308 109704 149796 109732
rect 104308 109692 104314 109704
rect 149790 109692 149796 109704
rect 149848 109692 149854 109744
rect 153838 109692 153844 109744
rect 153896 109732 153902 109744
rect 188246 109732 188252 109744
rect 153896 109704 188252 109732
rect 153896 109692 153902 109704
rect 188246 109692 188252 109704
rect 188304 109692 188310 109744
rect 225598 109692 225604 109744
rect 225656 109732 225662 109744
rect 252554 109732 252560 109744
rect 225656 109704 252560 109732
rect 225656 109692 225662 109704
rect 252554 109692 252560 109704
rect 252612 109732 252618 109744
rect 345658 109732 345664 109744
rect 252612 109704 345664 109732
rect 252612 109692 252618 109704
rect 345658 109692 345664 109704
rect 345716 109692 345722 109744
rect 48222 109012 48228 109064
rect 48280 109052 48286 109064
rect 52546 109052 52552 109064
rect 48280 109024 52552 109052
rect 48280 109012 48286 109024
rect 52546 109012 52552 109024
rect 52604 109052 52610 109064
rect 66898 109052 66904 109064
rect 52604 109024 66904 109052
rect 52604 109012 52610 109024
rect 66898 109012 66904 109024
rect 66956 109012 66962 109064
rect 53650 108944 53656 108996
rect 53708 108984 53714 108996
rect 66714 108984 66720 108996
rect 53708 108956 66720 108984
rect 53708 108944 53714 108956
rect 66714 108944 66720 108956
rect 66772 108944 66778 108996
rect 97902 108944 97908 108996
rect 97960 108984 97966 108996
rect 114646 108984 114652 108996
rect 97960 108956 114652 108984
rect 97960 108944 97966 108956
rect 114646 108944 114652 108956
rect 114704 108984 114710 108996
rect 115842 108984 115848 108996
rect 114704 108956 115848 108984
rect 114704 108944 114710 108956
rect 115842 108944 115848 108956
rect 115900 108944 115906 108996
rect 166442 108944 166448 108996
rect 166500 108984 166506 108996
rect 190270 108984 190276 108996
rect 166500 108956 190276 108984
rect 166500 108944 166506 108956
rect 190270 108944 190276 108956
rect 190328 108944 190334 108996
rect 226518 108944 226524 108996
rect 226576 108984 226582 108996
rect 245654 108984 245660 108996
rect 226576 108956 245660 108984
rect 226576 108944 226582 108956
rect 245654 108944 245660 108956
rect 245712 108944 245718 108996
rect 64782 108876 64788 108928
rect 64840 108916 64846 108928
rect 66438 108916 66444 108928
rect 64840 108888 66444 108916
rect 64840 108876 64846 108888
rect 66438 108876 66444 108888
rect 66496 108876 66502 108928
rect 183462 108876 183468 108928
rect 183520 108916 183526 108928
rect 191190 108916 191196 108928
rect 183520 108888 191196 108916
rect 183520 108876 183526 108888
rect 191190 108876 191196 108888
rect 191248 108876 191254 108928
rect 104894 108332 104900 108384
rect 104952 108372 104958 108384
rect 144178 108372 144184 108384
rect 104952 108344 144184 108372
rect 104952 108332 104958 108344
rect 144178 108332 144184 108344
rect 144236 108332 144242 108384
rect 115842 108264 115848 108316
rect 115900 108304 115906 108316
rect 180150 108304 180156 108316
rect 115900 108276 180156 108304
rect 115900 108264 115906 108276
rect 180150 108264 180156 108276
rect 180208 108264 180214 108316
rect 227070 108264 227076 108316
rect 227128 108304 227134 108316
rect 227714 108304 227720 108316
rect 227128 108276 227720 108304
rect 227128 108264 227134 108276
rect 227714 108264 227720 108276
rect 227772 108304 227778 108316
rect 270586 108304 270592 108316
rect 227772 108276 270592 108304
rect 227772 108264 227778 108276
rect 270586 108264 270592 108276
rect 270644 108264 270650 108316
rect 189074 107720 189080 107772
rect 189132 107760 189138 107772
rect 191190 107760 191196 107772
rect 189132 107732 191196 107760
rect 189132 107720 189138 107732
rect 191190 107720 191196 107732
rect 191248 107720 191254 107772
rect 163498 107584 163504 107636
rect 163556 107624 163562 107636
rect 191742 107624 191748 107636
rect 163556 107596 191748 107624
rect 163556 107584 163562 107596
rect 191742 107584 191748 107596
rect 191800 107584 191806 107636
rect 226702 107584 226708 107636
rect 226760 107624 226766 107636
rect 284386 107624 284392 107636
rect 226760 107596 284392 107624
rect 226760 107584 226766 107596
rect 284386 107584 284392 107596
rect 284444 107624 284450 107636
rect 285030 107624 285036 107636
rect 284444 107596 285036 107624
rect 284444 107584 284450 107596
rect 285030 107584 285036 107596
rect 285088 107584 285094 107636
rect 187602 107516 187608 107568
rect 187660 107556 187666 107568
rect 189074 107556 189080 107568
rect 187660 107528 189080 107556
rect 187660 107516 187666 107528
rect 189074 107516 189080 107528
rect 189132 107516 189138 107568
rect 7558 106904 7564 106956
rect 7616 106944 7622 106956
rect 66990 106944 66996 106956
rect 7616 106916 66996 106944
rect 7616 106904 7622 106916
rect 66990 106904 66996 106916
rect 67048 106904 67054 106956
rect 97810 106904 97816 106956
rect 97868 106944 97874 106956
rect 169110 106944 169116 106956
rect 97868 106916 169116 106944
rect 97868 106904 97874 106916
rect 169110 106904 169116 106916
rect 169168 106904 169174 106956
rect 284386 106904 284392 106956
rect 284444 106944 284450 106956
rect 349154 106944 349160 106956
rect 284444 106916 349160 106944
rect 284444 106904 284450 106916
rect 349154 106904 349160 106916
rect 349212 106904 349218 106956
rect 96982 106632 96988 106684
rect 97040 106672 97046 106684
rect 100018 106672 100024 106684
rect 97040 106644 100024 106672
rect 97040 106632 97046 106644
rect 100018 106632 100024 106644
rect 100076 106632 100082 106684
rect 97534 106020 97540 106072
rect 97592 106060 97598 106072
rect 101490 106060 101496 106072
rect 97592 106032 101496 106060
rect 97592 106020 97598 106032
rect 101490 106020 101496 106032
rect 101548 106020 101554 106072
rect 96890 105884 96896 105936
rect 96948 105924 96954 105936
rect 98730 105924 98736 105936
rect 96948 105896 98736 105924
rect 96948 105884 96954 105896
rect 98730 105884 98736 105896
rect 98788 105884 98794 105936
rect 188338 105884 188344 105936
rect 188396 105924 188402 105936
rect 191742 105924 191748 105936
rect 188396 105896 191748 105924
rect 188396 105884 188402 105896
rect 191742 105884 191748 105896
rect 191800 105884 191806 105936
rect 48130 105544 48136 105596
rect 48188 105584 48194 105596
rect 64782 105584 64788 105596
rect 48188 105556 64788 105584
rect 48188 105544 48194 105556
rect 64782 105544 64788 105556
rect 64840 105584 64846 105596
rect 66530 105584 66536 105596
rect 64840 105556 66536 105584
rect 64840 105544 64846 105556
rect 66530 105544 66536 105556
rect 66588 105544 66594 105596
rect 111058 104904 111064 104916
rect 110708 104876 111064 104904
rect 56410 104796 56416 104848
rect 56468 104836 56474 104848
rect 66346 104836 66352 104848
rect 56468 104808 66352 104836
rect 56468 104796 56474 104808
rect 66346 104796 66352 104808
rect 66404 104796 66410 104848
rect 97718 104796 97724 104848
rect 97776 104836 97782 104848
rect 110708 104836 110736 104876
rect 111058 104864 111064 104876
rect 111116 104904 111122 104916
rect 177298 104904 177304 104916
rect 111116 104876 177304 104904
rect 111116 104864 111122 104876
rect 177298 104864 177304 104876
rect 177356 104864 177362 104916
rect 186222 104864 186228 104916
rect 186280 104904 186286 104916
rect 191742 104904 191748 104916
rect 186280 104876 191748 104904
rect 186280 104864 186286 104876
rect 191742 104864 191748 104876
rect 191800 104864 191806 104916
rect 226702 104864 226708 104916
rect 226760 104904 226766 104916
rect 226760 104876 277394 104904
rect 226760 104864 226766 104876
rect 97776 104808 110736 104836
rect 277366 104836 277394 104876
rect 278038 104836 278044 104848
rect 277366 104808 278044 104836
rect 97776 104796 97782 104808
rect 278038 104796 278044 104808
rect 278096 104836 278102 104848
rect 285674 104836 285680 104848
rect 278096 104808 285680 104836
rect 278096 104796 278102 104808
rect 285674 104796 285680 104808
rect 285732 104796 285738 104848
rect 96522 103504 96528 103556
rect 96580 103544 96586 103556
rect 178770 103544 178776 103556
rect 96580 103516 178776 103544
rect 96580 103504 96586 103516
rect 178770 103504 178776 103516
rect 178828 103504 178834 103556
rect 226518 103504 226524 103556
rect 226576 103544 226582 103556
rect 231946 103544 231952 103556
rect 226576 103516 231952 103544
rect 226576 103504 226582 103516
rect 231946 103504 231952 103516
rect 232004 103544 232010 103556
rect 280798 103544 280804 103556
rect 232004 103516 280804 103544
rect 232004 103504 232010 103516
rect 280798 103504 280804 103516
rect 280856 103504 280862 103556
rect 64690 103436 64696 103488
rect 64748 103476 64754 103488
rect 66622 103476 66628 103488
rect 64748 103448 66628 103476
rect 64748 103436 64754 103448
rect 66622 103436 66628 103448
rect 66680 103436 66686 103488
rect 97902 103028 97908 103080
rect 97960 103068 97966 103080
rect 99558 103068 99564 103080
rect 97960 103040 99564 103068
rect 97960 103028 97966 103040
rect 99558 103028 99564 103040
rect 99616 103028 99622 103080
rect 99558 102756 99564 102808
rect 99616 102796 99622 102808
rect 188338 102796 188344 102808
rect 99616 102768 188344 102796
rect 99616 102756 99622 102768
rect 188338 102756 188344 102768
rect 188396 102756 188402 102808
rect 226702 102756 226708 102808
rect 226760 102796 226766 102808
rect 227806 102796 227812 102808
rect 226760 102768 227812 102796
rect 226760 102756 226766 102768
rect 227806 102756 227812 102768
rect 227864 102796 227870 102808
rect 281534 102796 281540 102808
rect 227864 102768 281540 102796
rect 227864 102756 227870 102768
rect 281534 102756 281540 102768
rect 281592 102796 281598 102808
rect 309778 102796 309784 102808
rect 281592 102768 309784 102796
rect 281592 102756 281598 102768
rect 309778 102756 309784 102768
rect 309836 102756 309842 102808
rect 63402 102212 63408 102264
rect 63460 102252 63466 102264
rect 66070 102252 66076 102264
rect 63460 102224 66076 102252
rect 63460 102212 63466 102224
rect 66070 102212 66076 102224
rect 66128 102252 66134 102264
rect 66530 102252 66536 102264
rect 66128 102224 66536 102252
rect 66128 102212 66134 102224
rect 66530 102212 66536 102224
rect 66588 102212 66594 102264
rect 67358 102144 67364 102196
rect 67416 102184 67422 102196
rect 67634 102184 67640 102196
rect 67416 102156 67640 102184
rect 67416 102144 67422 102156
rect 67634 102144 67640 102156
rect 67692 102144 67698 102196
rect 100662 102144 100668 102196
rect 100720 102184 100726 102196
rect 184290 102184 184296 102196
rect 100720 102156 184296 102184
rect 100720 102144 100726 102156
rect 184290 102144 184296 102156
rect 184348 102144 184354 102196
rect 186958 102144 186964 102196
rect 187016 102184 187022 102196
rect 191650 102184 191656 102196
rect 187016 102156 191656 102184
rect 187016 102144 187022 102156
rect 191650 102144 191656 102156
rect 191708 102144 191714 102196
rect 226702 102144 226708 102196
rect 226760 102184 226766 102196
rect 237558 102184 237564 102196
rect 226760 102156 237564 102184
rect 226760 102144 226766 102156
rect 237558 102144 237564 102156
rect 237616 102144 237622 102196
rect 226334 102076 226340 102128
rect 226392 102116 226398 102128
rect 266354 102116 266360 102128
rect 226392 102088 266360 102116
rect 226392 102076 226398 102088
rect 266354 102076 266360 102088
rect 266412 102076 266418 102128
rect 97902 102008 97908 102060
rect 97960 102048 97966 102060
rect 130562 102048 130568 102060
rect 97960 102020 130568 102048
rect 97960 102008 97966 102020
rect 130562 102008 130568 102020
rect 130620 102008 130626 102060
rect 130562 101464 130568 101516
rect 130620 101504 130626 101516
rect 148502 101504 148508 101516
rect 130620 101476 148508 101504
rect 130620 101464 130626 101476
rect 148502 101464 148508 101476
rect 148560 101464 148566 101516
rect 113910 101396 113916 101448
rect 113968 101436 113974 101448
rect 158622 101436 158628 101448
rect 113968 101408 158628 101436
rect 113968 101396 113974 101408
rect 158622 101396 158628 101408
rect 158680 101436 158686 101448
rect 181990 101436 181996 101448
rect 158680 101408 181996 101436
rect 158680 101396 158686 101408
rect 181990 101396 181996 101408
rect 182048 101396 182054 101448
rect 61930 100852 61936 100904
rect 61988 100892 61994 100904
rect 66806 100892 66812 100904
rect 61988 100864 66812 100892
rect 61988 100852 61994 100864
rect 66806 100852 66812 100864
rect 66864 100852 66870 100904
rect 181990 100716 181996 100768
rect 182048 100756 182054 100768
rect 191650 100756 191656 100768
rect 182048 100728 191656 100756
rect 182048 100716 182054 100728
rect 191650 100716 191656 100728
rect 191708 100716 191714 100768
rect 97902 100648 97908 100700
rect 97960 100688 97966 100700
rect 100662 100688 100668 100700
rect 97960 100660 100668 100688
rect 97960 100648 97966 100660
rect 100662 100648 100668 100660
rect 100720 100648 100726 100700
rect 185578 100648 185584 100700
rect 185636 100688 185642 100700
rect 190638 100688 190644 100700
rect 185636 100660 190644 100688
rect 185636 100648 185642 100660
rect 190638 100648 190644 100660
rect 190696 100648 190702 100700
rect 60642 99628 60648 99680
rect 60700 99668 60706 99680
rect 63402 99668 63408 99680
rect 60700 99640 63408 99668
rect 60700 99628 60706 99640
rect 63402 99628 63408 99640
rect 63460 99668 63466 99680
rect 66806 99668 66812 99680
rect 63460 99640 66812 99668
rect 63460 99628 63466 99640
rect 66806 99628 66812 99640
rect 66864 99628 66870 99680
rect 97534 99356 97540 99408
rect 97592 99396 97598 99408
rect 131022 99396 131028 99408
rect 97592 99368 131028 99396
rect 97592 99356 97598 99368
rect 131022 99356 131028 99368
rect 131080 99356 131086 99408
rect 226426 99356 226432 99408
rect 226484 99396 226490 99408
rect 229186 99396 229192 99408
rect 226484 99368 229192 99396
rect 226484 99356 226490 99368
rect 229186 99356 229192 99368
rect 229244 99396 229250 99408
rect 322198 99396 322204 99408
rect 229244 99368 322204 99396
rect 229244 99356 229250 99368
rect 322198 99356 322204 99368
rect 322256 99356 322262 99408
rect 62022 99288 62028 99340
rect 62080 99328 62086 99340
rect 66806 99328 66812 99340
rect 62080 99300 66812 99328
rect 62080 99288 62086 99300
rect 66806 99288 66812 99300
rect 66864 99288 66870 99340
rect 237374 98676 237380 98728
rect 237432 98716 237438 98728
rect 250530 98716 250536 98728
rect 237432 98688 250536 98716
rect 237432 98676 237438 98688
rect 250530 98676 250536 98688
rect 250588 98676 250594 98728
rect 226518 98608 226524 98660
rect 226576 98648 226582 98660
rect 264974 98648 264980 98660
rect 226576 98620 264980 98648
rect 226576 98608 226582 98620
rect 264974 98608 264980 98620
rect 265032 98608 265038 98660
rect 96890 98336 96896 98388
rect 96948 98376 96954 98388
rect 98914 98376 98920 98388
rect 96948 98348 98920 98376
rect 96948 98336 96954 98348
rect 98914 98336 98920 98348
rect 98972 98336 98978 98388
rect 100110 98064 100116 98116
rect 100168 98104 100174 98116
rect 164142 98104 164148 98116
rect 100168 98076 164148 98104
rect 100168 98064 100174 98076
rect 164142 98064 164148 98076
rect 164200 98104 164206 98116
rect 164878 98104 164884 98116
rect 164200 98076 164884 98104
rect 164200 98064 164206 98076
rect 164878 98064 164884 98076
rect 164936 98064 164942 98116
rect 184382 98064 184388 98116
rect 184440 98104 184446 98116
rect 191650 98104 191656 98116
rect 184440 98076 191656 98104
rect 184440 98064 184446 98076
rect 191650 98064 191656 98076
rect 191708 98064 191714 98116
rect 97350 97996 97356 98048
rect 97408 98036 97414 98048
rect 189810 98036 189816 98048
rect 97408 98008 189816 98036
rect 97408 97996 97414 98008
rect 189810 97996 189816 98008
rect 189868 97996 189874 98048
rect 181530 97928 181536 97980
rect 181588 97968 181594 97980
rect 190638 97968 190644 97980
rect 181588 97940 190644 97968
rect 181588 97928 181594 97940
rect 190638 97928 190644 97940
rect 190696 97928 190702 97980
rect 96890 96840 96896 96892
rect 96948 96880 96954 96892
rect 98822 96880 98828 96892
rect 96948 96852 98828 96880
rect 96948 96840 96954 96852
rect 98822 96840 98828 96852
rect 98880 96840 98886 96892
rect 3050 96636 3056 96688
rect 3108 96676 3114 96688
rect 62758 96676 62764 96688
rect 3108 96648 62764 96676
rect 3108 96636 3114 96648
rect 62758 96636 62764 96648
rect 62816 96636 62822 96688
rect 97902 96636 97908 96688
rect 97960 96676 97966 96688
rect 188430 96676 188436 96688
rect 97960 96648 188436 96676
rect 97960 96636 97966 96648
rect 188430 96636 188436 96648
rect 188488 96636 188494 96688
rect 226518 95956 226524 96008
rect 226576 95996 226582 96008
rect 228358 95996 228364 96008
rect 226576 95968 228364 95996
rect 226576 95956 226582 95968
rect 228358 95956 228364 95968
rect 228416 95956 228422 96008
rect 95418 95208 95424 95260
rect 95476 95248 95482 95260
rect 193122 95248 193128 95260
rect 95476 95220 193128 95248
rect 95476 95208 95482 95220
rect 193122 95208 193128 95220
rect 193180 95208 193186 95260
rect 52362 95140 52368 95192
rect 52420 95180 52426 95192
rect 66806 95180 66812 95192
rect 52420 95152 66812 95180
rect 52420 95140 52426 95152
rect 66806 95140 66812 95152
rect 66864 95140 66870 95192
rect 95970 95140 95976 95192
rect 96028 95180 96034 95192
rect 182082 95180 182088 95192
rect 96028 95152 182088 95180
rect 96028 95140 96034 95152
rect 182082 95140 182088 95152
rect 182140 95140 182146 95192
rect 96982 94460 96988 94512
rect 97040 94500 97046 94512
rect 102226 94500 102232 94512
rect 97040 94472 102232 94500
rect 97040 94460 97046 94472
rect 102226 94460 102232 94472
rect 102284 94460 102290 94512
rect 182082 94460 182088 94512
rect 182140 94500 182146 94512
rect 193398 94500 193404 94512
rect 182140 94472 193404 94500
rect 182140 94460 182146 94472
rect 193398 94460 193404 94472
rect 193456 94460 193462 94512
rect 227622 94460 227628 94512
rect 227680 94500 227686 94512
rect 263686 94500 263692 94512
rect 227680 94472 263692 94500
rect 227680 94460 227686 94472
rect 263686 94460 263692 94472
rect 263744 94460 263750 94512
rect 226610 94392 226616 94444
rect 226668 94432 226674 94444
rect 228358 94432 228364 94444
rect 226668 94404 228364 94432
rect 226668 94392 226674 94404
rect 228358 94392 228364 94404
rect 228416 94392 228422 94444
rect 53742 93780 53748 93832
rect 53800 93820 53806 93832
rect 68002 93820 68008 93832
rect 53800 93792 68008 93820
rect 53800 93780 53806 93792
rect 68002 93780 68008 93792
rect 68060 93780 68066 93832
rect 97902 93780 97908 93832
rect 97960 93820 97966 93832
rect 108390 93820 108396 93832
rect 97960 93792 108396 93820
rect 97960 93780 97966 93792
rect 108390 93780 108396 93792
rect 108448 93780 108454 93832
rect 171042 93100 171048 93152
rect 171100 93140 171106 93152
rect 183554 93140 183560 93152
rect 171100 93112 183560 93140
rect 171100 93100 171106 93112
rect 183554 93100 183560 93112
rect 183612 93140 183618 93152
rect 191742 93140 191748 93152
rect 183612 93112 191748 93140
rect 183612 93100 183618 93112
rect 191742 93100 191748 93112
rect 191800 93100 191806 93152
rect 231302 93100 231308 93152
rect 231360 93140 231366 93152
rect 249150 93140 249156 93152
rect 231360 93112 249156 93140
rect 231360 93100 231366 93112
rect 249150 93100 249156 93112
rect 249208 93100 249214 93152
rect 250530 93100 250536 93152
rect 250588 93140 250594 93152
rect 331214 93140 331220 93152
rect 250588 93112 331220 93140
rect 250588 93100 250594 93112
rect 331214 93100 331220 93112
rect 331272 93100 331278 93152
rect 69014 92896 69020 92948
rect 69072 92896 69078 92948
rect 67358 92828 67364 92880
rect 67416 92868 67422 92880
rect 68462 92868 68468 92880
rect 67416 92840 68468 92868
rect 67416 92828 67422 92840
rect 68462 92828 68468 92840
rect 68520 92828 68526 92880
rect 69032 92732 69060 92896
rect 70256 92732 70262 92744
rect 69032 92704 70262 92732
rect 70256 92692 70262 92704
rect 70314 92692 70320 92744
rect 91784 92692 91790 92744
rect 91842 92732 91848 92744
rect 95234 92732 95240 92744
rect 91842 92704 95240 92732
rect 91842 92692 91848 92704
rect 95234 92692 95240 92704
rect 95292 92692 95298 92744
rect 88656 92624 88662 92676
rect 88714 92664 88720 92676
rect 89622 92664 89628 92676
rect 88714 92636 89628 92664
rect 88714 92624 88720 92636
rect 89622 92624 89628 92636
rect 89680 92624 89686 92676
rect 90128 92624 90134 92676
rect 90186 92624 90192 92676
rect 74626 92556 74632 92608
rect 74684 92596 74690 92608
rect 75776 92596 75782 92608
rect 74684 92568 75782 92596
rect 74684 92556 74690 92568
rect 75776 92556 75782 92568
rect 75834 92556 75840 92608
rect 80146 92556 80152 92608
rect 80204 92596 80210 92608
rect 80928 92596 80934 92608
rect 80204 92568 80934 92596
rect 80204 92556 80210 92568
rect 80928 92556 80934 92568
rect 80986 92556 80992 92608
rect 50890 92352 50896 92404
rect 50948 92392 50954 92404
rect 72786 92392 72792 92404
rect 50948 92364 72792 92392
rect 50948 92352 50954 92364
rect 72786 92352 72792 92364
rect 72844 92352 72850 92404
rect 90146 92392 90174 92624
rect 126514 92488 126520 92540
rect 126572 92528 126578 92540
rect 218790 92528 218796 92540
rect 126572 92500 218796 92528
rect 126572 92488 126578 92500
rect 218790 92488 218796 92500
rect 218848 92488 218854 92540
rect 221918 92488 221924 92540
rect 221976 92528 221982 92540
rect 232498 92528 232504 92540
rect 221976 92500 232504 92528
rect 221976 92488 221982 92500
rect 232498 92488 232504 92500
rect 232556 92488 232562 92540
rect 126532 92392 126560 92488
rect 184290 92420 184296 92472
rect 184348 92460 184354 92472
rect 229186 92460 229192 92472
rect 184348 92432 229192 92460
rect 184348 92420 184354 92432
rect 229186 92420 229192 92432
rect 229244 92420 229250 92472
rect 90146 92364 126560 92392
rect 213178 92352 213184 92404
rect 213236 92392 213242 92404
rect 242250 92392 242256 92404
rect 213236 92364 242256 92392
rect 213236 92352 213242 92364
rect 242250 92352 242256 92364
rect 242308 92352 242314 92404
rect 67450 92284 67456 92336
rect 67508 92324 67514 92336
rect 184382 92324 184388 92336
rect 67508 92296 184388 92324
rect 67508 92284 67514 92296
rect 184382 92284 184388 92296
rect 184440 92284 184446 92336
rect 193122 91740 193128 91792
rect 193180 91780 193186 91792
rect 202138 91780 202144 91792
rect 193180 91752 202144 91780
rect 193180 91740 193186 91752
rect 202138 91740 202144 91752
rect 202196 91740 202202 91792
rect 65886 90992 65892 91044
rect 65944 91032 65950 91044
rect 71130 91032 71136 91044
rect 65944 91004 71136 91032
rect 65944 90992 65950 91004
rect 71130 90992 71136 91004
rect 71188 90992 71194 91044
rect 84654 90992 84660 91044
rect 84712 91032 84718 91044
rect 116118 91032 116124 91044
rect 84712 91004 116124 91032
rect 84712 90992 84718 91004
rect 116118 90992 116124 91004
rect 116176 91032 116182 91044
rect 212442 91032 212448 91044
rect 116176 91004 212448 91032
rect 116176 90992 116182 91004
rect 212442 90992 212448 91004
rect 212500 90992 212506 91044
rect 221366 90992 221372 91044
rect 221424 91032 221430 91044
rect 258074 91032 258080 91044
rect 221424 91004 258080 91032
rect 221424 90992 221430 91004
rect 258074 90992 258080 91004
rect 258132 90992 258138 91044
rect 85206 90312 85212 90364
rect 85264 90352 85270 90364
rect 94498 90352 94504 90364
rect 85264 90324 94504 90352
rect 85264 90312 85270 90324
rect 94498 90312 94504 90324
rect 94556 90312 94562 90364
rect 213454 90312 213460 90364
rect 213512 90352 213518 90364
rect 235258 90352 235264 90364
rect 213512 90324 235264 90352
rect 213512 90312 213518 90324
rect 235258 90312 235264 90324
rect 235316 90312 235322 90364
rect 68922 90244 68928 90296
rect 68980 90284 68986 90296
rect 71038 90284 71044 90296
rect 68980 90256 71044 90284
rect 68980 90244 68986 90256
rect 71038 90244 71044 90256
rect 71096 90244 71102 90296
rect 223758 90244 223764 90296
rect 223816 90284 223822 90296
rect 224862 90284 224868 90296
rect 223816 90256 224868 90284
rect 223816 90244 223822 90256
rect 224862 90244 224868 90256
rect 224920 90244 224926 90296
rect 105538 89700 105544 89752
rect 105596 89740 105602 89752
rect 106366 89740 106372 89752
rect 105596 89712 106372 89740
rect 105596 89700 105602 89712
rect 106366 89700 106372 89712
rect 106424 89700 106430 89752
rect 127618 89700 127624 89752
rect 127676 89740 127682 89752
rect 128354 89740 128360 89752
rect 127676 89712 128360 89740
rect 127676 89700 127682 89712
rect 128354 89700 128360 89712
rect 128412 89700 128418 89752
rect 245654 89700 245660 89752
rect 245712 89740 245718 89752
rect 246298 89740 246304 89752
rect 245712 89712 246304 89740
rect 245712 89700 245718 89712
rect 246298 89700 246304 89712
rect 246356 89740 246362 89752
rect 580258 89740 580264 89752
rect 246356 89712 580264 89740
rect 246356 89700 246362 89712
rect 580258 89700 580264 89712
rect 580316 89700 580322 89752
rect 49602 89632 49608 89684
rect 49660 89672 49666 89684
rect 79410 89672 79416 89684
rect 49660 89644 79416 89672
rect 49660 89632 49666 89644
rect 79410 89632 79416 89644
rect 79468 89632 79474 89684
rect 85574 89632 85580 89684
rect 85632 89672 85638 89684
rect 117314 89672 117320 89684
rect 85632 89644 117320 89672
rect 85632 89632 85638 89644
rect 117314 89632 117320 89644
rect 117372 89672 117378 89684
rect 117774 89672 117780 89684
rect 117372 89644 117780 89672
rect 117372 89632 117378 89644
rect 117774 89632 117780 89644
rect 117832 89632 117838 89684
rect 124122 89632 124128 89684
rect 124180 89672 124186 89684
rect 217686 89672 217692 89684
rect 124180 89644 217692 89672
rect 124180 89632 124186 89644
rect 217686 89632 217692 89644
rect 217744 89632 217750 89684
rect 220630 89632 220636 89684
rect 220688 89672 220694 89684
rect 273346 89672 273352 89684
rect 220688 89644 273352 89672
rect 220688 89632 220694 89644
rect 273346 89632 273352 89644
rect 273404 89632 273410 89684
rect 84102 89564 84108 89616
rect 84160 89604 84166 89616
rect 98730 89604 98736 89616
rect 84160 89576 98736 89604
rect 84160 89564 84166 89576
rect 98730 89564 98736 89576
rect 98788 89564 98794 89616
rect 193398 89564 193404 89616
rect 193456 89604 193462 89616
rect 199378 89604 199384 89616
rect 193456 89576 199384 89604
rect 193456 89564 193462 89576
rect 199378 89564 199384 89576
rect 199436 89564 199442 89616
rect 203702 89564 203708 89616
rect 203760 89604 203766 89616
rect 284294 89604 284300 89616
rect 203760 89576 284300 89604
rect 203760 89564 203766 89576
rect 284294 89564 284300 89576
rect 284352 89564 284358 89616
rect 123570 89224 123576 89276
rect 123628 89264 123634 89276
rect 124122 89264 124128 89276
rect 123628 89236 124128 89264
rect 123628 89224 123634 89236
rect 124122 89224 124128 89236
rect 124180 89224 124186 89276
rect 284294 88952 284300 89004
rect 284352 88992 284358 89004
rect 582834 88992 582840 89004
rect 284352 88964 582840 88992
rect 284352 88952 284358 88964
rect 582834 88952 582840 88964
rect 582892 88952 582898 89004
rect 67266 88272 67272 88324
rect 67324 88312 67330 88324
rect 113910 88312 113916 88324
rect 67324 88284 113916 88312
rect 67324 88272 67330 88284
rect 113910 88272 113916 88284
rect 113968 88272 113974 88324
rect 117774 88272 117780 88324
rect 117832 88312 117838 88324
rect 213454 88312 213460 88324
rect 117832 88284 213460 88312
rect 117832 88272 117838 88284
rect 213454 88272 213460 88284
rect 213512 88272 213518 88324
rect 214558 88272 214564 88324
rect 214616 88312 214622 88324
rect 262214 88312 262220 88324
rect 214616 88284 262220 88312
rect 214616 88272 214622 88284
rect 262214 88272 262220 88284
rect 262272 88272 262278 88324
rect 60458 88204 60464 88256
rect 60516 88244 60522 88256
rect 82630 88244 82636 88256
rect 60516 88216 82636 88244
rect 60516 88204 60522 88216
rect 82630 88204 82636 88216
rect 82688 88244 82694 88256
rect 83458 88244 83464 88256
rect 82688 88216 83464 88244
rect 82688 88204 82694 88216
rect 83458 88204 83464 88216
rect 83516 88204 83522 88256
rect 86678 88204 86684 88256
rect 86736 88244 86742 88256
rect 100754 88244 100760 88256
rect 86736 88216 100760 88244
rect 86736 88204 86742 88216
rect 100754 88204 100760 88216
rect 100812 88204 100818 88256
rect 188522 88204 188528 88256
rect 188580 88244 188586 88256
rect 196066 88244 196072 88256
rect 188580 88216 196072 88244
rect 188580 88204 188586 88216
rect 196066 88204 196072 88216
rect 196124 88204 196130 88256
rect 206370 88204 206376 88256
rect 206428 88244 206434 88256
rect 207382 88244 207388 88256
rect 206428 88216 207388 88244
rect 206428 88204 206434 88216
rect 207382 88204 207388 88216
rect 207440 88204 207446 88256
rect 215846 88204 215852 88256
rect 215904 88244 215910 88256
rect 216030 88244 216036 88256
rect 215904 88216 216036 88244
rect 215904 88204 215910 88216
rect 216030 88204 216036 88216
rect 216088 88244 216094 88256
rect 242158 88244 242164 88256
rect 216088 88216 242164 88244
rect 216088 88204 216094 88216
rect 242158 88204 242164 88216
rect 242216 88204 242222 88256
rect 89806 86912 89812 86964
rect 89864 86952 89870 86964
rect 124306 86952 124312 86964
rect 89864 86924 124312 86952
rect 89864 86912 89870 86924
rect 124306 86912 124312 86924
rect 124364 86952 124370 86964
rect 218238 86952 218244 86964
rect 124364 86924 218244 86952
rect 124364 86912 124370 86924
rect 218238 86912 218244 86924
rect 218296 86912 218302 86964
rect 219526 86912 219532 86964
rect 219584 86952 219590 86964
rect 220078 86952 220084 86964
rect 219584 86924 220084 86952
rect 219584 86912 219590 86924
rect 220078 86912 220084 86924
rect 220136 86952 220142 86964
rect 245654 86952 245660 86964
rect 220136 86924 245660 86952
rect 220136 86912 220142 86924
rect 245654 86912 245660 86924
rect 245712 86912 245718 86964
rect 73798 86844 73804 86896
rect 73856 86884 73862 86896
rect 73856 86856 84194 86884
rect 73856 86844 73862 86856
rect 84166 86816 84194 86856
rect 185118 86844 185124 86896
rect 185176 86884 185182 86896
rect 227714 86884 227720 86896
rect 185176 86856 227720 86884
rect 185176 86844 185182 86856
rect 227714 86844 227720 86856
rect 227772 86844 227778 86896
rect 95970 86816 95976 86828
rect 84166 86788 95976 86816
rect 95970 86776 95976 86788
rect 96028 86776 96034 86828
rect 228358 86232 228364 86284
rect 228416 86272 228422 86284
rect 241514 86272 241520 86284
rect 228416 86244 241520 86272
rect 228416 86232 228422 86244
rect 241514 86232 241520 86244
rect 241572 86232 241578 86284
rect 197354 85552 197360 85604
rect 197412 85592 197418 85604
rect 197998 85592 198004 85604
rect 197412 85564 198004 85592
rect 197412 85552 197418 85564
rect 197998 85552 198004 85564
rect 198056 85552 198062 85604
rect 52362 85484 52368 85536
rect 52420 85524 52426 85536
rect 52546 85524 52552 85536
rect 52420 85496 52552 85524
rect 52420 85484 52426 85496
rect 52546 85484 52552 85496
rect 52604 85484 52610 85536
rect 87230 85484 87236 85536
rect 87288 85524 87294 85536
rect 117958 85524 117964 85536
rect 87288 85496 117964 85524
rect 87288 85484 87294 85496
rect 117958 85484 117964 85496
rect 118016 85524 118022 85536
rect 215386 85524 215392 85536
rect 118016 85496 215392 85524
rect 118016 85484 118022 85496
rect 215386 85484 215392 85496
rect 215444 85484 215450 85536
rect 65978 85416 65984 85468
rect 66036 85456 66042 85468
rect 159358 85456 159364 85468
rect 66036 85428 159364 85456
rect 66036 85416 66042 85428
rect 159358 85416 159364 85428
rect 159416 85416 159422 85468
rect 238478 84872 238484 84924
rect 238536 84912 238542 84924
rect 307018 84912 307024 84924
rect 238536 84884 307024 84912
rect 238536 84872 238542 84884
rect 307018 84872 307024 84884
rect 307076 84872 307082 84924
rect 191742 84804 191748 84856
rect 191800 84844 191806 84856
rect 270586 84844 270592 84856
rect 191800 84816 270592 84844
rect 191800 84804 191806 84816
rect 270586 84804 270592 84816
rect 270644 84804 270650 84856
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 52362 84232 52368 84244
rect 3384 84204 52368 84232
rect 3384 84192 3390 84204
rect 52362 84192 52368 84204
rect 52420 84192 52426 84244
rect 69014 84124 69020 84176
rect 69072 84164 69078 84176
rect 169018 84164 169024 84176
rect 69072 84136 169024 84164
rect 69072 84124 69078 84136
rect 169018 84124 169024 84136
rect 169076 84164 169082 84176
rect 193306 84164 193312 84176
rect 169076 84136 193312 84164
rect 169076 84124 169082 84136
rect 193306 84124 193312 84136
rect 193364 84124 193370 84176
rect 216674 84124 216680 84176
rect 216732 84164 216738 84176
rect 261478 84164 261484 84176
rect 216732 84136 261484 84164
rect 216732 84124 216738 84136
rect 261478 84124 261484 84136
rect 261536 84124 261542 84176
rect 116026 84056 116032 84108
rect 116084 84096 116090 84108
rect 213914 84096 213920 84108
rect 116084 84068 213920 84096
rect 116084 84056 116090 84068
rect 213914 84056 213920 84068
rect 213972 84056 213978 84108
rect 222286 83036 222292 83088
rect 222344 83076 222350 83088
rect 222838 83076 222844 83088
rect 222344 83048 222844 83076
rect 222344 83036 222350 83048
rect 222838 83036 222844 83048
rect 222896 83036 222902 83088
rect 193306 82832 193312 82884
rect 193364 82872 193370 82884
rect 193950 82872 193956 82884
rect 193364 82844 193956 82872
rect 193364 82832 193370 82844
rect 193950 82832 193956 82844
rect 194008 82832 194014 82884
rect 216674 82832 216680 82884
rect 216732 82872 216738 82884
rect 217318 82872 217324 82884
rect 216732 82844 217324 82872
rect 216732 82832 216738 82844
rect 217318 82832 217324 82844
rect 217376 82832 217382 82884
rect 222838 82832 222844 82884
rect 222896 82872 222902 82884
rect 339494 82872 339500 82884
rect 222896 82844 339500 82872
rect 222896 82832 222902 82844
rect 339494 82832 339500 82844
rect 339552 82832 339558 82884
rect 88334 82764 88340 82816
rect 88392 82804 88398 82816
rect 123570 82804 123576 82816
rect 88392 82776 123576 82804
rect 88392 82764 88398 82776
rect 123570 82764 123576 82776
rect 123628 82764 123634 82816
rect 188338 82764 188344 82816
rect 188396 82804 188402 82816
rect 227806 82804 227812 82816
rect 188396 82776 227812 82804
rect 188396 82764 188402 82776
rect 227806 82764 227812 82776
rect 227864 82764 227870 82816
rect 80238 82696 80244 82748
rect 80296 82736 80302 82748
rect 105538 82736 105544 82748
rect 80296 82708 105544 82736
rect 80296 82696 80302 82708
rect 105538 82696 105544 82708
rect 105596 82696 105602 82748
rect 178034 82696 178040 82748
rect 178092 82736 178098 82748
rect 179322 82736 179328 82748
rect 178092 82708 179328 82736
rect 178092 82696 178098 82708
rect 179322 82696 179328 82708
rect 179380 82736 179386 82748
rect 200114 82736 200120 82748
rect 179380 82708 200120 82736
rect 179380 82696 179386 82708
rect 200114 82696 200120 82708
rect 200172 82736 200178 82748
rect 201402 82736 201408 82748
rect 200172 82708 201408 82736
rect 200172 82696 200178 82708
rect 201402 82696 201408 82708
rect 201460 82696 201466 82748
rect 201402 82084 201408 82136
rect 201460 82124 201466 82136
rect 245654 82124 245660 82136
rect 201460 82096 245660 82124
rect 201460 82084 201466 82096
rect 245654 82084 245660 82096
rect 245712 82084 245718 82136
rect 52362 81336 52368 81388
rect 52420 81376 52426 81388
rect 153838 81376 153844 81388
rect 52420 81348 153844 81376
rect 52420 81336 52426 81348
rect 153838 81336 153844 81348
rect 153896 81336 153902 81388
rect 178770 81336 178776 81388
rect 178828 81376 178834 81388
rect 231946 81376 231952 81388
rect 178828 81348 231952 81376
rect 178828 81336 178834 81348
rect 231946 81336 231952 81348
rect 232004 81336 232010 81388
rect 71866 81268 71872 81320
rect 71924 81308 71930 81320
rect 172514 81308 172520 81320
rect 71924 81280 172520 81308
rect 71924 81268 71930 81280
rect 172514 81268 172520 81280
rect 172572 81308 172578 81320
rect 173802 81308 173808 81320
rect 172572 81280 173808 81308
rect 172572 81268 172578 81280
rect 173802 81268 173808 81280
rect 173860 81268 173866 81320
rect 164142 81200 164148 81252
rect 164200 81240 164206 81252
rect 195974 81240 195980 81252
rect 164200 81212 195980 81240
rect 164200 81200 164206 81212
rect 195974 81200 195980 81212
rect 196032 81200 196038 81252
rect 210510 80656 210516 80708
rect 210568 80696 210574 80708
rect 582926 80696 582932 80708
rect 210568 80668 582932 80696
rect 210568 80656 210574 80668
rect 582926 80656 582932 80668
rect 582984 80656 582990 80708
rect 195974 80044 195980 80096
rect 196032 80084 196038 80096
rect 196618 80084 196624 80096
rect 196032 80056 196624 80084
rect 196032 80044 196038 80056
rect 196618 80044 196624 80056
rect 196676 80044 196682 80096
rect 80054 79976 80060 80028
rect 80112 80016 80118 80028
rect 161474 80016 161480 80028
rect 80112 79988 161480 80016
rect 80112 79976 80118 79988
rect 161446 79976 161480 79988
rect 161532 79976 161538 80028
rect 177298 79976 177304 80028
rect 177356 80016 177362 80028
rect 224954 80016 224960 80028
rect 177356 79988 224960 80016
rect 177356 79976 177362 79988
rect 224954 79976 224960 79988
rect 225012 79976 225018 80028
rect 62758 79908 62764 79960
rect 62816 79948 62822 79960
rect 96614 79948 96620 79960
rect 62816 79920 96620 79948
rect 62816 79908 62822 79920
rect 96614 79908 96620 79920
rect 96672 79908 96678 79960
rect 161446 79948 161474 79976
rect 205634 79948 205640 79960
rect 161446 79920 205640 79948
rect 205634 79908 205640 79920
rect 205692 79908 205698 79960
rect 205634 79500 205640 79552
rect 205692 79540 205698 79552
rect 206278 79540 206284 79552
rect 205692 79512 206284 79540
rect 205692 79500 205698 79512
rect 206278 79500 206284 79512
rect 206336 79500 206342 79552
rect 98638 79296 98644 79348
rect 98696 79336 98702 79348
rect 113818 79336 113824 79348
rect 98696 79308 113824 79336
rect 98696 79296 98702 79308
rect 113818 79296 113824 79308
rect 113876 79296 113882 79348
rect 75822 78616 75828 78668
rect 75880 78656 75886 78668
rect 178034 78656 178040 78668
rect 75880 78628 178040 78656
rect 75880 78616 75886 78628
rect 178034 78616 178040 78628
rect 178092 78616 178098 78668
rect 180150 78616 180156 78668
rect 180208 78656 180214 78668
rect 225046 78656 225052 78668
rect 180208 78628 225052 78656
rect 180208 78616 180214 78628
rect 225046 78616 225052 78628
rect 225104 78616 225110 78668
rect 173802 78548 173808 78600
rect 173860 78588 173866 78600
rect 197446 78588 197452 78600
rect 173860 78560 197452 78588
rect 173860 78548 173866 78560
rect 197446 78548 197452 78560
rect 197504 78588 197510 78600
rect 197998 78588 198004 78600
rect 197504 78560 198004 78588
rect 197504 78548 197510 78560
rect 197998 78548 198004 78560
rect 198056 78548 198062 78600
rect 198734 77936 198740 77988
rect 198792 77976 198798 77988
rect 240134 77976 240140 77988
rect 198792 77948 240140 77976
rect 198792 77936 198798 77948
rect 240134 77936 240140 77948
rect 240192 77936 240198 77988
rect 288342 77936 288348 77988
rect 288400 77976 288406 77988
rect 345014 77976 345020 77988
rect 288400 77948 345020 77976
rect 288400 77936 288406 77948
rect 345014 77936 345020 77948
rect 345072 77936 345078 77988
rect 92474 77188 92480 77240
rect 92532 77228 92538 77240
rect 127618 77228 127624 77240
rect 92532 77200 127624 77228
rect 92532 77188 92538 77200
rect 127618 77188 127624 77200
rect 127676 77188 127682 77240
rect 148502 77188 148508 77240
rect 148560 77228 148566 77240
rect 237558 77228 237564 77240
rect 148560 77200 237564 77228
rect 148560 77188 148566 77200
rect 237558 77188 237564 77200
rect 237616 77228 237622 77240
rect 238018 77228 238024 77240
rect 237616 77200 238024 77228
rect 237616 77188 237622 77200
rect 238018 77188 238024 77200
rect 238076 77188 238082 77240
rect 173250 77120 173256 77172
rect 173308 77160 173314 77172
rect 244274 77160 244280 77172
rect 173308 77132 244280 77160
rect 173308 77120 173314 77132
rect 244274 77120 244280 77132
rect 244332 77120 244338 77172
rect 70302 76508 70308 76560
rect 70360 76548 70366 76560
rect 166350 76548 166356 76560
rect 70360 76520 166356 76548
rect 70360 76508 70366 76520
rect 166350 76508 166356 76520
rect 166408 76508 166414 76560
rect 280062 76508 280068 76560
rect 280120 76548 280126 76560
rect 292666 76548 292672 76560
rect 280120 76520 292672 76548
rect 280120 76508 280126 76520
rect 292666 76508 292672 76520
rect 292724 76508 292730 76560
rect 244274 76304 244280 76356
rect 244332 76344 244338 76356
rect 245010 76344 245016 76356
rect 244332 76316 245016 76344
rect 244332 76304 244338 76316
rect 245010 76304 245016 76316
rect 245068 76304 245074 76356
rect 169110 75828 169116 75880
rect 169168 75868 169174 75880
rect 229094 75868 229100 75880
rect 169168 75840 229100 75868
rect 169168 75828 169174 75840
rect 229094 75828 229100 75840
rect 229152 75828 229158 75880
rect 193214 75760 193220 75812
rect 193272 75800 193278 75812
rect 193858 75800 193864 75812
rect 193272 75772 193864 75800
rect 193272 75760 193278 75772
rect 193858 75760 193864 75772
rect 193916 75800 193922 75812
rect 244918 75800 244924 75812
rect 193916 75772 244924 75800
rect 193916 75760 193922 75772
rect 244918 75760 244924 75772
rect 244976 75760 244982 75812
rect 74534 75148 74540 75200
rect 74592 75188 74598 75200
rect 167638 75188 167644 75200
rect 74592 75160 167644 75188
rect 74592 75148 74598 75160
rect 167638 75148 167644 75160
rect 167696 75148 167702 75200
rect 255222 74536 255228 74588
rect 255280 74576 255286 74588
rect 318058 74576 318064 74588
rect 255280 74548 318064 74576
rect 255280 74536 255286 74548
rect 318058 74536 318064 74548
rect 318116 74536 318122 74588
rect 61930 74468 61936 74520
rect 61988 74508 61994 74520
rect 186958 74508 186964 74520
rect 61988 74480 186964 74508
rect 61988 74468 61994 74480
rect 186958 74468 186964 74480
rect 187016 74468 187022 74520
rect 201494 74468 201500 74520
rect 201552 74508 201558 74520
rect 255240 74508 255268 74536
rect 201552 74480 255268 74508
rect 201552 74468 201558 74480
rect 166350 74400 166356 74452
rect 166408 74440 166414 74452
rect 194594 74440 194600 74452
rect 166408 74412 194600 74440
rect 166408 74400 166414 74412
rect 194594 74400 194600 74412
rect 194652 74400 194658 74452
rect 85574 73788 85580 73840
rect 85632 73828 85638 73840
rect 160830 73828 160836 73840
rect 85632 73800 160836 73828
rect 85632 73788 85638 73800
rect 160830 73788 160836 73800
rect 160888 73788 160894 73840
rect 61378 73176 61384 73228
rect 61436 73216 61442 73228
rect 61930 73216 61936 73228
rect 61436 73188 61936 73216
rect 61436 73176 61442 73188
rect 61930 73176 61936 73188
rect 61988 73176 61994 73228
rect 194594 73176 194600 73228
rect 194652 73216 194658 73228
rect 195238 73216 195244 73228
rect 194652 73188 195244 73216
rect 194652 73176 194658 73188
rect 195238 73176 195244 73188
rect 195296 73176 195302 73228
rect 80146 73108 80152 73160
rect 80204 73148 80210 73160
rect 103514 73148 103520 73160
rect 80204 73120 103520 73148
rect 80204 73108 80210 73120
rect 103514 73108 103520 73120
rect 103572 73148 103578 73160
rect 207014 73148 207020 73160
rect 103572 73120 207020 73148
rect 103572 73108 103578 73120
rect 207014 73108 207020 73120
rect 207072 73108 207078 73160
rect 249794 73148 249800 73160
rect 238726 73120 249800 73148
rect 197354 73040 197360 73092
rect 197412 73080 197418 73092
rect 238726 73080 238754 73120
rect 249794 73108 249800 73120
rect 249852 73148 249858 73160
rect 583018 73148 583024 73160
rect 249852 73120 583024 73148
rect 249852 73108 249858 73120
rect 583018 73108 583024 73120
rect 583076 73108 583082 73160
rect 197412 73052 238754 73080
rect 197412 73040 197418 73052
rect 88334 72428 88340 72480
rect 88392 72468 88398 72480
rect 184934 72468 184940 72480
rect 88392 72440 184940 72468
rect 88392 72428 88398 72440
rect 184934 72428 184940 72440
rect 184992 72428 184998 72480
rect 207014 72428 207020 72480
rect 207072 72468 207078 72480
rect 269022 72468 269028 72480
rect 207072 72440 269028 72468
rect 207072 72428 207078 72440
rect 269022 72428 269028 72440
rect 269080 72468 269086 72480
rect 269758 72468 269764 72480
rect 269080 72440 269764 72468
rect 269080 72428 269086 72440
rect 269758 72428 269764 72440
rect 269816 72428 269822 72480
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 95326 71720 95332 71732
rect 3568 71692 95332 71720
rect 3568 71680 3574 71692
rect 95326 71680 95332 71692
rect 95384 71680 95390 71732
rect 131022 71680 131028 71732
rect 131080 71720 131086 71732
rect 226426 71720 226432 71732
rect 131080 71692 226432 71720
rect 131080 71680 131086 71692
rect 226426 71680 226432 71692
rect 226484 71680 226490 71732
rect 92474 71000 92480 71052
rect 92532 71040 92538 71052
rect 164970 71040 164976 71052
rect 92532 71012 164976 71040
rect 92532 71000 92538 71012
rect 164970 71000 164976 71012
rect 165028 71000 165034 71052
rect 192846 71000 192852 71052
rect 192904 71040 192910 71052
rect 281534 71040 281540 71052
rect 192904 71012 281540 71040
rect 192904 71000 192910 71012
rect 281534 71000 281540 71012
rect 281592 71000 281598 71052
rect 226426 70388 226432 70440
rect 226484 70428 226490 70440
rect 226978 70428 226984 70440
rect 226484 70400 226984 70428
rect 226484 70388 226490 70400
rect 226978 70388 226984 70400
rect 227036 70388 227042 70440
rect 66070 70320 66076 70372
rect 66128 70360 66134 70372
rect 185578 70360 185584 70372
rect 66128 70332 185584 70360
rect 66128 70320 66134 70332
rect 185578 70320 185584 70332
rect 185636 70320 185642 70372
rect 160738 70252 160744 70304
rect 160796 70292 160802 70304
rect 233326 70292 233332 70304
rect 160796 70264 233332 70292
rect 160796 70252 160802 70264
rect 233326 70252 233332 70264
rect 233384 70252 233390 70304
rect 94682 68960 94688 69012
rect 94740 69000 94746 69012
rect 222838 69000 222844 69012
rect 94740 68972 222844 69000
rect 94740 68960 94746 68972
rect 222838 68960 222844 68972
rect 222896 68960 222902 69012
rect 170490 68892 170496 68944
rect 170548 68932 170554 68944
rect 233878 68932 233884 68944
rect 170548 68904 233884 68932
rect 170548 68892 170554 68904
rect 233878 68892 233884 68904
rect 233936 68892 233942 68944
rect 93854 68280 93860 68332
rect 93912 68320 93918 68332
rect 106918 68320 106924 68332
rect 93912 68292 106924 68320
rect 93912 68280 93918 68292
rect 106918 68280 106924 68292
rect 106976 68280 106982 68332
rect 109034 68280 109040 68332
rect 109092 68320 109098 68332
rect 126330 68320 126336 68332
rect 109092 68292 126336 68320
rect 109092 68280 109098 68292
rect 126330 68280 126336 68292
rect 126388 68280 126394 68332
rect 235258 68280 235264 68332
rect 235316 68320 235322 68332
rect 287054 68320 287060 68332
rect 235316 68292 287060 68320
rect 235316 68280 235322 68292
rect 287054 68280 287060 68292
rect 287112 68280 287118 68332
rect 74626 67532 74632 67584
rect 74684 67572 74690 67584
rect 201494 67572 201500 67584
rect 74684 67544 201500 67572
rect 74684 67532 74690 67544
rect 201494 67532 201500 67544
rect 201552 67532 201558 67584
rect 112438 67464 112444 67516
rect 112496 67504 112502 67516
rect 230474 67504 230480 67516
rect 112496 67476 230480 67504
rect 112496 67464 112502 67476
rect 230474 67464 230480 67476
rect 230532 67464 230538 67516
rect 87046 66172 87052 66224
rect 87104 66212 87110 66224
rect 87104 66184 200114 66212
rect 87104 66172 87110 66184
rect 200086 66144 200114 66184
rect 215294 66144 215300 66156
rect 200086 66116 215300 66144
rect 215294 66104 215300 66116
rect 215352 66144 215358 66156
rect 215938 66144 215944 66156
rect 215352 66116 215944 66144
rect 215352 66104 215358 66116
rect 215938 66104 215944 66116
rect 215996 66104 216002 66156
rect 188890 65492 188896 65544
rect 188948 65532 188954 65544
rect 220078 65532 220084 65544
rect 188948 65504 220084 65532
rect 188948 65492 188954 65504
rect 220078 65492 220084 65504
rect 220136 65492 220142 65544
rect 97258 64812 97264 64864
rect 97316 64852 97322 64864
rect 241514 64852 241520 64864
rect 97316 64824 241520 64852
rect 97316 64812 97322 64824
rect 241514 64812 241520 64824
rect 241572 64812 241578 64864
rect 108390 64132 108396 64184
rect 108448 64172 108454 64184
rect 124858 64172 124864 64184
rect 108448 64144 124864 64172
rect 108448 64132 108454 64144
rect 124858 64132 124864 64144
rect 124916 64132 124922 64184
rect 202966 63520 202972 63572
rect 203024 63560 203030 63572
rect 322290 63560 322296 63572
rect 203024 63532 322296 63560
rect 203024 63520 203030 63532
rect 322290 63520 322296 63532
rect 322348 63520 322354 63572
rect 71038 63452 71044 63504
rect 71096 63492 71102 63504
rect 193858 63492 193864 63504
rect 71096 63464 193864 63492
rect 71096 63452 71102 63464
rect 193858 63452 193864 63464
rect 193916 63452 193922 63504
rect 86954 63384 86960 63436
rect 87012 63424 87018 63436
rect 121546 63424 121552 63436
rect 87012 63396 121552 63424
rect 87012 63384 87018 63396
rect 121546 63384 121552 63396
rect 121604 63384 121610 63436
rect 190362 62772 190368 62824
rect 190420 62812 190426 62824
rect 249794 62812 249800 62824
rect 190420 62784 249800 62812
rect 190420 62772 190426 62784
rect 249794 62772 249800 62784
rect 249852 62772 249858 62824
rect 215202 62500 215208 62552
rect 215260 62540 215266 62552
rect 216030 62540 216036 62552
rect 215260 62512 216036 62540
rect 215260 62500 215266 62512
rect 216030 62500 216036 62512
rect 216088 62500 216094 62552
rect 127618 62024 127624 62076
rect 127676 62064 127682 62076
rect 222194 62064 222200 62076
rect 127676 62036 222200 62064
rect 127676 62024 127682 62036
rect 222194 62024 222200 62036
rect 222252 62024 222258 62076
rect 240778 61344 240784 61396
rect 240836 61384 240842 61396
rect 269758 61384 269764 61396
rect 240836 61356 269764 61384
rect 240836 61344 240842 61356
rect 269758 61344 269764 61356
rect 269816 61344 269822 61396
rect 222194 60732 222200 60784
rect 222252 60772 222258 60784
rect 222838 60772 222844 60784
rect 222252 60744 222844 60772
rect 222252 60732 222258 60744
rect 222838 60732 222844 60744
rect 222896 60732 222902 60784
rect 89622 60664 89628 60716
rect 89680 60704 89686 60716
rect 217318 60704 217324 60716
rect 89680 60676 217324 60704
rect 89680 60664 89686 60676
rect 217318 60664 217324 60676
rect 217376 60664 217382 60716
rect 181990 59984 181996 60036
rect 182048 60024 182054 60036
rect 233878 60024 233884 60036
rect 182048 59996 233884 60024
rect 182048 59984 182054 59996
rect 233878 59984 233884 59996
rect 233936 59984 233942 60036
rect 94498 59304 94504 59356
rect 94556 59344 94562 59356
rect 213178 59344 213184 59356
rect 94556 59316 213184 59344
rect 94556 59304 94562 59316
rect 213178 59304 213184 59316
rect 213236 59304 213242 59356
rect 193950 58624 193956 58676
rect 194008 58664 194014 58676
rect 264974 58664 264980 58676
rect 194008 58636 264980 58664
rect 194008 58624 194014 58636
rect 264974 58624 264980 58636
rect 265032 58624 265038 58676
rect 77202 57876 77208 57928
rect 77260 57916 77266 57928
rect 202966 57916 202972 57928
rect 77260 57888 202972 57916
rect 77260 57876 77266 57888
rect 202966 57876 202972 57888
rect 203024 57876 203030 57928
rect 199378 57196 199384 57248
rect 199436 57236 199442 57248
rect 244274 57236 244280 57248
rect 199436 57208 244280 57236
rect 199436 57196 199442 57208
rect 244274 57196 244280 57208
rect 244332 57196 244338 57248
rect 83458 56516 83464 56568
rect 83516 56556 83522 56568
rect 210418 56556 210424 56568
rect 83516 56528 210424 56556
rect 83516 56516 83522 56528
rect 210418 56516 210424 56528
rect 210476 56516 210482 56568
rect 105538 56448 105544 56500
rect 105596 56488 105602 56500
rect 206370 56488 206376 56500
rect 105596 56460 206376 56488
rect 105596 56448 105602 56460
rect 206370 56448 206376 56460
rect 206428 56448 206434 56500
rect 46934 54476 46940 54528
rect 46992 54516 46998 54528
rect 135898 54516 135904 54528
rect 46992 54488 135904 54516
rect 46992 54476 46998 54488
rect 135898 54476 135904 54488
rect 135956 54476 135962 54528
rect 184290 54476 184296 54528
rect 184348 54516 184354 54528
rect 320266 54516 320272 54528
rect 184348 54488 320272 54516
rect 184348 54476 184354 54488
rect 320266 54476 320272 54488
rect 320324 54476 320330 54528
rect 87598 53048 87604 53100
rect 87656 53088 87662 53100
rect 140038 53088 140044 53100
rect 87656 53060 140044 53088
rect 87656 53048 87662 53060
rect 140038 53048 140044 53060
rect 140096 53048 140102 53100
rect 192938 53048 192944 53100
rect 192996 53088 193002 53100
rect 270494 53088 270500 53100
rect 192996 53060 270500 53088
rect 192996 53048 193002 53060
rect 270494 53048 270500 53060
rect 270552 53048 270558 53100
rect 75178 51756 75184 51808
rect 75236 51796 75242 51808
rect 108298 51796 108304 51808
rect 75236 51768 108304 51796
rect 75236 51756 75242 51768
rect 108298 51756 108304 51768
rect 108356 51756 108362 51808
rect 97258 51688 97264 51740
rect 97316 51728 97322 51740
rect 143534 51728 143540 51740
rect 97316 51700 143540 51728
rect 97316 51688 97322 51700
rect 143534 51688 143540 51700
rect 143592 51688 143598 51740
rect 239398 51688 239404 51740
rect 239456 51728 239462 51740
rect 259454 51728 259460 51740
rect 239456 51700 259460 51728
rect 239456 51688 239462 51700
rect 259454 51688 259460 51700
rect 259512 51688 259518 51740
rect 2866 50328 2872 50380
rect 2924 50368 2930 50380
rect 146938 50368 146944 50380
rect 2924 50340 146944 50368
rect 2924 50328 2930 50340
rect 146938 50328 146944 50340
rect 146996 50328 147002 50380
rect 202138 50328 202144 50380
rect 202196 50368 202202 50380
rect 286318 50368 286324 50380
rect 202196 50340 286324 50368
rect 202196 50328 202202 50340
rect 286318 50328 286324 50340
rect 286376 50328 286382 50380
rect 71774 48968 71780 49020
rect 71832 49008 71838 49020
rect 138658 49008 138664 49020
rect 71832 48980 138664 49008
rect 71832 48968 71838 48980
rect 138658 48968 138664 48980
rect 138716 48968 138722 49020
rect 189718 48968 189724 49020
rect 189776 49008 189782 49020
rect 580166 49008 580172 49020
rect 189776 48980 580172 49008
rect 189776 48968 189782 48980
rect 580166 48968 580172 48980
rect 580224 48968 580230 49020
rect 53834 47540 53840 47592
rect 53892 47580 53898 47592
rect 149698 47580 149704 47592
rect 53892 47552 149704 47580
rect 53892 47540 53898 47552
rect 149698 47540 149704 47552
rect 149756 47540 149762 47592
rect 187510 47540 187516 47592
rect 187568 47580 187574 47592
rect 298094 47580 298100 47592
rect 187568 47552 298100 47580
rect 187568 47540 187574 47552
rect 298094 47540 298100 47552
rect 298152 47540 298158 47592
rect 3510 46180 3516 46232
rect 3568 46220 3574 46232
rect 61378 46220 61384 46232
rect 3568 46192 61384 46220
rect 3568 46180 3574 46192
rect 61378 46180 61384 46192
rect 61436 46180 61442 46232
rect 217318 46180 217324 46232
rect 217376 46220 217382 46232
rect 291930 46220 291936 46232
rect 217376 46192 291936 46220
rect 217376 46180 217382 46192
rect 291930 46180 291936 46192
rect 291988 46180 291994 46232
rect 291838 45568 291844 45620
rect 291896 45608 291902 45620
rect 296806 45608 296812 45620
rect 291896 45580 296812 45608
rect 291896 45568 291902 45580
rect 296806 45568 296812 45580
rect 296864 45568 296870 45620
rect 64874 44820 64880 44872
rect 64932 44860 64938 44872
rect 142890 44860 142896 44872
rect 64932 44832 142896 44860
rect 64932 44820 64938 44832
rect 142890 44820 142896 44832
rect 142948 44820 142954 44872
rect 193030 44820 193036 44872
rect 193088 44860 193094 44872
rect 309134 44860 309140 44872
rect 193088 44832 309140 44860
rect 193088 44820 193094 44832
rect 309134 44820 309140 44832
rect 309192 44820 309198 44872
rect 99374 43392 99380 43444
rect 99432 43432 99438 43444
rect 141418 43432 141424 43444
rect 99432 43404 141424 43432
rect 99432 43392 99438 43404
rect 141418 43392 141424 43404
rect 141476 43392 141482 43444
rect 210418 43392 210424 43444
rect 210476 43432 210482 43444
rect 322934 43432 322940 43444
rect 210476 43404 322940 43432
rect 210476 43392 210482 43404
rect 322934 43392 322940 43404
rect 322992 43392 322998 43444
rect 66254 42032 66260 42084
rect 66312 42072 66318 42084
rect 123478 42072 123484 42084
rect 66312 42044 123484 42072
rect 66312 42032 66318 42044
rect 123478 42032 123484 42044
rect 123536 42032 123542 42084
rect 213178 40672 213184 40724
rect 213236 40712 213242 40724
rect 334066 40712 334072 40724
rect 213236 40684 334072 40712
rect 213236 40672 213242 40684
rect 334066 40672 334072 40684
rect 334124 40672 334130 40724
rect 75914 39312 75920 39364
rect 75972 39352 75978 39364
rect 155310 39352 155316 39364
rect 75972 39324 155316 39352
rect 75972 39312 75978 39324
rect 155310 39312 155316 39324
rect 155368 39312 155374 39364
rect 97994 37884 98000 37936
rect 98052 37924 98058 37936
rect 148410 37924 148416 37936
rect 98052 37896 148416 37924
rect 98052 37884 98058 37896
rect 148410 37884 148416 37896
rect 148468 37884 148474 37936
rect 204898 37204 204904 37256
rect 204956 37244 204962 37256
rect 296714 37244 296720 37256
rect 204956 37216 296720 37244
rect 204956 37204 204962 37216
rect 296714 37204 296720 37216
rect 296772 37244 296778 37256
rect 298002 37244 298008 37256
rect 296772 37216 298008 37244
rect 296772 37204 296778 37216
rect 298002 37204 298008 37216
rect 298060 37204 298066 37256
rect 45554 36524 45560 36576
rect 45612 36564 45618 36576
rect 166258 36564 166264 36576
rect 45612 36536 166264 36564
rect 45612 36524 45618 36536
rect 166258 36524 166264 36536
rect 166316 36524 166322 36576
rect 298002 36524 298008 36576
rect 298060 36564 298066 36576
rect 343634 36564 343640 36576
rect 298060 36536 343640 36564
rect 298060 36524 298066 36536
rect 343634 36524 343640 36536
rect 343692 36524 343698 36576
rect 42794 35164 42800 35216
rect 42852 35204 42858 35216
rect 170398 35204 170404 35216
rect 42852 35176 170404 35204
rect 42852 35164 42858 35176
rect 170398 35164 170404 35176
rect 170456 35164 170462 35216
rect 195238 35164 195244 35216
rect 195296 35204 195302 35216
rect 311894 35204 311900 35216
rect 195296 35176 311900 35204
rect 195296 35164 195302 35176
rect 311894 35164 311900 35176
rect 311952 35164 311958 35216
rect 23474 33736 23480 33788
rect 23532 33776 23538 33788
rect 173158 33776 173164 33788
rect 23532 33748 173164 33776
rect 23532 33736 23538 33748
rect 173158 33736 173164 33748
rect 173216 33736 173222 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 57238 33096 57244 33108
rect 3568 33068 57244 33096
rect 3568 33056 3574 33068
rect 57238 33056 57244 33068
rect 57296 33056 57302 33108
rect 117314 32444 117320 32496
rect 117372 32484 117378 32496
rect 156598 32484 156604 32496
rect 117372 32456 156604 32484
rect 117372 32444 117378 32456
rect 156598 32444 156604 32456
rect 156656 32444 156662 32496
rect 55214 32376 55220 32428
rect 55272 32416 55278 32428
rect 134610 32416 134616 32428
rect 55272 32388 134616 32416
rect 55272 32376 55278 32388
rect 134610 32376 134616 32388
rect 134668 32376 134674 32428
rect 208394 32376 208400 32428
rect 208452 32416 208458 32428
rect 278774 32416 278780 32428
rect 208452 32388 278780 32416
rect 208452 32376 208458 32388
rect 278774 32376 278780 32388
rect 278832 32376 278838 32428
rect 113174 31016 113180 31068
rect 113232 31056 113238 31068
rect 157978 31056 157984 31068
rect 113232 31028 157984 31056
rect 113232 31016 113238 31028
rect 157978 31016 157984 31028
rect 158036 31016 158042 31068
rect 215938 31016 215944 31068
rect 215996 31056 216002 31068
rect 266354 31056 266360 31068
rect 215996 31028 266360 31056
rect 215996 31016 216002 31028
rect 266354 31016 266360 31028
rect 266412 31016 266418 31068
rect 81434 29588 81440 29640
rect 81492 29628 81498 29640
rect 179414 29628 179420 29640
rect 81492 29600 179420 29628
rect 81492 29588 81498 29600
rect 179414 29588 179420 29600
rect 179472 29588 179478 29640
rect 183370 29588 183376 29640
rect 183428 29628 183434 29640
rect 263686 29628 263692 29640
rect 183428 29600 263692 29628
rect 183428 29588 183434 29600
rect 263686 29588 263692 29600
rect 263744 29588 263750 29640
rect 67634 28228 67640 28280
rect 67692 28268 67698 28280
rect 171134 28268 171140 28280
rect 67692 28240 171140 28268
rect 67692 28228 67698 28240
rect 171134 28228 171140 28240
rect 171192 28228 171198 28280
rect 226978 28228 226984 28280
rect 227036 28268 227042 28280
rect 277394 28268 277400 28280
rect 227036 28240 277400 28268
rect 227036 28228 227042 28240
rect 277394 28228 277400 28240
rect 277452 28228 277458 28280
rect 82814 26868 82820 26920
rect 82872 26908 82878 26920
rect 151078 26908 151084 26920
rect 82872 26880 151084 26908
rect 82872 26868 82878 26880
rect 151078 26868 151084 26880
rect 151136 26868 151142 26920
rect 193858 25508 193864 25560
rect 193916 25548 193922 25560
rect 291194 25548 291200 25560
rect 193916 25520 291200 25548
rect 193916 25508 193922 25520
rect 291194 25508 291200 25520
rect 291252 25508 291258 25560
rect 96614 24148 96620 24200
rect 96672 24188 96678 24200
rect 130470 24188 130476 24200
rect 96672 24160 130476 24188
rect 96672 24148 96678 24160
rect 130470 24148 130476 24160
rect 130528 24148 130534 24200
rect 59354 24080 59360 24132
rect 59412 24120 59418 24132
rect 131758 24120 131764 24132
rect 59412 24092 131764 24120
rect 59412 24080 59418 24092
rect 131758 24080 131764 24092
rect 131816 24080 131822 24132
rect 78674 22720 78680 22772
rect 78732 22760 78738 22772
rect 145558 22760 145564 22772
rect 78732 22732 145564 22760
rect 78732 22720 78738 22732
rect 145558 22720 145564 22732
rect 145616 22720 145622 22772
rect 57974 21360 57980 21412
rect 58032 21400 58038 21412
rect 137370 21400 137376 21412
rect 58032 21372 137376 21400
rect 58032 21360 58038 21372
rect 137370 21360 137376 21372
rect 137428 21360 137434 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 90358 20652 90364 20664
rect 3476 20624 90364 20652
rect 3476 20612 3482 20624
rect 90358 20612 90364 20624
rect 90416 20612 90422 20664
rect 95234 19932 95240 19984
rect 95292 19972 95298 19984
rect 162854 19972 162860 19984
rect 95292 19944 162860 19972
rect 95292 19932 95298 19944
rect 162854 19932 162860 19944
rect 162912 19932 162918 19984
rect 205542 19932 205548 19984
rect 205600 19972 205606 19984
rect 288434 19972 288440 19984
rect 205600 19944 288440 19972
rect 205600 19932 205606 19944
rect 288434 19932 288440 19944
rect 288492 19932 288498 19984
rect 63494 18572 63500 18624
rect 63552 18612 63558 18624
rect 178678 18612 178684 18624
rect 63552 18584 178684 18612
rect 63552 18572 63558 18584
rect 178678 18572 178684 18584
rect 178736 18572 178742 18624
rect 215202 18572 215208 18624
rect 215260 18612 215266 18624
rect 284386 18612 284392 18624
rect 215260 18584 284392 18612
rect 215260 18572 215266 18584
rect 284386 18572 284392 18584
rect 284444 18572 284450 18624
rect 322198 18572 322204 18624
rect 322256 18612 322262 18624
rect 332594 18612 332600 18624
rect 322256 18584 332600 18612
rect 322256 18572 322262 18584
rect 332594 18572 332600 18584
rect 332652 18572 332658 18624
rect 309778 17960 309784 18012
rect 309836 18000 309842 18012
rect 316126 18000 316132 18012
rect 309836 17972 316132 18000
rect 309836 17960 309842 17972
rect 316126 17960 316132 17972
rect 316184 17960 316190 18012
rect 233878 17280 233884 17332
rect 233936 17320 233942 17332
rect 251266 17320 251272 17332
rect 233936 17292 251272 17320
rect 233936 17280 233942 17292
rect 251266 17280 251272 17292
rect 251324 17280 251330 17332
rect 49694 17212 49700 17264
rect 49752 17252 49758 17264
rect 162118 17252 162124 17264
rect 49752 17224 162124 17252
rect 49752 17212 49758 17224
rect 162118 17212 162124 17224
rect 162176 17212 162182 17264
rect 206278 17212 206284 17264
rect 206336 17252 206342 17264
rect 233970 17252 233976 17264
rect 206336 17224 233976 17252
rect 206336 17212 206342 17224
rect 233970 17212 233976 17224
rect 234028 17212 234034 17264
rect 260098 17212 260104 17264
rect 260156 17252 260162 17264
rect 336734 17252 336740 17264
rect 260156 17224 336740 17252
rect 260156 17212 260162 17224
rect 336734 17212 336740 17224
rect 336792 17212 336798 17264
rect 91554 15852 91560 15904
rect 91612 15892 91618 15904
rect 129090 15892 129096 15904
rect 91612 15864 129096 15892
rect 91612 15852 91618 15864
rect 129090 15852 129096 15864
rect 129148 15852 129154 15904
rect 245010 15852 245016 15904
rect 245068 15892 245074 15904
rect 256694 15892 256700 15904
rect 245068 15864 256700 15892
rect 245068 15852 245074 15864
rect 256694 15852 256700 15864
rect 256752 15852 256758 15904
rect 302878 15852 302884 15904
rect 302936 15892 302942 15904
rect 314654 15892 314660 15904
rect 302936 15864 314660 15892
rect 302936 15852 302942 15864
rect 314654 15852 314660 15864
rect 314712 15852 314718 15904
rect 106 14492 112 14544
rect 164 14532 170 14544
rect 96706 14532 96712 14544
rect 164 14504 96712 14532
rect 164 14492 170 14504
rect 96706 14492 96712 14504
rect 96764 14492 96770 14544
rect 222838 14492 222844 14544
rect 222896 14532 222902 14544
rect 302878 14532 302884 14544
rect 222896 14504 302884 14532
rect 222896 14492 222902 14504
rect 302878 14492 302884 14504
rect 302936 14492 302942 14544
rect 87506 14424 87512 14476
rect 87564 14464 87570 14476
rect 231118 14464 231124 14476
rect 87564 14436 231124 14464
rect 87564 14424 87570 14436
rect 231118 14424 231124 14436
rect 231176 14424 231182 14476
rect 89898 13064 89904 13116
rect 89956 13104 89962 13116
rect 155218 13104 155224 13116
rect 89956 13076 155224 13104
rect 89956 13064 89962 13076
rect 155218 13064 155224 13076
rect 155276 13064 155282 13116
rect 200758 13064 200764 13116
rect 200816 13104 200822 13116
rect 340966 13104 340972 13116
rect 200816 13076 340972 13104
rect 200816 13064 200822 13076
rect 340966 13064 340972 13076
rect 341024 13064 341030 13116
rect 61562 11704 61568 11756
rect 61620 11744 61626 11756
rect 133138 11744 133144 11756
rect 61620 11716 133144 11744
rect 61620 11704 61626 11716
rect 133138 11704 133144 11716
rect 133196 11704 133202 11756
rect 188982 11704 188988 11756
rect 189040 11744 189046 11756
rect 280706 11744 280712 11756
rect 189040 11716 280712 11744
rect 189040 11704 189046 11716
rect 280706 11704 280712 11716
rect 280764 11704 280770 11756
rect 324406 11704 324412 11756
rect 324464 11744 324470 11756
rect 325602 11744 325608 11756
rect 324464 11716 325608 11744
rect 324464 11704 324470 11716
rect 325602 11704 325608 11716
rect 325660 11704 325666 11756
rect 108114 10412 108120 10464
rect 108172 10452 108178 10464
rect 142798 10452 142804 10464
rect 108172 10424 142804 10452
rect 108172 10412 108178 10424
rect 142798 10412 142804 10424
rect 142856 10412 142862 10464
rect 73338 10344 73344 10396
rect 73396 10384 73402 10396
rect 108390 10384 108396 10396
rect 73396 10356 108396 10384
rect 73396 10344 73402 10356
rect 108390 10344 108396 10356
rect 108448 10344 108454 10396
rect 86402 10276 86408 10328
rect 86460 10316 86466 10328
rect 126238 10316 126244 10328
rect 86460 10288 126244 10316
rect 86460 10276 86466 10288
rect 126238 10276 126244 10288
rect 126296 10276 126302 10328
rect 197998 10276 198004 10328
rect 198056 10316 198062 10328
rect 342898 10316 342904 10328
rect 198056 10288 342904 10316
rect 198056 10276 198062 10288
rect 342898 10276 342904 10288
rect 342956 10276 342962 10328
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 87598 9024 87604 9036
rect 1728 8996 87604 9024
rect 1728 8984 1734 8996
rect 87598 8984 87604 8996
rect 87656 8984 87662 9036
rect 78582 8916 78588 8968
rect 78640 8956 78646 8968
rect 168374 8956 168380 8968
rect 78640 8928 168380 8956
rect 78640 8916 78646 8928
rect 168374 8916 168380 8928
rect 168432 8916 168438 8968
rect 196618 8916 196624 8968
rect 196676 8956 196682 8968
rect 258258 8956 258264 8968
rect 196676 8928 258264 8956
rect 196676 8916 196682 8928
rect 258258 8916 258264 8928
rect 258316 8916 258322 8968
rect 258718 8236 258724 8288
rect 258776 8276 258782 8288
rect 261754 8276 261760 8288
rect 258776 8248 261760 8276
rect 258776 8236 258782 8248
rect 261754 8236 261760 8248
rect 261812 8236 261818 8288
rect 111610 7624 111616 7676
rect 111668 7664 111674 7676
rect 148318 7664 148324 7676
rect 111668 7636 148324 7664
rect 111668 7624 111674 7636
rect 148318 7624 148324 7636
rect 148376 7624 148382 7676
rect 67726 7556 67732 7608
rect 67784 7596 67790 7608
rect 125870 7596 125876 7608
rect 67784 7568 125876 7596
rect 67784 7556 67790 7568
rect 125870 7556 125876 7568
rect 125928 7556 125934 7608
rect 224862 7556 224868 7608
rect 224920 7596 224926 7608
rect 254670 7596 254676 7608
rect 224920 7568 254676 7596
rect 224920 7556 224926 7568
rect 254670 7556 254676 7568
rect 254728 7556 254734 7608
rect 280798 7556 280804 7608
rect 280856 7596 280862 7608
rect 330386 7596 330392 7608
rect 280856 7568 330392 7596
rect 280856 7556 280862 7568
rect 330386 7556 330392 7568
rect 330444 7556 330450 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 7558 6848 7564 6860
rect 3476 6820 7564 6848
rect 3476 6808 3482 6820
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 80882 6128 80888 6180
rect 80940 6168 80946 6180
rect 130378 6168 130384 6180
rect 80940 6140 130384 6168
rect 80940 6128 80946 6140
rect 130378 6128 130384 6140
rect 130436 6128 130442 6180
rect 206370 6128 206376 6180
rect 206428 6168 206434 6180
rect 247586 6168 247592 6180
rect 206428 6140 247592 6168
rect 206428 6128 206434 6140
rect 247586 6128 247592 6140
rect 247644 6128 247650 6180
rect 286318 6128 286324 6180
rect 286376 6168 286382 6180
rect 329190 6168 329196 6180
rect 286376 6140 329196 6168
rect 286376 6128 286382 6140
rect 329190 6128 329196 6140
rect 329248 6128 329254 6180
rect 134518 5516 134524 5568
rect 134576 5556 134582 5568
rect 136450 5556 136456 5568
rect 134576 5528 136456 5556
rect 134576 5516 134582 5528
rect 136450 5516 136456 5528
rect 136508 5516 136514 5568
rect 305638 5516 305644 5568
rect 305696 5556 305702 5568
rect 309042 5556 309048 5568
rect 305696 5528 309048 5556
rect 305696 5516 305702 5528
rect 309042 5516 309048 5528
rect 309100 5516 309106 5568
rect 346946 5516 346952 5568
rect 347004 5556 347010 5568
rect 349154 5556 349160 5568
rect 347004 5528 349160 5556
rect 347004 5516 347010 5528
rect 349154 5516 349160 5528
rect 349212 5516 349218 5568
rect 69106 4768 69112 4820
rect 69164 4808 69170 4820
rect 152550 4808 152556 4820
rect 69164 4780 152556 4808
rect 69164 4768 69170 4780
rect 152550 4768 152556 4780
rect 152608 4768 152614 4820
rect 220078 4768 220084 4820
rect 220136 4808 220142 4820
rect 244090 4808 244096 4820
rect 220136 4780 244096 4808
rect 220136 4768 220142 4780
rect 244090 4768 244096 4780
rect 244148 4768 244154 4820
rect 238018 4360 238024 4412
rect 238076 4400 238082 4412
rect 239306 4400 239312 4412
rect 238076 4372 239312 4400
rect 238076 4360 238082 4372
rect 239306 4360 239312 4372
rect 239364 4360 239370 4412
rect 276014 4360 276020 4412
rect 276072 4400 276078 4412
rect 278038 4400 278044 4412
rect 276072 4372 278044 4400
rect 276072 4360 276078 4372
rect 278038 4360 278044 4372
rect 278096 4360 278102 4412
rect 228358 4088 228364 4140
rect 228416 4128 228422 4140
rect 248782 4128 248788 4140
rect 228416 4100 248788 4128
rect 228416 4088 228422 4100
rect 248782 4088 248788 4100
rect 248840 4128 248846 4140
rect 249058 4128 249064 4140
rect 248840 4100 249064 4128
rect 248840 4088 248846 4100
rect 249058 4088 249064 4100
rect 249116 4088 249122 4140
rect 266998 4088 267004 4140
rect 267056 4128 267062 4140
rect 267734 4128 267740 4140
rect 267056 4100 267740 4128
rect 267056 4088 267062 4100
rect 267734 4088 267740 4100
rect 267792 4088 267798 4140
rect 302970 3952 302976 4004
rect 303028 3992 303034 4004
rect 306742 3992 306748 4004
rect 303028 3964 306748 3992
rect 303028 3952 303034 3964
rect 306742 3952 306748 3964
rect 306800 3952 306806 4004
rect 323578 3952 323584 4004
rect 323636 3992 323642 4004
rect 326798 3992 326804 4004
rect 323636 3964 326804 3992
rect 323636 3952 323642 3964
rect 326798 3952 326804 3964
rect 326856 3952 326862 4004
rect 150618 3612 150624 3664
rect 150676 3652 150682 3664
rect 152458 3652 152464 3664
rect 150676 3624 152464 3652
rect 150676 3612 150682 3624
rect 152458 3612 152464 3624
rect 152516 3612 152522 3664
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 252370 3584 252376 3596
rect 251232 3556 252376 3584
rect 251232 3544 251238 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 316126 3544 316132 3596
rect 316184 3584 316190 3596
rect 317322 3584 317328 3596
rect 316184 3556 317328 3584
rect 316184 3544 316190 3556
rect 317322 3544 317328 3556
rect 317380 3544 317386 3596
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 4062 3516 4068 3528
rect 2832 3488 4068 3516
rect 2832 3476 2838 3488
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 22738 3516 22744 3528
rect 19484 3488 22744 3516
rect 19484 3476 19490 3488
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 37182 3516 37188 3528
rect 35952 3488 37188 3516
rect 35952 3476 35958 3488
rect 37182 3476 37188 3488
rect 37240 3476 37246 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 98638 3516 98644 3528
rect 84528 3488 98644 3516
rect 84528 3476 84534 3488
rect 98638 3476 98644 3488
rect 98696 3476 98702 3528
rect 101398 3476 101404 3528
rect 101456 3516 101462 3528
rect 102226 3516 102232 3528
rect 101456 3488 102232 3516
rect 101456 3476 101462 3488
rect 102226 3476 102232 3488
rect 102284 3476 102290 3528
rect 118694 3476 118700 3528
rect 118752 3516 118758 3528
rect 119890 3516 119896 3528
rect 118752 3488 119896 3516
rect 118752 3476 118758 3488
rect 119890 3476 119896 3488
rect 119948 3476 119954 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144730 3516 144736 3528
rect 143592 3488 144736 3516
rect 143592 3476 143598 3488
rect 144730 3476 144736 3488
rect 144788 3476 144794 3528
rect 270034 3476 270040 3528
rect 270092 3516 270098 3528
rect 270586 3516 270592 3528
rect 270092 3488 270592 3516
rect 270092 3476 270098 3488
rect 270586 3476 270592 3488
rect 270644 3476 270650 3528
rect 289078 3476 289084 3528
rect 289136 3516 289142 3528
rect 290182 3516 290188 3528
rect 289136 3488 290188 3516
rect 289136 3476 289142 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 291930 3476 291936 3528
rect 291988 3516 291994 3528
rect 294874 3516 294880 3528
rect 291988 3488 294880 3516
rect 291988 3476 291994 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 298738 3476 298744 3528
rect 298796 3516 298802 3528
rect 305546 3516 305552 3528
rect 298796 3488 305552 3516
rect 298796 3476 298802 3488
rect 305546 3476 305552 3488
rect 305604 3476 305610 3528
rect 307018 3476 307024 3528
rect 307076 3516 307082 3528
rect 311434 3516 311440 3528
rect 307076 3488 311440 3516
rect 307076 3476 307082 3488
rect 311434 3476 311440 3488
rect 311492 3476 311498 3528
rect 319714 3476 319720 3528
rect 319772 3516 319778 3528
rect 320174 3516 320180 3528
rect 319772 3488 320180 3516
rect 319772 3476 319778 3488
rect 320174 3476 320180 3488
rect 320232 3476 320238 3528
rect 351638 3476 351644 3528
rect 351696 3516 351702 3528
rect 353294 3516 353300 3528
rect 351696 3488 353300 3516
rect 351696 3476 351702 3488
rect 353294 3476 353300 3488
rect 353352 3476 353358 3528
rect 63218 3408 63224 3460
rect 63276 3448 63282 3460
rect 75178 3448 75184 3460
rect 63276 3420 75184 3448
rect 63276 3408 63282 3420
rect 75178 3408 75184 3420
rect 75236 3408 75242 3460
rect 77386 3408 77392 3460
rect 77444 3448 77450 3460
rect 104250 3448 104256 3460
rect 77444 3420 104256 3448
rect 77444 3408 77450 3420
rect 104250 3408 104256 3420
rect 104308 3408 104314 3460
rect 140038 3408 140044 3460
rect 140096 3448 140102 3460
rect 184198 3448 184204 3460
rect 140096 3420 184204 3448
rect 140096 3408 140102 3420
rect 184198 3408 184204 3420
rect 184256 3408 184262 3460
rect 233970 3408 233976 3460
rect 234028 3448 234034 3460
rect 242894 3448 242900 3460
rect 234028 3420 242900 3448
rect 234028 3408 234034 3420
rect 242894 3408 242900 3420
rect 242952 3408 242958 3460
rect 276750 3408 276756 3460
rect 276808 3448 276814 3460
rect 286594 3448 286600 3460
rect 276808 3420 286600 3448
rect 276808 3408 276814 3420
rect 286594 3408 286600 3420
rect 286652 3408 286658 3460
rect 580994 3272 581000 3324
rect 581052 3312 581058 3324
rect 582558 3312 582564 3324
rect 581052 3284 582564 3312
rect 581052 3272 581058 3284
rect 582558 3272 582564 3284
rect 582616 3272 582622 3324
rect 318150 3204 318156 3256
rect 318208 3244 318214 3256
rect 322106 3244 322112 3256
rect 318208 3216 322112 3244
rect 318208 3204 318214 3216
rect 322106 3204 322112 3216
rect 322164 3204 322170 3256
rect 348050 3204 348056 3256
rect 348108 3244 348114 3256
rect 351914 3244 351920 3256
rect 348108 3216 351920 3244
rect 348108 3204 348114 3216
rect 351914 3204 351920 3216
rect 351972 3204 351978 3256
rect 260650 3136 260656 3188
rect 260708 3176 260714 3188
rect 263594 3176 263600 3188
rect 260708 3148 263600 3176
rect 260708 3136 260714 3148
rect 263594 3136 263600 3148
rect 263652 3136 263658 3188
rect 269758 3136 269764 3188
rect 269816 3176 269822 3188
rect 272426 3176 272432 3188
rect 269816 3148 272432 3176
rect 269816 3136 269822 3148
rect 272426 3136 272432 3148
rect 272484 3136 272490 3188
rect 322290 3136 322296 3188
rect 322348 3176 322354 3188
rect 324406 3176 324412 3188
rect 322348 3148 324412 3176
rect 322348 3136 322354 3148
rect 324406 3136 324412 3148
rect 324464 3136 324470 3188
rect 345658 3136 345664 3188
rect 345716 3176 345722 3188
rect 349246 3176 349252 3188
rect 345716 3148 349252 3176
rect 345716 3136 345722 3148
rect 349246 3136 349252 3148
rect 349304 3136 349310 3188
rect 287698 3000 287704 3052
rect 287756 3040 287762 3052
rect 292574 3040 292580 3052
rect 287756 3012 292580 3040
rect 287756 3000 287762 3012
rect 292574 3000 292580 3012
rect 292632 3000 292638 3052
rect 282178 2932 282184 2984
rect 282236 2972 282242 2984
rect 283098 2972 283104 2984
rect 282236 2944 283104 2972
rect 282236 2932 282242 2944
rect 283098 2932 283104 2944
rect 283156 2932 283162 2984
rect 299474 2592 299480 2644
rect 299532 2632 299538 2644
rect 300762 2632 300768 2644
rect 299532 2604 300768 2632
rect 299532 2592 299538 2604
rect 300762 2592 300768 2604
rect 300820 2592 300826 2644
rect 93946 2116 93952 2168
rect 94004 2156 94010 2168
rect 137278 2156 137284 2168
rect 94004 2128 137284 2156
rect 94004 2116 94010 2128
rect 137278 2116 137284 2128
rect 137336 2116 137342 2168
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 33778 2088 33784 2100
rect 7708 2060 33784 2088
rect 7708 2048 7714 2060
rect 33778 2048 33784 2060
rect 33836 2048 33842 2100
rect 51350 2048 51356 2100
rect 51408 2088 51414 2100
rect 97258 2088 97264 2100
rect 51408 2060 97264 2088
rect 51408 2048 51414 2060
rect 97258 2048 97264 2060
rect 97316 2048 97322 2100
<< via1 >>
rect 242808 703128 242860 703180
rect 348792 703128 348844 703180
rect 274548 703060 274600 703112
rect 413652 703060 413704 703112
rect 184296 702992 184348 703044
rect 332508 702992 332560 703044
rect 201500 702924 201552 702976
rect 202788 702924 202840 702976
rect 280804 702924 280856 702976
rect 429844 702924 429896 702976
rect 188896 702856 188948 702908
rect 364984 702856 365036 702908
rect 218980 702788 219032 702840
rect 269304 702788 269356 702840
rect 285588 702788 285640 702840
rect 462320 702788 462372 702840
rect 169760 702720 169812 702772
rect 170312 702720 170364 702772
rect 224224 702720 224276 702772
rect 248420 702720 248472 702772
rect 494796 702720 494848 702772
rect 206284 702652 206336 702704
rect 397368 702652 397420 702704
rect 24308 702584 24360 702636
rect 85580 702584 85632 702636
rect 137836 702584 137888 702636
rect 215300 702584 215352 702636
rect 222844 702584 222896 702636
rect 478512 702584 478564 702636
rect 8116 702516 8168 702568
rect 96620 702516 96672 702568
rect 154120 702516 154172 702568
rect 233240 702516 233292 702568
rect 271144 702516 271196 702568
rect 527180 702516 527232 702568
rect 67640 702448 67692 702500
rect 169760 702448 169812 702500
rect 180064 702448 180116 702500
rect 235172 702448 235224 702500
rect 255964 702448 256016 702500
rect 543464 702448 543516 702500
rect 62028 700340 62080 700392
rect 72976 700340 73028 700392
rect 84108 700340 84160 700392
rect 89168 700340 89220 700392
rect 71688 700272 71740 700324
rect 105452 700272 105504 700324
rect 251824 700272 251876 700324
rect 283840 700272 283892 700324
rect 559656 700272 559708 700324
rect 582840 700272 582892 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 3424 683136 3476 683188
rect 33784 683136 33836 683188
rect 3516 670692 3568 670744
rect 15844 670692 15896 670744
rect 3424 656888 3476 656940
rect 36544 656888 36596 656940
rect 144828 622412 144880 622464
rect 241520 622412 241572 622464
rect 151728 619624 151780 619676
rect 251180 619624 251232 619676
rect 251824 619624 251876 619676
rect 205640 619556 205692 619608
rect 206284 619556 206336 619608
rect 3516 618604 3568 618656
rect 7564 618604 7616 618656
rect 178776 618332 178828 618384
rect 236000 618332 236052 618384
rect 129648 618264 129700 618316
rect 205640 618264 205692 618316
rect 177488 616904 177540 616956
rect 242900 616904 242952 616956
rect 141976 616836 142028 616888
rect 219440 616836 219492 616888
rect 233240 615952 233292 616004
rect 233884 615952 233936 616004
rect 184848 615544 184900 615596
rect 233240 615544 233292 615596
rect 142068 615476 142120 615528
rect 213920 615476 213972 615528
rect 140688 614184 140740 614236
rect 207664 614184 207716 614236
rect 152556 614116 152608 614168
rect 232320 614116 232372 614168
rect 153844 612824 153896 612876
rect 221648 612824 221700 612876
rect 71780 612756 71832 612808
rect 258080 612756 258132 612808
rect 188988 611396 189040 611448
rect 230480 611396 230532 611448
rect 67548 611328 67600 611380
rect 254032 611328 254084 611380
rect 187516 610036 187568 610088
rect 217232 610036 217284 610088
rect 123484 609968 123536 610020
rect 256700 609968 256752 610020
rect 201500 609220 201552 609272
rect 222292 609220 222344 609272
rect 182088 608676 182140 608728
rect 226340 608676 226392 608728
rect 139308 608608 139360 608660
rect 200672 608608 200724 608660
rect 188344 607248 188396 607300
rect 196716 607248 196768 607300
rect 177396 607180 177448 607232
rect 209412 607180 209464 607232
rect 215668 606432 215720 606484
rect 582380 606432 582432 606484
rect 184388 605888 184440 605940
rect 215668 605888 215720 605940
rect 3516 605820 3568 605872
rect 94688 605820 94740 605872
rect 98644 605820 98696 605872
rect 144736 605820 144788 605872
rect 180708 605820 180760 605872
rect 214380 605820 214432 605872
rect 183468 604528 183520 604580
rect 206100 604528 206152 604580
rect 169024 604460 169076 604512
rect 216956 604460 217008 604512
rect 241796 604460 241848 604512
rect 242808 604460 242860 604512
rect 274824 604460 274876 604512
rect 289728 604460 289780 604512
rect 582840 604460 582892 604512
rect 246212 603168 246264 603220
rect 254584 603168 254636 603220
rect 177304 603100 177356 603152
rect 203708 603100 203760 603152
rect 241060 603100 241112 603152
rect 281540 603100 281592 603152
rect 222200 602148 222252 602200
rect 223028 602148 223080 602200
rect 191748 601740 191800 601792
rect 263692 601740 263744 601792
rect 104164 601672 104216 601724
rect 211252 601672 211304 601724
rect 252468 601672 252520 601724
rect 259460 601672 259512 601724
rect 224224 601604 224276 601656
rect 225236 601604 225288 601656
rect 233884 601536 233936 601588
rect 235356 601536 235408 601588
rect 192576 600380 192628 600432
rect 204260 600380 204312 600432
rect 239772 600380 239824 600432
rect 271880 600380 271932 600432
rect 148968 600312 149020 600364
rect 200396 600312 200448 600364
rect 216680 600312 216732 600364
rect 227812 600312 227864 600364
rect 251180 600312 251232 600364
rect 299480 600312 299532 600364
rect 180156 599020 180208 599072
rect 192484 599156 192536 599208
rect 197636 599156 197688 599208
rect 193404 599088 193456 599140
rect 66076 598952 66128 599004
rect 187608 598952 187660 599004
rect 192668 598952 192720 599004
rect 195612 598952 195664 599004
rect 229008 599020 229060 599072
rect 247684 599020 247736 599072
rect 257344 599020 257396 599072
rect 205180 598952 205232 599004
rect 222936 598952 222988 599004
rect 280160 598952 280212 599004
rect 192944 598884 192996 598936
rect 195060 598884 195112 598936
rect 197360 598884 197412 598936
rect 245200 598884 245252 598936
rect 256056 598884 256108 598936
rect 193312 598816 193364 598868
rect 246764 598408 246816 598460
rect 112444 597592 112496 597644
rect 189724 597592 189776 597644
rect 161388 597524 161440 597576
rect 192944 597524 192996 597576
rect 255412 597592 255464 597644
rect 287060 597592 287112 597644
rect 273352 597524 273404 597576
rect 150440 596776 150492 596828
rect 184388 596776 184440 596828
rect 253388 596776 253440 596828
rect 293960 596776 294012 596828
rect 86960 596164 87012 596216
rect 150440 596164 150492 596216
rect 255412 596164 255464 596216
rect 267740 596164 267792 596216
rect 92480 595416 92532 595468
rect 165528 595416 165580 595468
rect 165528 594872 165580 594924
rect 166264 594872 166316 594924
rect 170404 594872 170456 594924
rect 190644 594872 190696 594924
rect 159364 594804 159416 594856
rect 191748 594804 191800 594856
rect 175188 594124 175240 594176
rect 192760 594124 192812 594176
rect 143356 594056 143408 594108
rect 192668 594056 192720 594108
rect 255320 594056 255372 594108
rect 285680 594056 285732 594108
rect 69848 593376 69900 593428
rect 143356 593376 143408 593428
rect 285680 593376 285732 593428
rect 582656 593376 582708 593428
rect 175096 592628 175148 592680
rect 192576 592628 192628 592680
rect 256332 592628 256384 592680
rect 256700 592628 256752 592680
rect 284300 592628 284352 592680
rect 299572 592628 299624 592680
rect 164884 592084 164936 592136
rect 191748 592084 191800 592136
rect 89720 592016 89772 592068
rect 175096 592016 175148 592068
rect 95148 591268 95200 591320
rect 192484 591268 192536 591320
rect 253480 591268 253532 591320
rect 298100 591268 298152 591320
rect 163504 590656 163556 590708
rect 191012 590656 191064 590708
rect 255412 590656 255464 590708
rect 265072 590656 265124 590708
rect 77392 589976 77444 590028
rect 84108 589976 84160 590028
rect 122840 589976 122892 590028
rect 36544 589908 36596 589960
rect 74632 589908 74684 589960
rect 116584 589908 116636 589960
rect 190552 589908 190604 589960
rect 254584 589908 254636 589960
rect 292580 589908 292632 589960
rect 255412 589296 255464 589348
rect 261024 589296 261076 589348
rect 40040 589228 40092 589280
rect 95148 589228 95200 589280
rect 133788 588548 133840 588600
rect 177396 588548 177448 588600
rect 85488 587868 85540 587920
rect 133788 587868 133840 587920
rect 255412 587868 255464 587920
rect 287152 587868 287204 587920
rect 81808 587120 81860 587172
rect 186964 587120 187016 587172
rect 256056 587120 256108 587172
rect 270500 587120 270552 587172
rect 150348 586508 150400 586560
rect 191196 586576 191248 586628
rect 187056 586508 187108 586560
rect 190460 586508 190512 586560
rect 71688 585760 71740 585812
rect 106924 585760 106976 585812
rect 67364 585148 67416 585200
rect 71688 585148 71740 585200
rect 92112 585148 92164 585200
rect 118700 585148 118752 585200
rect 168288 585148 168340 585200
rect 191748 585148 191800 585200
rect 255320 584400 255372 584452
rect 258080 584400 258132 584452
rect 277492 584400 277544 584452
rect 582380 584400 582432 584452
rect 73528 583788 73580 583840
rect 111064 583788 111116 583840
rect 157156 583788 157208 583840
rect 191748 583788 191800 583840
rect 79048 583720 79100 583772
rect 158720 583720 158772 583772
rect 255412 583652 255464 583704
rect 274548 583652 274600 583704
rect 88248 583380 88300 583432
rect 88984 583380 89036 583432
rect 94412 583380 94464 583432
rect 98644 583380 98696 583432
rect 148692 582972 148744 583024
rect 191288 582972 191340 583024
rect 274548 582972 274600 583024
rect 284392 582972 284444 583024
rect 77208 582768 77260 582820
rect 79324 582768 79376 582820
rect 76288 582428 76340 582480
rect 95148 582428 95200 582480
rect 93768 582360 93820 582412
rect 177396 582360 177448 582412
rect 182824 582360 182876 582412
rect 191748 582360 191800 582412
rect 158536 581612 158588 581664
rect 177488 581612 177540 581664
rect 67456 581068 67508 581120
rect 124864 581068 124916 581120
rect 3332 580932 3384 580984
rect 80244 581000 80296 581052
rect 176568 581000 176620 581052
rect 191748 581000 191800 581052
rect 69020 580660 69072 580712
rect 86592 580660 86644 580712
rect 91008 580660 91060 580712
rect 98644 580660 98696 580712
rect 63408 579708 63460 579760
rect 66628 579708 66680 579760
rect 53748 579640 53800 579692
rect 255964 580252 256016 580304
rect 278780 580252 278832 580304
rect 161480 579708 161532 579760
rect 188344 579708 188396 579760
rect 98644 579640 98696 579692
rect 169760 579640 169812 579692
rect 95148 578892 95200 578944
rect 108304 578892 108356 578944
rect 158720 578892 158772 578944
rect 159916 578892 159968 578944
rect 184296 578892 184348 578944
rect 55128 578212 55180 578264
rect 66444 578212 66496 578264
rect 96804 578212 96856 578264
rect 134524 578212 134576 578264
rect 186964 578212 187016 578264
rect 191564 578212 191616 578264
rect 98552 578144 98604 578196
rect 191748 578144 191800 578196
rect 137928 577464 137980 577516
rect 187056 577464 187108 577516
rect 255412 577464 255464 577516
rect 298192 577464 298244 577516
rect 255412 576852 255464 576904
rect 264980 576852 265032 576904
rect 3424 576784 3476 576836
rect 67548 576784 67600 576836
rect 97908 576784 97960 576836
rect 123484 576784 123536 576836
rect 94688 576036 94740 576088
rect 96712 576036 96764 576088
rect 181904 575560 181956 575612
rect 191012 575560 191064 575612
rect 67548 575492 67600 575544
rect 67824 575492 67876 575544
rect 119436 575492 119488 575544
rect 191196 575492 191248 575544
rect 255412 575492 255464 575544
rect 270592 575492 270644 575544
rect 172428 574744 172480 574796
rect 185584 574744 185636 574796
rect 96804 574064 96856 574116
rect 151084 574064 151136 574116
rect 166356 574064 166408 574116
rect 191288 574064 191340 574116
rect 255412 574064 255464 574116
rect 273444 574064 273496 574116
rect 98000 573316 98052 573368
rect 137100 573316 137152 573368
rect 163596 572772 163648 572824
rect 191012 572772 191064 572824
rect 64604 572704 64656 572756
rect 66628 572704 66680 572756
rect 96896 572704 96948 572756
rect 111800 572704 111852 572756
rect 136640 572704 136692 572756
rect 137100 572704 137152 572756
rect 191564 572704 191616 572756
rect 255412 572704 255464 572756
rect 283564 572704 283616 572756
rect 97908 572636 97960 572688
rect 112444 572636 112496 572688
rect 184296 572636 184348 572688
rect 191288 572636 191340 572688
rect 111800 571956 111852 572008
rect 183376 571956 183428 572008
rect 60648 571344 60700 571396
rect 66628 571344 66680 571396
rect 97724 571344 97776 571396
rect 101404 571344 101456 571396
rect 255412 571344 255464 571396
rect 278872 571344 278924 571396
rect 188344 571276 188396 571328
rect 190920 571276 190972 571328
rect 157248 570596 157300 570648
rect 182824 570664 182876 570716
rect 182916 570596 182968 570648
rect 183376 570596 183428 570648
rect 191564 570596 191616 570648
rect 255412 570596 255464 570648
rect 255688 570596 255740 570648
rect 582564 570596 582616 570648
rect 57888 569916 57940 569968
rect 66628 569916 66680 569968
rect 97908 569916 97960 569968
rect 146944 569916 146996 569968
rect 97448 569168 97500 569220
rect 178868 569168 178920 569220
rect 255412 568896 255464 568948
rect 258080 568896 258132 568948
rect 255412 568556 255464 568608
rect 289912 568556 289964 568608
rect 96804 568488 96856 568540
rect 129648 568488 129700 568540
rect 129004 567808 129056 567860
rect 186964 567808 187016 567860
rect 255504 567808 255556 567860
rect 281632 567808 281684 567860
rect 255780 567264 255832 567316
rect 258172 567264 258224 567316
rect 188804 567196 188856 567248
rect 191748 567196 191800 567248
rect 289728 566448 289780 566500
rect 582472 566448 582524 566500
rect 255688 565904 255740 565956
rect 274916 565904 274968 565956
rect 52368 565836 52420 565888
rect 67640 565836 67692 565888
rect 255596 565836 255648 565888
rect 288624 565836 288676 565888
rect 289728 565836 289780 565888
rect 187700 565768 187752 565820
rect 188896 565768 188948 565820
rect 190828 565768 190880 565820
rect 169208 565088 169260 565140
rect 187700 565088 187752 565140
rect 39948 564408 40000 564460
rect 66812 564408 66864 564460
rect 187700 564408 187752 564460
rect 191104 564408 191156 564460
rect 255596 564408 255648 564460
rect 269120 564408 269172 564460
rect 124864 563660 124916 563712
rect 191012 563660 191064 563712
rect 64696 563048 64748 563100
rect 66720 563048 66772 563100
rect 255596 563048 255648 563100
rect 277400 563048 277452 563100
rect 169576 561688 169628 561740
rect 191748 561688 191800 561740
rect 255596 561688 255648 561740
rect 259644 561688 259696 561740
rect 259368 561008 259420 561060
rect 266360 561008 266412 561060
rect 96896 560940 96948 560992
rect 180156 560940 180208 560992
rect 185676 560396 185728 560448
rect 191104 560396 191156 560448
rect 170956 560260 171008 560312
rect 191196 560260 191248 560312
rect 255596 560260 255648 560312
rect 260932 560260 260984 560312
rect 98092 559512 98144 559564
rect 115204 559512 115256 559564
rect 61936 558900 61988 558952
rect 66812 558900 66864 558952
rect 96988 558900 97040 558952
rect 113824 558900 113876 558952
rect 255596 558900 255648 558952
rect 273260 558900 273312 558952
rect 115204 558832 115256 558884
rect 160744 558832 160796 558884
rect 162768 558152 162820 558204
rect 187700 558152 187752 558204
rect 188344 557608 188396 557660
rect 190920 557608 190972 557660
rect 181996 557540 182048 557592
rect 191748 557540 191800 557592
rect 255596 557540 255648 557592
rect 266360 557540 266412 557592
rect 97908 556792 97960 556844
rect 115296 556792 115348 556844
rect 166448 556180 166500 556232
rect 191748 556180 191800 556232
rect 255596 556180 255648 556232
rect 288440 556180 288492 556232
rect 257344 555432 257396 555484
rect 280252 555432 280304 555484
rect 182824 554820 182876 554872
rect 188344 554820 188396 554872
rect 159456 554752 159508 554804
rect 180156 554752 180208 554804
rect 184664 554752 184716 554804
rect 190828 554752 190880 554804
rect 2780 553800 2832 553852
rect 4804 553800 4856 553852
rect 255596 553460 255648 553512
rect 260840 553460 260892 553512
rect 57796 553392 57848 553444
rect 66720 553392 66772 553444
rect 171784 553392 171836 553444
rect 190920 553392 190972 553444
rect 255688 553392 255740 553444
rect 277584 553392 277636 553444
rect 255596 552644 255648 552696
rect 259368 552644 259420 552696
rect 269212 552644 269264 552696
rect 97908 552304 97960 552356
rect 100760 552304 100812 552356
rect 167644 552032 167696 552084
rect 191748 552032 191800 552084
rect 105544 551284 105596 551336
rect 162216 551284 162268 551336
rect 255596 550672 255648 550724
rect 259552 550672 259604 550724
rect 161572 550604 161624 550656
rect 162216 550604 162268 550656
rect 191380 550604 191432 550656
rect 255596 550536 255648 550588
rect 269304 550536 269356 550588
rect 276112 550536 276164 550588
rect 97908 549856 97960 549908
rect 160100 549856 160152 549908
rect 160100 549244 160152 549296
rect 160744 549244 160796 549296
rect 188344 549312 188396 549364
rect 187700 549244 187752 549296
rect 191748 549244 191800 549296
rect 100760 548496 100812 548548
rect 112444 548496 112496 548548
rect 173624 548496 173676 548548
rect 187700 548496 187752 548548
rect 187424 547884 187476 547936
rect 191564 547884 191616 547936
rect 255596 547884 255648 547936
rect 263600 547884 263652 547936
rect 178684 546524 178736 546576
rect 191564 546524 191616 546576
rect 99380 546456 99432 546508
rect 191288 546456 191340 546508
rect 255596 546456 255648 546508
rect 271972 546456 272024 546508
rect 146944 545708 146996 545760
rect 188436 545708 188488 545760
rect 255596 545232 255648 545284
rect 258264 545232 258316 545284
rect 176476 545096 176528 545148
rect 191196 545096 191248 545148
rect 180156 545028 180208 545080
rect 190644 545028 190696 545080
rect 50988 543736 51040 543788
rect 66812 543736 66864 543788
rect 97540 543736 97592 543788
rect 104256 543736 104308 543788
rect 150256 543736 150308 543788
rect 191104 543736 191156 543788
rect 255596 543736 255648 543788
rect 266452 543736 266504 543788
rect 33784 542988 33836 543040
rect 65984 542988 66036 543040
rect 66536 542988 66588 543040
rect 165068 542444 165120 542496
rect 191564 542444 191616 542496
rect 97540 542376 97592 542428
rect 146116 542376 146168 542428
rect 189080 542376 189132 542428
rect 169760 542308 169812 542360
rect 179420 542308 179472 542360
rect 180064 542308 180116 542360
rect 278044 542308 278096 542360
rect 285864 542308 285916 542360
rect 97908 541628 97960 541680
rect 116584 541628 116636 541680
rect 155776 541628 155828 541680
rect 169760 541628 169812 541680
rect 166540 540948 166592 541000
rect 190828 540948 190880 541000
rect 255596 540948 255648 541000
rect 262312 540948 262364 541000
rect 7564 540200 7616 540252
rect 188344 540200 188396 540252
rect 191564 540200 191616 540252
rect 73160 539860 73212 539912
rect 67272 539792 67324 539844
rect 71780 539792 71832 539844
rect 59084 539588 59136 539640
rect 66628 539588 66680 539640
rect 91744 539588 91796 539640
rect 162860 539588 162912 539640
rect 170496 539588 170548 539640
rect 191472 539588 191524 539640
rect 253112 539316 253164 539368
rect 255688 539316 255740 539368
rect 122104 538840 122156 538892
rect 146944 538840 146996 538892
rect 43444 538296 43496 538348
rect 94596 538296 94648 538348
rect 104164 538296 104216 538348
rect 189080 538296 189132 538348
rect 221372 538296 221424 538348
rect 252100 538296 252152 538348
rect 258172 538296 258224 538348
rect 85856 538228 85908 538280
rect 96436 538228 96488 538280
rect 99380 538228 99432 538280
rect 177396 538228 177448 538280
rect 238668 538228 238720 538280
rect 255596 538228 255648 538280
rect 282920 538228 282972 538280
rect 4804 538160 4856 538212
rect 70952 538160 71004 538212
rect 79232 538160 79284 538212
rect 119436 538160 119488 538212
rect 178868 538160 178920 538212
rect 244372 538160 244424 538212
rect 62028 537480 62080 537532
rect 73160 537480 73212 537532
rect 144644 537480 144696 537532
rect 222108 537480 222160 537532
rect 244280 537480 244332 537532
rect 582380 537480 582432 537532
rect 79232 537004 79284 537056
rect 79968 537004 80020 537056
rect 59176 536800 59228 536852
rect 62028 536800 62080 536852
rect 88248 536800 88300 536852
rect 95424 536800 95476 536852
rect 244372 536800 244424 536852
rect 244832 536800 244884 536852
rect 249708 536800 249760 536852
rect 254124 536800 254176 536852
rect 73160 536732 73212 536784
rect 76748 536732 76800 536784
rect 93400 536732 93452 536784
rect 246764 536732 246816 536784
rect 285588 536800 285640 536852
rect 291200 536800 291252 536852
rect 82176 536664 82228 536716
rect 91744 536664 91796 536716
rect 239220 536664 239272 536716
rect 244280 536664 244332 536716
rect 68928 536528 68980 536580
rect 72424 536528 72476 536580
rect 195980 536188 196032 536240
rect 197636 536188 197688 536240
rect 244924 536120 244976 536172
rect 245936 536120 245988 536172
rect 3424 536052 3476 536104
rect 41328 536052 41380 536104
rect 69388 536052 69440 536104
rect 70952 536052 71004 536104
rect 86224 536052 86276 536104
rect 189816 536052 189868 536104
rect 193588 536052 193640 536104
rect 225236 536052 225288 536104
rect 226984 536052 227036 536104
rect 86684 535916 86736 535968
rect 87604 535916 87656 535968
rect 214656 535508 214708 535560
rect 216404 535508 216456 535560
rect 91008 535440 91060 535492
rect 91836 535440 91888 535492
rect 215944 535440 215996 535492
rect 216956 535440 217008 535492
rect 231676 535440 231728 535492
rect 233884 535440 233936 535492
rect 246304 535440 246356 535492
rect 247500 535440 247552 535492
rect 106924 535372 106976 535424
rect 143540 535372 143592 535424
rect 144644 535372 144696 535424
rect 163872 535372 163924 535424
rect 197360 535372 197412 535424
rect 206376 535236 206428 535288
rect 209964 535236 210016 535288
rect 217324 534828 217376 534880
rect 239772 534828 239824 534880
rect 231216 534760 231268 534812
rect 254032 534760 254084 534812
rect 48136 534692 48188 534744
rect 96896 534692 96948 534744
rect 178776 534692 178828 534744
rect 230388 534692 230440 534744
rect 251916 534692 251968 534744
rect 281724 534692 281776 534744
rect 162860 534420 162912 534472
rect 163872 534420 163924 534472
rect 67364 534012 67416 534064
rect 158720 534012 158772 534064
rect 180616 534012 180668 534064
rect 209412 534012 209464 534064
rect 158720 533536 158772 533588
rect 159456 533536 159508 533588
rect 195980 533400 196032 533452
rect 196900 533400 196952 533452
rect 197360 533400 197412 533452
rect 198188 533400 198240 533452
rect 82728 533332 82780 533384
rect 94688 533332 94740 533384
rect 187700 533332 187752 533384
rect 200396 533400 200448 533452
rect 211804 533400 211856 533452
rect 212540 533400 212592 533452
rect 213184 533400 213236 533452
rect 222660 533400 222712 533452
rect 227812 533400 227864 533452
rect 239404 533400 239456 533452
rect 244556 533400 244608 533452
rect 245016 533400 245068 533452
rect 248420 533400 248472 533452
rect 248972 533400 249024 533452
rect 250444 533400 250496 533452
rect 259644 533400 259696 533452
rect 201500 533332 201552 533384
rect 202052 533332 202104 533384
rect 206284 533332 206336 533384
rect 233240 533332 233292 533384
rect 233700 533332 233752 533384
rect 238668 533332 238720 533384
rect 273536 533332 273588 533384
rect 236644 533264 236696 533316
rect 209044 532924 209096 532976
rect 211252 532924 211304 532976
rect 240140 532856 240192 532908
rect 240692 532856 240744 532908
rect 112444 532652 112496 532704
rect 113088 532652 113140 532704
rect 187700 532652 187752 532704
rect 179328 532584 179380 532636
rect 206836 532584 206888 532636
rect 75828 532040 75880 532092
rect 96804 532040 96856 532092
rect 73436 531972 73488 532024
rect 102784 531972 102836 532024
rect 246212 531972 246264 532024
rect 281816 531972 281868 532024
rect 64696 531224 64748 531276
rect 223580 531224 223632 531276
rect 93124 531156 93176 531208
rect 94044 531156 94096 531208
rect 190368 530544 190420 530596
rect 200212 530544 200264 530596
rect 228364 530544 228416 530596
rect 247592 530544 247644 530596
rect 247684 530544 247736 530596
rect 256700 530544 256752 530596
rect 214564 529932 214616 529984
rect 219624 529932 219676 529984
rect 191656 529864 191708 529916
rect 198832 529864 198884 529916
rect 213920 529728 213972 529780
rect 214748 529728 214800 529780
rect 71872 529252 71924 529304
rect 122104 529252 122156 529304
rect 193128 529252 193180 529304
rect 207204 529252 207256 529304
rect 67456 529184 67508 529236
rect 126888 529184 126940 529236
rect 166540 529184 166592 529236
rect 204536 529184 204588 529236
rect 238024 529184 238076 529236
rect 242900 529184 242952 529236
rect 291292 529184 291344 529236
rect 3148 528504 3200 528556
rect 98000 528504 98052 528556
rect 104256 528504 104308 528556
rect 104808 528504 104860 528556
rect 197636 528504 197688 528556
rect 164976 527892 165028 527944
rect 205640 527892 205692 527944
rect 244924 527892 244976 527944
rect 266544 527892 266596 527944
rect 201592 527824 201644 527876
rect 248604 527824 248656 527876
rect 62028 526396 62080 526448
rect 96712 526396 96764 526448
rect 196072 526396 196124 526448
rect 219440 526396 219492 526448
rect 226248 526260 226300 526312
rect 229284 526260 229336 526312
rect 218704 525036 218756 525088
rect 237472 525036 237524 525088
rect 248512 525036 248564 525088
rect 265164 525036 265216 525088
rect 60648 524356 60700 524408
rect 165620 524356 165672 524408
rect 166448 524356 166500 524408
rect 187332 523744 187384 523796
rect 197452 523744 197504 523796
rect 196624 523676 196676 523728
rect 222200 523676 222252 523728
rect 146944 522928 146996 522980
rect 147404 522928 147456 522980
rect 214656 522928 214708 522980
rect 226984 522928 227036 522980
rect 229100 522928 229152 522980
rect 3424 522248 3476 522300
rect 93124 522248 93176 522300
rect 94504 522248 94556 522300
rect 244556 522248 244608 522300
rect 270684 522248 270736 522300
rect 203524 520956 203576 521008
rect 258172 520956 258224 521008
rect 141884 520888 141936 520940
rect 204260 520888 204312 520940
rect 128268 519596 128320 519648
rect 200120 519596 200172 519648
rect 178868 519528 178920 519580
rect 261024 519528 261076 519580
rect 171048 518236 171100 518288
rect 215944 518236 215996 518288
rect 72424 518168 72476 518220
rect 99472 518168 99524 518220
rect 137836 518168 137888 518220
rect 189816 518168 189868 518220
rect 195244 518168 195296 518220
rect 206376 518168 206428 518220
rect 65800 517148 65852 517200
rect 69664 517148 69716 517200
rect 204904 515448 204956 515500
rect 240232 515448 240284 515500
rect 63408 515380 63460 515432
rect 92572 515380 92624 515432
rect 147588 515380 147640 515432
rect 213184 515380 213236 515432
rect 233332 515380 233384 515432
rect 251456 515380 251508 515432
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 193496 514088 193548 514140
rect 202880 514088 202932 514140
rect 153016 514020 153068 514072
rect 251272 514020 251324 514072
rect 50988 513272 51040 513324
rect 169208 513272 169260 513324
rect 177396 512592 177448 512644
rect 208400 512592 208452 512644
rect 186228 511232 186280 511284
rect 205640 511232 205692 511284
rect 213184 511232 213236 511284
rect 230480 511232 230532 511284
rect 187516 510892 187568 510944
rect 191932 510892 191984 510944
rect 204996 509940 205048 509992
rect 253204 509940 253256 509992
rect 146208 509872 146260 509924
rect 205088 509872 205140 509924
rect 76012 509192 76064 509244
rect 212448 509192 212500 509244
rect 212448 508512 212500 508564
rect 222200 508512 222252 508564
rect 76012 508308 76064 508360
rect 76564 508308 76616 508360
rect 206376 507152 206428 507204
rect 258080 507152 258132 507204
rect 143264 507084 143316 507136
rect 247684 507084 247736 507136
rect 169484 505724 169536 505776
rect 254216 505724 254268 505776
rect 136548 504432 136600 504484
rect 195980 504432 196032 504484
rect 168104 504364 168156 504416
rect 232504 504364 232556 504416
rect 237380 504364 237432 504416
rect 253204 504364 253256 504416
rect 173532 502936 173584 502988
rect 244464 502936 244516 502988
rect 170772 501576 170824 501628
rect 253940 501576 253992 501628
rect 210424 500284 210476 500336
rect 253296 500284 253348 500336
rect 161204 500216 161256 500268
rect 217324 500216 217376 500268
rect 186964 498856 187016 498908
rect 216772 498856 216824 498908
rect 162676 498788 162728 498840
rect 195244 498788 195296 498840
rect 233884 497496 233936 497548
rect 277860 497496 277912 497548
rect 172244 497428 172296 497480
rect 250444 497428 250496 497480
rect 187424 496136 187476 496188
rect 214656 496136 214708 496188
rect 217324 496136 217376 496188
rect 231216 496136 231268 496188
rect 108948 496068 109000 496120
rect 277676 496068 277728 496120
rect 108304 495456 108356 495508
rect 108948 495456 109000 495508
rect 185584 494776 185636 494828
rect 214012 494776 214064 494828
rect 220912 494776 220964 494828
rect 256792 494776 256844 494828
rect 154488 494708 154540 494760
rect 222936 494708 222988 494760
rect 98000 492668 98052 492720
rect 210240 492668 210292 492720
rect 210516 492668 210568 492720
rect 157064 491988 157116 492040
rect 171784 491988 171836 492040
rect 165528 491920 165580 491972
rect 197360 491920 197412 491972
rect 227628 491920 227680 491972
rect 248420 491920 248472 491972
rect 184756 489132 184808 489184
rect 203524 489132 203576 489184
rect 222108 489132 222160 489184
rect 246304 489132 246356 489184
rect 166540 487840 166592 487892
rect 220084 487840 220136 487892
rect 187516 487772 187568 487824
rect 251824 487772 251876 487824
rect 236000 486684 236052 486736
rect 238116 486684 238168 486736
rect 210516 486480 210568 486532
rect 232504 486480 232556 486532
rect 160008 486412 160060 486464
rect 184664 486412 184716 486464
rect 218152 486412 218204 486464
rect 199476 485052 199528 485104
rect 241612 485052 241664 485104
rect 155684 484440 155736 484492
rect 182916 484440 182968 484492
rect 183376 484440 183428 484492
rect 122748 484372 122800 484424
rect 223580 484372 223632 484424
rect 183376 484304 183428 484356
rect 579804 484304 579856 484356
rect 178960 483624 179012 483676
rect 195428 483624 195480 483676
rect 233240 483624 233292 483676
rect 249800 483624 249852 483676
rect 242900 482944 242952 482996
rect 243544 482944 243596 482996
rect 177488 482264 177540 482316
rect 217324 482264 217376 482316
rect 239404 482264 239456 482316
rect 276204 482264 276256 482316
rect 133788 481652 133840 481704
rect 242900 481652 242952 481704
rect 181904 480292 181956 480344
rect 267924 480292 267976 480344
rect 126244 480224 126296 480276
rect 240784 480224 240836 480276
rect 176384 479476 176436 479528
rect 213920 479476 213972 479528
rect 218060 479476 218112 479528
rect 254124 479476 254176 479528
rect 132408 478932 132460 478984
rect 199476 478932 199528 478984
rect 198740 478864 198792 478916
rect 199384 478864 199436 478916
rect 215300 478864 215352 478916
rect 148784 478184 148836 478236
rect 198740 478184 198792 478236
rect 111064 478116 111116 478168
rect 251456 478116 251508 478168
rect 110420 477504 110472 477556
rect 111064 477504 111116 477556
rect 251456 477504 251508 477556
rect 251916 477504 251968 477556
rect 85488 476756 85540 476808
rect 94136 476756 94188 476808
rect 224960 476756 225012 476808
rect 269764 476756 269816 476808
rect 198740 476552 198792 476604
rect 199476 476552 199528 476604
rect 141424 476076 141476 476128
rect 258264 476076 258316 476128
rect 3332 475328 3384 475380
rect 43444 475328 43496 475380
rect 206468 475328 206520 475380
rect 222844 475328 222896 475380
rect 226340 474784 226392 474836
rect 226984 474784 227036 474836
rect 302240 474784 302292 474836
rect 164056 474716 164108 474768
rect 251364 474716 251416 474768
rect 146944 474648 146996 474700
rect 147404 474648 147456 474700
rect 146944 473424 146996 473476
rect 253480 473424 253532 473476
rect 108856 473356 108908 473408
rect 249064 473356 249116 473408
rect 93952 472608 94004 472660
rect 94596 472608 94648 472660
rect 209780 472608 209832 472660
rect 217324 472608 217376 472660
rect 269212 472608 269264 472660
rect 287060 472608 287112 472660
rect 287612 472608 287664 472660
rect 582472 472608 582524 472660
rect 151084 471996 151136 472048
rect 186044 471996 186096 472048
rect 229100 471996 229152 472048
rect 102140 471928 102192 471980
rect 102784 471928 102836 471980
rect 79968 471248 80020 471300
rect 101404 471248 101456 471300
rect 246948 471248 247000 471300
rect 249708 471248 249760 471300
rect 287060 471248 287112 471300
rect 251180 471112 251232 471164
rect 251824 471112 251876 471164
rect 135904 470636 135956 470688
rect 251180 470636 251232 470688
rect 102140 470568 102192 470620
rect 240232 470568 240284 470620
rect 180616 469820 180668 469872
rect 206284 469820 206336 469872
rect 228456 469820 228508 469872
rect 239404 469820 239456 469872
rect 174544 469208 174596 469260
rect 175004 469208 175056 469260
rect 242164 469208 242216 469260
rect 241428 469140 241480 469192
rect 259552 469140 259604 469192
rect 195336 468528 195388 468580
rect 213184 468528 213236 468580
rect 223580 468528 223632 468580
rect 246948 468528 247000 468580
rect 79324 468460 79376 468512
rect 91192 468460 91244 468512
rect 93860 468460 93912 468512
rect 160744 468460 160796 468512
rect 227720 468460 227772 468512
rect 240232 468460 240284 468512
rect 241428 468460 241480 468512
rect 197360 467100 197412 467152
rect 255504 467100 255556 467152
rect 140596 466488 140648 466540
rect 204260 466488 204312 466540
rect 68928 466420 68980 466472
rect 188344 466420 188396 466472
rect 224960 466420 225012 466472
rect 226248 466420 226300 466472
rect 299572 466420 299624 466472
rect 158444 465672 158496 465724
rect 165068 465672 165120 465724
rect 183284 465672 183336 465724
rect 191932 465672 191984 465724
rect 193036 465672 193088 465724
rect 212724 465672 212776 465724
rect 94504 465536 94556 465588
rect 95148 465536 95200 465588
rect 95148 465060 95200 465112
rect 216680 465060 216732 465112
rect 237380 465060 237432 465112
rect 238024 465060 238076 465112
rect 290004 465060 290056 465112
rect 201500 464992 201552 465044
rect 207112 464992 207164 465044
rect 77300 464312 77352 464364
rect 110512 464312 110564 464364
rect 130384 464312 130436 464364
rect 197360 464312 197412 464364
rect 273904 464312 273956 464364
rect 280252 464312 280304 464364
rect 165620 464176 165672 464228
rect 166448 464176 166500 464228
rect 226340 463768 226392 463820
rect 227628 463768 227680 463820
rect 274732 463768 274784 463820
rect 106280 463700 106332 463752
rect 165620 463700 165672 463752
rect 167644 463700 167696 463752
rect 248420 463700 248472 463752
rect 248604 463700 248656 463752
rect 204260 463632 204312 463684
rect 273444 463632 273496 463684
rect 87604 462952 87656 463004
rect 104900 462952 104952 463004
rect 190276 462952 190328 463004
rect 204996 462952 205048 463004
rect 3424 462408 3476 462460
rect 7564 462408 7616 462460
rect 104900 462340 104952 462392
rect 242992 462340 243044 462392
rect 82820 462272 82872 462324
rect 108856 462272 108908 462324
rect 109040 462272 109092 462324
rect 251180 462272 251232 462324
rect 251916 462272 251968 462324
rect 216680 461660 216732 461712
rect 231860 461660 231912 461712
rect 67640 461592 67692 461644
rect 83464 461592 83516 461644
rect 110512 461592 110564 461644
rect 117320 461592 117372 461644
rect 213828 461592 213880 461644
rect 270592 461592 270644 461644
rect 216680 461524 216732 461576
rect 217324 461524 217376 461576
rect 184664 460980 184716 461032
rect 216680 460980 216732 461032
rect 104808 460912 104860 460964
rect 188160 460912 188212 460964
rect 251180 460912 251232 460964
rect 292672 460912 292724 460964
rect 66168 460164 66220 460216
rect 85672 460164 85724 460216
rect 86224 460164 86276 460216
rect 114560 460164 114612 460216
rect 142804 460164 142856 460216
rect 249800 460164 249852 460216
rect 259552 460164 259604 460216
rect 112444 459552 112496 459604
rect 113088 459552 113140 459604
rect 129648 459552 129700 459604
rect 249616 459552 249668 459604
rect 187792 459484 187844 459536
rect 211804 459484 211856 459536
rect 253204 458872 253256 458924
rect 262404 458872 262456 458924
rect 241520 458804 241572 458856
rect 254032 458804 254084 458856
rect 276296 458668 276348 458720
rect 277308 458668 277360 458720
rect 278872 458668 278924 458720
rect 160744 458260 160796 458312
rect 197360 458260 197412 458312
rect 198004 458260 198056 458312
rect 75184 458192 75236 458244
rect 75828 458192 75880 458244
rect 187700 458192 187752 458244
rect 100024 457444 100076 457496
rect 142896 457444 142948 457496
rect 154028 457444 154080 457496
rect 187608 457444 187660 457496
rect 188160 457444 188212 457496
rect 246396 457444 246448 457496
rect 247500 457444 247552 457496
rect 277676 457444 277728 457496
rect 156604 457376 156656 457428
rect 163504 457376 163556 457428
rect 184204 456764 184256 456816
rect 213276 456764 213328 456816
rect 213828 456764 213880 456816
rect 237472 456764 237524 456816
rect 238116 456764 238168 456816
rect 253572 456764 253624 456816
rect 187516 456084 187568 456136
rect 188344 456084 188396 456136
rect 218152 456084 218204 456136
rect 218980 456084 219032 456136
rect 251272 456084 251324 456136
rect 252100 456084 252152 456136
rect 187700 456016 187752 456068
rect 196072 456016 196124 456068
rect 240140 456016 240192 456068
rect 254216 456016 254268 456068
rect 288348 456016 288400 456068
rect 580172 456016 580224 456068
rect 225052 455744 225104 455796
rect 226984 455744 227036 455796
rect 82084 455404 82136 455456
rect 82728 455404 82780 455456
rect 211160 455404 211212 455456
rect 233976 455404 234028 455456
rect 258080 455404 258132 455456
rect 73160 455336 73212 455388
rect 112996 455336 113048 455388
rect 129004 455336 129056 455388
rect 214656 455336 214708 455388
rect 242992 455336 243044 455388
rect 243544 455336 243596 455388
rect 276112 455336 276164 455388
rect 276388 455336 276440 455388
rect 221648 455268 221700 455320
rect 222108 455268 222160 455320
rect 63408 454656 63460 454708
rect 74540 454656 74592 454708
rect 154396 454656 154448 454708
rect 178868 454656 178920 454708
rect 276388 454656 276440 454708
rect 280252 454656 280304 454708
rect 188436 454112 188488 454164
rect 207112 454112 207164 454164
rect 187056 454044 187108 454096
rect 209872 454044 209924 454096
rect 210424 454044 210476 454096
rect 221648 454044 221700 454096
rect 261116 454044 261168 454096
rect 221188 453976 221240 454028
rect 223488 453976 223540 454028
rect 227812 453976 227864 454028
rect 228732 453976 228784 454028
rect 249616 453976 249668 454028
rect 253388 453976 253440 454028
rect 260104 453976 260156 454028
rect 262312 453976 262364 454028
rect 198832 453908 198884 453960
rect 200396 453908 200448 453960
rect 194508 453296 194560 453348
rect 241428 453296 241480 453348
rect 122196 452684 122248 452736
rect 195244 452684 195296 452736
rect 77944 452616 77996 452668
rect 166448 452616 166500 452668
rect 204168 452616 204220 452668
rect 218704 452616 218756 452668
rect 223028 452616 223080 452668
rect 260104 452616 260156 452668
rect 75828 451868 75880 451920
rect 98736 451868 98788 451920
rect 105544 451868 105596 451920
rect 158812 451868 158864 451920
rect 279424 451868 279476 451920
rect 287152 451868 287204 451920
rect 182180 451324 182232 451376
rect 195612 451324 195664 451376
rect 227720 451324 227772 451376
rect 272064 451324 272116 451376
rect 116584 451256 116636 451308
rect 240140 451256 240192 451308
rect 241336 451256 241388 451308
rect 261024 451256 261076 451308
rect 240692 451188 240744 451240
rect 251824 450984 251876 451036
rect 256976 450984 257028 451036
rect 113824 450644 113876 450696
rect 114468 450644 114520 450696
rect 180064 450576 180116 450628
rect 188804 450576 188856 450628
rect 4804 450508 4856 450560
rect 104164 450508 104216 450560
rect 184296 450508 184348 450560
rect 204168 450508 204220 450560
rect 193220 450236 193272 450288
rect 193496 450236 193548 450288
rect 114468 449964 114520 450016
rect 172336 449964 172388 450016
rect 78680 449896 78732 449948
rect 175004 449896 175056 449948
rect 188804 449896 188856 449948
rect 250904 449896 250956 449948
rect 258172 449896 258224 449948
rect 192760 449760 192812 449812
rect 195336 449760 195388 449812
rect 172336 449692 172388 449744
rect 194508 449692 194560 449744
rect 251916 449692 251968 449744
rect 95240 449216 95292 449268
rect 151084 449216 151136 449268
rect 57888 449148 57940 449200
rect 169024 449148 169076 449200
rect 268016 449148 268068 449200
rect 184848 449080 184900 449132
rect 191564 449080 191616 449132
rect 3148 448536 3200 448588
rect 36544 448536 36596 448588
rect 66076 448536 66128 448588
rect 70492 448536 70544 448588
rect 95148 448536 95200 448588
rect 95884 448536 95936 448588
rect 177580 447856 177632 447908
rect 188436 447856 188488 447908
rect 66168 447788 66220 447840
rect 191564 447788 191616 447840
rect 176108 447040 176160 447092
rect 176476 447040 176528 447092
rect 191012 447040 191064 447092
rect 67180 446428 67232 446480
rect 165068 446428 165120 446480
rect 76656 446360 76708 446412
rect 176108 446360 176160 446412
rect 255596 446360 255648 446412
rect 269212 446360 269264 446412
rect 173716 445748 173768 445800
rect 177304 445748 177356 445800
rect 160100 445680 160152 445732
rect 160744 445680 160796 445732
rect 191012 445680 191064 445732
rect 143356 445000 143408 445052
rect 184204 445000 184256 445052
rect 269764 445000 269816 445052
rect 278872 445000 278924 445052
rect 83464 444456 83516 444508
rect 142896 444456 142948 444508
rect 143356 444456 143408 444508
rect 72424 444388 72476 444440
rect 160100 444388 160152 444440
rect 86960 444320 87012 444372
rect 88248 444320 88300 444372
rect 255504 443844 255556 443896
rect 88248 443708 88300 443760
rect 184296 443708 184348 443760
rect 68928 443640 68980 443692
rect 80060 443640 80112 443692
rect 184572 443640 184624 443692
rect 187148 443640 187200 443692
rect 258264 443640 258316 443692
rect 269304 443640 269356 443692
rect 71136 442960 71188 443012
rect 193036 443028 193088 443080
rect 257344 442280 257396 442332
rect 263692 442280 263744 442332
rect 163964 442212 164016 442264
rect 190276 442212 190328 442264
rect 191564 442212 191616 442264
rect 255504 442212 255556 442264
rect 259644 442212 259696 442264
rect 285772 442212 285824 442264
rect 61844 441668 61896 441720
rect 138664 441668 138716 441720
rect 68284 441600 68336 441652
rect 163964 441600 164016 441652
rect 173624 441532 173676 441584
rect 191564 441532 191616 441584
rect 104164 441464 104216 441516
rect 174544 441464 174596 441516
rect 69756 440852 69808 440904
rect 122196 440852 122248 440904
rect 190276 440852 190328 440904
rect 193312 440852 193364 440904
rect 183376 440240 183428 440292
rect 186964 440240 187016 440292
rect 76840 439560 76892 439612
rect 89720 439560 89772 439612
rect 50988 439492 51040 439544
rect 83740 439492 83792 439544
rect 255504 439492 255556 439544
rect 288716 439492 288768 439544
rect 183468 438948 183520 439000
rect 186964 438948 187016 439000
rect 104808 438880 104860 438932
rect 107660 438880 107712 438932
rect 186044 438880 186096 438932
rect 187700 438880 187752 438932
rect 147680 438812 147732 438864
rect 148692 438812 148744 438864
rect 191656 438812 191708 438864
rect 255504 438812 255556 438864
rect 263784 438812 263836 438864
rect 255964 438744 256016 438796
rect 260196 438744 260248 438796
rect 73896 438200 73948 438252
rect 77944 438200 77996 438252
rect 67364 438132 67416 438184
rect 76656 438132 76708 438184
rect 81440 438132 81492 438184
rect 88984 438132 89036 438184
rect 90640 438132 90692 438184
rect 147680 438132 147732 438184
rect 78588 437452 78640 437504
rect 176476 437452 176528 437504
rect 177580 437452 177632 437504
rect 183468 437452 183520 437504
rect 184572 437452 184624 437504
rect 263784 437452 263836 437504
rect 266636 437452 266688 437504
rect 76564 437384 76616 437436
rect 82912 437384 82964 437436
rect 101404 437384 101456 437436
rect 104164 437384 104216 437436
rect 102508 437316 102560 437368
rect 105544 437316 105596 437368
rect 110788 436704 110840 436756
rect 180064 436704 180116 436756
rect 95884 436296 95936 436348
rect 96988 436296 97040 436348
rect 52276 436160 52328 436212
rect 68928 436228 68980 436280
rect 41236 436092 41288 436144
rect 70492 436160 70544 436212
rect 68652 436092 68704 436144
rect 71780 436160 71832 436212
rect 72700 436160 72752 436212
rect 71688 436092 71740 436144
rect 72424 436092 72476 436144
rect 96344 436092 96396 436144
rect 100024 436092 100076 436144
rect 103888 436092 103940 436144
rect 104164 436092 104216 436144
rect 116032 436092 116084 436144
rect 116584 436092 116636 436144
rect 188344 436092 188396 436144
rect 191656 436092 191708 436144
rect 255504 436024 255556 436076
rect 267924 436024 267976 436076
rect 276296 436024 276348 436076
rect 170404 435344 170456 435396
rect 181536 435344 181588 435396
rect 264244 435344 264296 435396
rect 274824 435344 274876 435396
rect 3424 434800 3476 434852
rect 112260 434800 112312 434852
rect 62028 434732 62080 434784
rect 191656 434732 191708 434784
rect 115756 434664 115808 434716
rect 126244 434664 126296 434716
rect 68192 433984 68244 434036
rect 191656 433984 191708 434036
rect 255504 433984 255556 434036
rect 262864 433984 262916 434036
rect 67272 433780 67324 433832
rect 71136 433780 71188 433832
rect 70676 433644 70728 433696
rect 53748 433304 53800 433356
rect 57704 433304 57756 433356
rect 66812 433304 66864 433356
rect 67732 433236 67784 433288
rect 276020 433304 276072 433356
rect 115848 433236 115900 433288
rect 146944 433236 146996 433288
rect 155592 433236 155644 433288
rect 155776 433236 155828 433288
rect 269028 433236 269080 433288
rect 67548 433168 67600 433220
rect 68284 433168 68336 433220
rect 155592 432556 155644 432608
rect 191656 432556 191708 432608
rect 262864 432556 262916 432608
rect 267924 432556 267976 432608
rect 269028 432556 269080 432608
rect 65708 432488 65760 432540
rect 66168 432488 66220 432540
rect 63316 431944 63368 431996
rect 178960 431944 179012 431996
rect 254216 431944 254268 431996
rect 263784 431944 263836 431996
rect 56508 431196 56560 431248
rect 67364 431196 67416 431248
rect 165436 431196 165488 431248
rect 191748 431196 191800 431248
rect 255412 431196 255464 431248
rect 262496 431196 262548 431248
rect 138664 430516 138716 430568
rect 164976 430516 165028 430568
rect 165436 430516 165488 430568
rect 178960 430516 179012 430568
rect 191012 430516 191064 430568
rect 114928 430448 114980 430500
rect 141424 430448 141476 430500
rect 155776 429836 155828 429888
rect 188344 429836 188396 429888
rect 255412 429496 255464 429548
rect 259552 429496 259604 429548
rect 64696 429360 64748 429412
rect 67272 429360 67324 429412
rect 48228 429156 48280 429208
rect 66812 429156 66864 429208
rect 115848 429088 115900 429140
rect 154028 429088 154080 429140
rect 154396 429088 154448 429140
rect 190828 429088 190880 429140
rect 65800 427320 65852 427372
rect 67548 427320 67600 427372
rect 122196 427048 122248 427100
rect 133144 427048 133196 427100
rect 169024 427048 169076 427100
rect 178040 427048 178092 427100
rect 284392 427048 284444 427100
rect 291384 427048 291436 427100
rect 582564 427048 582616 427100
rect 115848 426436 115900 426488
rect 125600 426436 125652 426488
rect 178040 426436 178092 426488
rect 179328 426436 179380 426488
rect 191748 426436 191800 426488
rect 255412 426436 255464 426488
rect 284392 426436 284444 426488
rect 67548 426368 67600 426420
rect 68192 426368 68244 426420
rect 115756 426368 115808 426420
rect 117504 426368 117556 426420
rect 119344 426368 119396 426420
rect 49608 425688 49660 425740
rect 66996 425688 67048 425740
rect 256608 425688 256660 425740
rect 273536 425688 273588 425740
rect 165620 425076 165672 425128
rect 191748 425076 191800 425128
rect 115848 425008 115900 425060
rect 130384 425008 130436 425060
rect 151728 425008 151780 425060
rect 182088 425008 182140 425060
rect 191012 425008 191064 425060
rect 115112 424940 115164 424992
rect 117320 424940 117372 424992
rect 169392 424464 169444 424516
rect 182088 424464 182140 424516
rect 169576 424328 169628 424380
rect 182824 424328 182876 424380
rect 256608 424328 256660 424380
rect 274824 424328 274876 424380
rect 59268 423648 59320 423700
rect 66720 423648 66772 423700
rect 60740 423580 60792 423632
rect 62028 423580 62080 423632
rect 66812 423580 66864 423632
rect 115848 423580 115900 423632
rect 170404 423580 170456 423632
rect 146116 423512 146168 423564
rect 151084 423512 151136 423564
rect 253572 423376 253624 423428
rect 256976 423376 257028 423428
rect 44088 422900 44140 422952
rect 60740 422900 60792 422952
rect 151084 422288 151136 422340
rect 191748 422288 191800 422340
rect 255504 422288 255556 422340
rect 277768 422288 277820 422340
rect 152924 421540 152976 421592
rect 177396 421540 177448 421592
rect 65984 420996 66036 421048
rect 67548 420996 67600 421048
rect 50988 420928 51040 420980
rect 66812 420928 66864 420980
rect 146116 420928 146168 420980
rect 152556 420928 152608 420980
rect 153108 420928 153160 420980
rect 255504 420928 255556 420980
rect 298284 420928 298336 420980
rect 61844 420860 61896 420912
rect 66904 420860 66956 420912
rect 57888 420180 57940 420232
rect 66812 420180 66864 420232
rect 186964 420180 187016 420232
rect 192484 420180 192536 420232
rect 174636 419500 174688 419552
rect 192392 419500 192444 419552
rect 255504 419500 255556 419552
rect 280436 419500 280488 419552
rect 285864 419500 285916 419552
rect 115848 419432 115900 419484
rect 142804 419432 142856 419484
rect 255412 419432 255464 419484
rect 281540 419432 281592 419484
rect 122104 419364 122156 419416
rect 123024 419364 123076 419416
rect 281540 418752 281592 418804
rect 285864 418752 285916 418804
rect 582380 418752 582432 418804
rect 63224 418276 63276 418328
rect 66444 418276 66496 418328
rect 63408 418072 63460 418124
rect 66444 418072 66496 418124
rect 153108 417392 153160 417444
rect 155684 417392 155736 417444
rect 179420 417392 179472 417444
rect 283656 417392 283708 417444
rect 582656 417392 582708 417444
rect 117412 417188 117464 417240
rect 122196 417188 122248 417240
rect 126244 417188 126296 417240
rect 126888 417188 126940 417240
rect 57796 416780 57848 416832
rect 115848 416780 115900 416832
rect 117412 416780 117464 416832
rect 126888 416780 126940 416832
rect 148324 416780 148376 416832
rect 177304 416780 177356 416832
rect 191748 416780 191800 416832
rect 255504 416780 255556 416832
rect 283196 416780 283248 416832
rect 283656 416780 283708 416832
rect 61844 416712 61896 416764
rect 179420 416712 179472 416764
rect 191656 416712 191708 416764
rect 255412 416712 255464 416764
rect 278964 416712 279016 416764
rect 279332 416712 279384 416764
rect 122104 416032 122156 416084
rect 189724 416032 189776 416084
rect 115848 415624 115900 415676
rect 120080 415624 120132 415676
rect 61844 415420 61896 415472
rect 66904 415420 66956 415472
rect 114928 414672 114980 414724
rect 124864 414672 124916 414724
rect 176568 414672 176620 414724
rect 189724 414672 189776 414724
rect 54852 413992 54904 414044
rect 66812 413992 66864 414044
rect 154028 413992 154080 414044
rect 191196 413992 191248 414044
rect 57980 413244 58032 413296
rect 66628 413244 66680 413296
rect 123024 412700 123076 412752
rect 142804 412700 142856 412752
rect 115848 412632 115900 412684
rect 147036 412632 147088 412684
rect 115756 412564 115808 412616
rect 123024 412564 123076 412616
rect 255504 412564 255556 412616
rect 281816 412564 281868 412616
rect 52184 411884 52236 411936
rect 55036 411884 55088 411936
rect 57980 411884 58032 411936
rect 165436 411884 165488 411936
rect 191748 411884 191800 411936
rect 64788 411272 64840 411324
rect 66904 411272 66956 411324
rect 115848 411204 115900 411256
rect 126244 411204 126296 411256
rect 60004 410524 60056 410576
rect 66812 410524 66864 410576
rect 154396 410524 154448 410576
rect 161480 410524 161532 410576
rect 183192 410524 183244 410576
rect 191748 410524 191800 410576
rect 115940 409844 115992 409896
rect 154396 409844 154448 409896
rect 135996 409776 136048 409828
rect 141884 409776 141936 409828
rect 177304 409776 177356 409828
rect 115848 409708 115900 409760
rect 122104 409708 122156 409760
rect 39856 409096 39908 409148
rect 52368 409096 52420 409148
rect 60004 409096 60056 409148
rect 129004 409096 129056 409148
rect 135996 409096 136048 409148
rect 153844 409096 153896 409148
rect 184296 409096 184348 409148
rect 271788 409096 271840 409148
rect 280160 409096 280212 409148
rect 63316 408484 63368 408536
rect 66444 408484 66496 408536
rect 115848 408484 115900 408536
rect 141424 408484 141476 408536
rect 255412 408484 255464 408536
rect 270776 408484 270828 408536
rect 271788 408484 271840 408536
rect 255412 407804 255464 407856
rect 262404 407804 262456 407856
rect 48136 407736 48188 407788
rect 66812 407736 66864 407788
rect 186136 407736 186188 407788
rect 193312 407736 193364 407788
rect 255504 407736 255556 407788
rect 267832 407736 267884 407788
rect 124864 407124 124916 407176
rect 185584 407124 185636 407176
rect 113088 407056 113140 407108
rect 135904 407056 135956 407108
rect 50896 406376 50948 406428
rect 64604 406376 64656 406428
rect 66444 406376 66496 406428
rect 119344 406376 119396 406428
rect 143264 406376 143316 406428
rect 177396 406376 177448 406428
rect 186136 405968 186188 406020
rect 187056 405968 187108 406020
rect 191012 405696 191064 405748
rect 255504 405696 255556 405748
rect 281816 405696 281868 405748
rect 153016 405628 153068 405680
rect 161480 405628 161532 405680
rect 181628 405628 181680 405680
rect 181996 405628 182048 405680
rect 191748 405628 191800 405680
rect 62028 404336 62080 404388
rect 66904 404336 66956 404388
rect 115848 404336 115900 404388
rect 146944 404336 146996 404388
rect 178868 404336 178920 404388
rect 181628 404336 181680 404388
rect 154304 404268 154356 404320
rect 158720 404268 158772 404320
rect 162768 404268 162820 404320
rect 191748 404268 191800 404320
rect 262864 403588 262916 403640
rect 270500 403588 270552 403640
rect 119988 403044 120040 403096
rect 154304 403044 154356 403096
rect 54760 402976 54812 403028
rect 66444 402976 66496 403028
rect 115848 402976 115900 403028
rect 151176 402976 151228 403028
rect 157984 402976 158036 403028
rect 162768 402976 162820 403028
rect 255412 402976 255464 403028
rect 291384 402976 291436 403028
rect 55128 402908 55180 402960
rect 67640 402908 67692 402960
rect 161388 402296 161440 402348
rect 176660 402296 176712 402348
rect 115940 402228 115992 402280
rect 184756 402228 184808 402280
rect 184756 401684 184808 401736
rect 186964 401684 187016 401736
rect 176660 401616 176712 401668
rect 177948 401616 178000 401668
rect 191012 401616 191064 401668
rect 255412 401616 255464 401668
rect 259552 401616 259604 401668
rect 169024 401548 169076 401600
rect 173532 401548 173584 401600
rect 191748 401548 191800 401600
rect 114836 400936 114888 400988
rect 119988 400936 120040 400988
rect 118792 400868 118844 400920
rect 143540 400868 143592 400920
rect 177856 400596 177908 400648
rect 178776 400596 178828 400648
rect 58992 400188 59044 400240
rect 66444 400188 66496 400240
rect 115388 400188 115440 400240
rect 122104 400188 122156 400240
rect 129004 400188 129056 400240
rect 177856 400188 177908 400240
rect 255412 400188 255464 400240
rect 280344 400188 280396 400240
rect 147036 399440 147088 399492
rect 180248 399440 180300 399492
rect 53656 398828 53708 398880
rect 66812 398828 66864 398880
rect 188344 398828 188396 398880
rect 191012 398828 191064 398880
rect 61936 398760 61988 398812
rect 67088 398760 67140 398812
rect 276480 398760 276532 398812
rect 277492 398760 277544 398812
rect 115848 398284 115900 398336
rect 116124 398284 116176 398336
rect 118792 398284 118844 398336
rect 253572 398148 253624 398200
rect 262496 398148 262548 398200
rect 118792 398080 118844 398132
rect 149060 398080 149112 398132
rect 255412 398080 255464 398132
rect 276020 398080 276072 398132
rect 276480 398080 276532 398132
rect 168104 397536 168156 397588
rect 169760 397536 169812 397588
rect 190828 397536 190880 397588
rect 4804 397468 4856 397520
rect 64604 397468 64656 397520
rect 66812 397468 66864 397520
rect 126244 397468 126296 397520
rect 178684 397468 178736 397520
rect 162124 397264 162176 397316
rect 162676 397264 162728 397316
rect 115756 397060 115808 397112
rect 118792 397060 118844 397112
rect 41328 396720 41380 396772
rect 60740 396720 60792 396772
rect 130384 396720 130436 396772
rect 137928 396720 137980 396772
rect 180892 396720 180944 396772
rect 258724 396720 258776 396772
rect 276204 396720 276256 396772
rect 60740 396040 60792 396092
rect 61936 396040 61988 396092
rect 66260 396040 66312 396092
rect 115848 396040 115900 396092
rect 124956 396040 125008 396092
rect 162124 396040 162176 396092
rect 192668 396040 192720 396092
rect 153016 395972 153068 396024
rect 156604 395972 156656 396024
rect 162216 395972 162268 396024
rect 170864 395972 170916 396024
rect 191748 395972 191800 396024
rect 259000 395292 259052 395344
rect 273444 395292 273496 395344
rect 115848 394748 115900 394800
rect 144184 394748 144236 394800
rect 115848 394612 115900 394664
rect 153016 394680 153068 394732
rect 255412 394680 255464 394732
rect 272156 394680 272208 394732
rect 117228 394000 117280 394052
rect 136640 394000 136692 394052
rect 137284 394000 137336 394052
rect 159364 394000 159416 394052
rect 118608 393932 118660 393984
rect 163872 393932 163924 393984
rect 171968 393932 172020 393984
rect 178684 393932 178736 393984
rect 187976 393932 188028 393984
rect 256700 393932 256752 393984
rect 278872 393932 278924 393984
rect 60556 393320 60608 393372
rect 67732 393320 67784 393372
rect 166356 393320 166408 393372
rect 177488 393320 177540 393372
rect 255412 393320 255464 393372
rect 278872 393320 278924 393372
rect 115940 392708 115992 392760
rect 117228 392708 117280 392760
rect 142988 392572 143040 392624
rect 158536 392572 158588 392624
rect 179420 392572 179472 392624
rect 254032 392096 254084 392148
rect 255504 392096 255556 392148
rect 60556 391960 60608 392012
rect 66628 391960 66680 392012
rect 115848 391960 115900 392012
rect 141608 391960 141660 392012
rect 168196 391960 168248 392012
rect 186320 391960 186372 392012
rect 68560 391892 68612 391944
rect 161204 391892 161256 391944
rect 177488 391280 177540 391332
rect 193220 391280 193272 391332
rect 259276 391280 259328 391332
rect 298192 391280 298244 391332
rect 43444 391212 43496 391264
rect 189724 391212 189776 391264
rect 93952 390940 94004 390992
rect 193220 390940 193272 390992
rect 194140 390940 194192 390992
rect 218336 390940 218388 390992
rect 218796 390940 218848 390992
rect 251732 390940 251784 390992
rect 273904 391212 273956 391264
rect 283564 391212 283616 391264
rect 291476 391212 291528 391264
rect 582380 391212 582432 391264
rect 89904 390600 89956 390652
rect 90456 390600 90508 390652
rect 100392 390532 100444 390584
rect 179144 390532 179196 390584
rect 179512 390532 179564 390584
rect 67824 390124 67876 390176
rect 68790 390124 68842 390176
rect 96712 390124 96764 390176
rect 97862 390124 97914 390176
rect 100806 390124 100858 390176
rect 101956 390124 102008 390176
rect 104808 389784 104860 389836
rect 114836 389784 114888 389836
rect 156696 389784 156748 389836
rect 168380 389784 168432 389836
rect 179236 389784 179288 389836
rect 180892 389784 180944 389836
rect 277308 389784 277360 389836
rect 281540 389784 281592 389836
rect 36544 389240 36596 389292
rect 100760 389240 100812 389292
rect 168380 389240 168432 389292
rect 169484 389240 169536 389292
rect 202052 389240 202104 389292
rect 230572 389240 230624 389292
rect 256700 389240 256752 389292
rect 3516 389172 3568 389224
rect 107660 389172 107712 389224
rect 118608 389172 118660 389224
rect 187976 389172 188028 389224
rect 240140 389172 240192 389224
rect 241060 389172 241112 389224
rect 241520 389172 241572 389224
rect 264244 389172 264296 389224
rect 157156 389104 157208 389156
rect 161572 389104 161624 389156
rect 176384 389104 176436 389156
rect 197268 389104 197320 389156
rect 250444 389104 250496 389156
rect 281632 389104 281684 389156
rect 253388 389036 253440 389088
rect 271972 389036 272024 389088
rect 59176 388424 59228 388476
rect 71688 388424 71740 388476
rect 72332 388424 72384 388476
rect 128360 388424 128412 388476
rect 180616 388424 180668 388476
rect 184848 388424 184900 388476
rect 93952 388288 94004 388340
rect 94228 388288 94280 388340
rect 232596 387948 232648 388000
rect 236276 387948 236328 388000
rect 166264 387880 166316 387932
rect 167736 387880 167788 387932
rect 231216 387880 231268 387932
rect 234252 387880 234304 387932
rect 71688 387812 71740 387864
rect 72516 387812 72568 387864
rect 128360 387812 128412 387864
rect 129004 387812 129056 387864
rect 173624 387812 173676 387864
rect 196072 387812 196124 387864
rect 197268 387812 197320 387864
rect 221464 387812 221516 387864
rect 223948 387812 224000 387864
rect 233332 387812 233384 387864
rect 235264 387812 235316 387864
rect 249156 387812 249208 387864
rect 252284 387812 252336 387864
rect 103888 387744 103940 387796
rect 126244 387744 126296 387796
rect 187424 387744 187476 387796
rect 188436 387744 188488 387796
rect 188528 387744 188580 387796
rect 215944 387744 215996 387796
rect 238116 387744 238168 387796
rect 284300 387744 284352 387796
rect 184388 387676 184440 387728
rect 184848 387676 184900 387728
rect 202972 387676 203024 387728
rect 149704 387132 149756 387184
rect 168196 387132 168248 387184
rect 86868 387064 86920 387116
rect 106188 387064 106240 387116
rect 110420 387064 110472 387116
rect 187148 387064 187200 387116
rect 228364 387064 228416 387116
rect 253388 387064 253440 387116
rect 265716 387064 265768 387116
rect 582380 387064 582432 387116
rect 69020 386996 69072 387048
rect 69756 386996 69808 387048
rect 70400 386996 70452 387048
rect 71228 386996 71280 387048
rect 74540 386996 74592 387048
rect 75276 386996 75328 387048
rect 78680 386996 78732 387048
rect 79508 386996 79560 387048
rect 109040 386996 109092 387048
rect 109500 386996 109552 387048
rect 205640 386996 205692 387048
rect 206468 386996 206520 387048
rect 208400 386996 208452 387048
rect 209228 386996 209280 387048
rect 83188 386928 83240 386980
rect 84108 386928 84160 386980
rect 93952 386860 94004 386912
rect 94780 386860 94832 386912
rect 85120 386248 85172 386300
rect 124864 386316 124916 386368
rect 194140 386316 194192 386368
rect 252560 386316 252612 386368
rect 224868 386248 224920 386300
rect 258724 386248 258776 386300
rect 85396 385840 85448 385892
rect 88432 385840 88484 385892
rect 77208 385772 77260 385824
rect 78036 385772 78088 385824
rect 141976 385704 142028 385756
rect 147036 385704 147088 385756
rect 99564 385636 99616 385688
rect 170496 385636 170548 385688
rect 177396 385636 177448 385688
rect 180064 385636 180116 385688
rect 195888 385636 195940 385688
rect 267004 385636 267056 385688
rect 270500 385636 270552 385688
rect 188988 385364 189040 385416
rect 191196 385364 191248 385416
rect 158076 385024 158128 385076
rect 162124 385024 162176 385076
rect 185584 384956 185636 385008
rect 215300 384956 215352 385008
rect 239404 384956 239456 385008
rect 251732 384956 251784 385008
rect 251824 384956 251876 385008
rect 254032 384956 254084 385008
rect 192576 384888 192628 384940
rect 222844 384888 222896 384940
rect 226432 384344 226484 384396
rect 227628 384344 227680 384396
rect 73804 384276 73856 384328
rect 93124 384276 93176 384328
rect 215300 384276 215352 384328
rect 216036 384276 216088 384328
rect 106188 383732 106240 383784
rect 150440 383732 150492 383784
rect 3516 383664 3568 383716
rect 113456 383664 113508 383716
rect 150256 383664 150308 383716
rect 153936 383664 153988 383716
rect 227628 383664 227680 383716
rect 280160 383664 280212 383716
rect 109132 382984 109184 383036
rect 126244 382984 126296 383036
rect 175188 382984 175240 383036
rect 182088 382984 182140 383036
rect 208492 382984 208544 383036
rect 252468 382984 252520 383036
rect 263692 382984 263744 383036
rect 97724 382916 97776 382968
rect 124220 382916 124272 382968
rect 231860 382916 231912 382968
rect 281632 382916 281684 382968
rect 67364 382168 67416 382220
rect 150808 382168 150860 382220
rect 151084 382168 151136 382220
rect 177856 382168 177908 382220
rect 211160 382168 211212 382220
rect 102048 381488 102100 381540
rect 113364 381488 113416 381540
rect 150808 381488 150860 381540
rect 158720 381488 158772 381540
rect 173624 381488 173676 381540
rect 216680 381488 216732 381540
rect 227628 381488 227680 381540
rect 256792 381488 256844 381540
rect 211160 380876 211212 380928
rect 211804 380876 211856 380928
rect 231124 380876 231176 380928
rect 277676 380876 277728 380928
rect 48136 380808 48188 380860
rect 154028 380808 154080 380860
rect 236368 380808 236420 380860
rect 236644 380808 236696 380860
rect 281724 380808 281776 380860
rect 77300 380740 77352 380792
rect 130384 380740 130436 380792
rect 187700 380196 187752 380248
rect 226432 380196 226484 380248
rect 129740 380128 129792 380180
rect 138756 380128 138808 380180
rect 207020 380128 207072 380180
rect 221556 380128 221608 380180
rect 269396 380128 269448 380180
rect 270684 380128 270736 380180
rect 67272 379448 67324 379500
rect 157340 379448 157392 379500
rect 235264 379448 235316 379500
rect 235908 379448 235960 379500
rect 291292 379448 291344 379500
rect 157340 378972 157392 379024
rect 157984 378972 158036 379024
rect 188436 378836 188488 378888
rect 197452 378836 197504 378888
rect 121644 378768 121696 378820
rect 187700 378768 187752 378820
rect 241428 378768 241480 378820
rect 253940 378768 253992 378820
rect 111984 378088 112036 378140
rect 112444 378088 112496 378140
rect 179236 378020 179288 378072
rect 205732 378020 205784 378072
rect 227812 378088 227864 378140
rect 283196 378088 283248 378140
rect 228364 378020 228416 378072
rect 243084 378020 243136 378072
rect 262220 378020 262272 378072
rect 262864 378020 262916 378072
rect 97632 377408 97684 377460
rect 130384 377408 130436 377460
rect 94228 376660 94280 376712
rect 121644 376660 121696 376712
rect 148968 376660 149020 376712
rect 251272 376660 251324 376712
rect 108948 375980 109000 376032
rect 116124 375980 116176 376032
rect 88248 375300 88300 375352
rect 91928 375300 91980 375352
rect 213184 375300 213236 375352
rect 245752 375368 245804 375420
rect 263968 375368 264020 375420
rect 171968 375232 172020 375284
rect 218060 374008 218112 374060
rect 265164 374008 265216 374060
rect 82820 373940 82872 373992
rect 187148 373940 187200 373992
rect 250444 373940 250496 373992
rect 161572 373872 161624 373924
rect 162768 373872 162820 373924
rect 213920 373872 213972 373924
rect 187148 373396 187200 373448
rect 187608 373396 187660 373448
rect 107568 373260 107620 373312
rect 115940 373260 115992 373312
rect 242348 373260 242400 373312
rect 263784 373260 263836 373312
rect 137836 372716 137888 372768
rect 141516 372716 141568 372768
rect 61936 372512 61988 372564
rect 169760 372512 169812 372564
rect 188344 372512 188396 372564
rect 273260 372512 273312 372564
rect 93952 372444 94004 372496
rect 141240 372444 141292 372496
rect 141240 371832 141292 371884
rect 142068 371832 142120 371884
rect 178776 371832 178828 371884
rect 182824 371832 182876 371884
rect 187056 371832 187108 371884
rect 209044 371832 209096 371884
rect 234528 371832 234580 371884
rect 298100 371832 298152 371884
rect 169760 371220 169812 371272
rect 170404 371220 170456 371272
rect 67824 371152 67876 371204
rect 158076 371152 158128 371204
rect 161388 371152 161440 371204
rect 231216 371152 231268 371204
rect 150348 371084 150400 371136
rect 218060 371084 218112 371136
rect 232504 370472 232556 370524
rect 265256 370472 265308 370524
rect 101956 369792 102008 369844
rect 236644 369792 236696 369844
rect 110420 369724 110472 369776
rect 111064 369724 111116 369776
rect 148968 369724 149020 369776
rect 151176 369724 151228 369776
rect 255412 369724 255464 369776
rect 114468 368432 114520 368484
rect 281816 368432 281868 368484
rect 69112 368364 69164 368416
rect 165712 368364 165764 368416
rect 166356 368364 166408 368416
rect 168288 368364 168340 368416
rect 227720 368364 227772 368416
rect 228548 368364 228600 368416
rect 98368 367752 98420 367804
rect 113364 367752 113416 367804
rect 114468 367752 114520 367804
rect 228364 367752 228416 367804
rect 288440 367752 288492 367804
rect 67732 367004 67784 367056
rect 180800 367004 180852 367056
rect 181536 367004 181588 367056
rect 97264 366936 97316 366988
rect 161480 366936 161532 366988
rect 162216 366936 162268 366988
rect 183376 366324 183428 366376
rect 190552 366324 190604 366376
rect 218704 366324 218756 366376
rect 263600 366324 263652 366376
rect 93124 365644 93176 365696
rect 171232 365644 171284 365696
rect 171876 365644 171928 365696
rect 163872 365576 163924 365628
rect 221464 365576 221516 365628
rect 249708 365100 249760 365152
rect 252560 365100 252612 365152
rect 211804 364964 211856 365016
rect 256792 364964 256844 365016
rect 241520 364352 241572 364404
rect 249064 364352 249116 364404
rect 104716 364284 104768 364336
rect 60556 364216 60608 364268
rect 142988 364216 143040 364268
rect 153016 364216 153068 364268
rect 272156 364216 272208 364268
rect 123484 362856 123536 362908
rect 226340 362856 226392 362908
rect 240140 362244 240192 362296
rect 263600 362244 263652 362296
rect 93860 362176 93912 362228
rect 103520 362176 103572 362228
rect 212816 362176 212868 362228
rect 247776 362176 247828 362228
rect 226340 361564 226392 361616
rect 226984 361564 227036 361616
rect 155224 361496 155276 361548
rect 249156 361496 249208 361548
rect 249616 361496 249668 361548
rect 74632 361428 74684 361480
rect 156696 361428 156748 361480
rect 231216 360816 231268 360868
rect 253204 360816 253256 360868
rect 156052 360612 156104 360664
rect 156696 360612 156748 360664
rect 141608 360136 141660 360188
rect 255504 360136 255556 360188
rect 84108 360068 84160 360120
rect 155868 360068 155920 360120
rect 179512 360068 179564 360120
rect 179512 359660 179564 359712
rect 180156 359660 180208 359712
rect 255504 359660 255556 359712
rect 255964 359660 256016 359712
rect 195980 359456 196032 359508
rect 240140 359456 240192 359508
rect 69020 358708 69072 358760
rect 69664 358708 69716 358760
rect 142804 358708 142856 358760
rect 285864 358708 285916 358760
rect 194600 358640 194652 358692
rect 2780 358436 2832 358488
rect 4804 358436 4856 358488
rect 247776 358028 247828 358080
rect 253940 358028 253992 358080
rect 103428 356668 103480 356720
rect 110420 356668 110472 356720
rect 126244 356668 126296 356720
rect 155868 356668 155920 356720
rect 212816 356668 212868 356720
rect 242164 356668 242216 356720
rect 292580 356668 292632 356720
rect 110420 356056 110472 356108
rect 239404 356056 239456 356108
rect 75920 355988 75972 356040
rect 76564 355988 76616 356040
rect 202972 355988 203024 356040
rect 102232 355920 102284 355972
rect 103428 355920 103480 355972
rect 218796 355920 218848 355972
rect 222844 355308 222896 355360
rect 244924 355308 244976 355360
rect 249616 355308 249668 355360
rect 260380 355308 260432 355360
rect 137284 354628 137336 354680
rect 205640 354628 205692 354680
rect 100760 353948 100812 354000
rect 118792 353948 118844 354000
rect 236644 353948 236696 354000
rect 262404 353948 262456 354000
rect 118792 353268 118844 353320
rect 238116 353268 238168 353320
rect 74540 353200 74592 353252
rect 184296 353200 184348 353252
rect 205640 352588 205692 352640
rect 252836 352588 252888 352640
rect 108948 352520 109000 352572
rect 280344 352520 280396 352572
rect 119988 351840 120040 351892
rect 274824 351840 274876 351892
rect 172336 351160 172388 351212
rect 181444 351160 181496 351212
rect 204996 351160 205048 351212
rect 222936 351160 222988 351212
rect 180708 349868 180760 349920
rect 254584 349868 254636 349920
rect 107568 349800 107620 349852
rect 278872 349800 278924 349852
rect 130384 349052 130436 349104
rect 130660 349052 130712 349104
rect 231124 349052 231176 349104
rect 188988 348372 189040 348424
rect 253480 348372 253532 348424
rect 259368 347692 259420 347744
rect 261116 347692 261168 347744
rect 216036 347080 216088 347132
rect 261208 347080 261260 347132
rect 180156 347012 180208 347064
rect 242348 347012 242400 347064
rect 3148 346332 3200 346384
rect 42708 346332 42760 346384
rect 42708 345856 42760 345908
rect 43444 345856 43496 345908
rect 72516 345720 72568 345772
rect 73068 345720 73120 345772
rect 175556 345108 175608 345160
rect 198740 345108 198792 345160
rect 72516 345040 72568 345092
rect 231124 345040 231176 345092
rect 247684 344292 247736 344344
rect 251916 344292 251968 344344
rect 130384 343680 130436 343732
rect 228456 343680 228508 343732
rect 129096 343612 129148 343664
rect 129648 343612 129700 343664
rect 246488 343612 246540 343664
rect 209136 342864 209188 342916
rect 277400 342864 277452 342916
rect 175096 342320 175148 342372
rect 202144 342320 202196 342372
rect 95148 342252 95200 342304
rect 294052 342252 294104 342304
rect 143448 341572 143500 341624
rect 155408 341572 155460 341624
rect 177948 341572 178000 341624
rect 253296 341572 253348 341624
rect 101404 341504 101456 341556
rect 268016 341504 268068 341556
rect 183192 340144 183244 340196
rect 246396 340144 246448 340196
rect 67548 339464 67600 339516
rect 291476 339464 291528 339516
rect 239404 339396 239456 339448
rect 246304 339396 246356 339448
rect 215944 338784 215996 338836
rect 243544 338784 243596 338836
rect 33140 338716 33192 338768
rect 175096 338716 175148 338768
rect 191748 338716 191800 338768
rect 222200 338716 222252 338768
rect 246948 338716 247000 338768
rect 258080 338716 258132 338768
rect 148876 338104 148928 338156
rect 150440 338104 150492 338156
rect 215300 338104 215352 338156
rect 142804 337356 142856 337408
rect 188896 337356 188948 337408
rect 215576 337356 215628 337408
rect 221464 337356 221516 337408
rect 274640 337356 274692 337408
rect 141608 336744 141660 336796
rect 247776 336744 247828 336796
rect 165528 335996 165580 336048
rect 215484 335996 215536 336048
rect 244280 335792 244332 335844
rect 245016 335792 245068 335844
rect 143080 335316 143132 335368
rect 244280 335316 244332 335368
rect 222292 334636 222344 334688
rect 260840 334636 260892 334688
rect 151636 334568 151688 334620
rect 160192 334568 160244 334620
rect 177396 334568 177448 334620
rect 187516 334568 187568 334620
rect 242900 334568 242952 334620
rect 160192 333956 160244 334008
rect 160744 333956 160796 334008
rect 205640 333956 205692 334008
rect 205640 333276 205692 333328
rect 245752 333276 245804 333328
rect 246488 333276 246540 333328
rect 273536 333276 273588 333328
rect 30380 333208 30432 333260
rect 154028 333208 154080 333260
rect 172428 333208 172480 333260
rect 190368 333208 190420 333260
rect 247040 333208 247092 333260
rect 234620 332528 234672 332580
rect 240784 332528 240836 332580
rect 158076 331848 158128 331900
rect 173716 331848 173768 331900
rect 243176 331848 243228 331900
rect 148508 331236 148560 331288
rect 234620 331236 234672 331288
rect 94504 330488 94556 330540
rect 153200 330488 153252 330540
rect 172244 329876 172296 329928
rect 201592 329876 201644 329928
rect 166264 329808 166316 329860
rect 233884 329808 233936 329860
rect 252376 329740 252428 329792
rect 254032 329740 254084 329792
rect 164884 328516 164936 328568
rect 240140 328516 240192 328568
rect 116676 328448 116728 328500
rect 252376 328448 252428 328500
rect 218152 328380 218204 328432
rect 218704 328380 218756 328432
rect 260380 328380 260432 328432
rect 266728 328380 266780 328432
rect 209780 327700 209832 327752
rect 266360 327700 266412 327752
rect 190368 327156 190420 327208
rect 192484 327156 192536 327208
rect 121460 327088 121512 327140
rect 218152 327088 218204 327140
rect 123576 326340 123628 326392
rect 154488 326340 154540 326392
rect 160928 326340 160980 326392
rect 169392 326340 169444 326392
rect 241520 326340 241572 326392
rect 242256 326340 242308 326392
rect 256700 326340 256752 326392
rect 96712 325660 96764 325712
rect 250444 325660 250496 325712
rect 232596 324912 232648 324964
rect 271880 324912 271932 324964
rect 138664 324368 138716 324420
rect 209780 324368 209832 324420
rect 210240 324368 210292 324420
rect 41236 324300 41288 324352
rect 154488 324300 154540 324352
rect 175924 324300 175976 324352
rect 176476 324300 176528 324352
rect 258724 324300 258776 324352
rect 260840 323756 260892 323808
rect 261208 323756 261260 323808
rect 151176 323008 151228 323060
rect 260840 323008 260892 323060
rect 155316 322940 155368 322992
rect 269304 322940 269356 322992
rect 35900 322328 35952 322380
rect 153292 322328 153344 322380
rect 157064 322260 157116 322312
rect 233608 322260 233660 322312
rect 104808 322192 104860 322244
rect 277400 322192 277452 322244
rect 277768 322192 277820 322244
rect 153844 321580 153896 321632
rect 157064 321580 157116 321632
rect 154488 320832 154540 320884
rect 292580 320832 292632 320884
rect 185584 320152 185636 320204
rect 259736 320152 259788 320204
rect 84844 320084 84896 320136
rect 85488 320084 85540 320136
rect 150164 320084 150216 320136
rect 247132 320084 247184 320136
rect 4068 319404 4120 319456
rect 41236 319404 41288 319456
rect 252284 319404 252336 319456
rect 292672 319404 292724 319456
rect 188436 318792 188488 318844
rect 266636 318792 266688 318844
rect 44272 318044 44324 318096
rect 94504 318044 94556 318096
rect 178684 317500 178736 317552
rect 179328 317500 179380 317552
rect 249156 317500 249208 317552
rect 176016 317432 176068 317484
rect 266544 317432 266596 317484
rect 280252 317364 280304 317416
rect 280436 317364 280488 317416
rect 87604 316752 87656 316804
rect 88248 316752 88300 316804
rect 34428 316684 34480 316736
rect 165436 316684 165488 316736
rect 264980 316684 265032 316736
rect 87604 316004 87656 316056
rect 116584 316004 116636 316056
rect 148876 316004 148928 316056
rect 149796 316004 149848 316056
rect 188344 316004 188396 316056
rect 280436 316004 280488 316056
rect 155408 315460 155460 315512
rect 162216 315460 162268 315512
rect 154028 315324 154080 315376
rect 188436 315324 188488 315376
rect 40040 315256 40092 315308
rect 154120 315256 154172 315308
rect 231124 315256 231176 315308
rect 262864 315256 262916 315308
rect 170588 314712 170640 314764
rect 224224 314712 224276 314764
rect 187792 314644 187844 314696
rect 281540 314644 281592 314696
rect 281816 314644 281868 314696
rect 184204 313352 184256 313404
rect 240784 313352 240836 313404
rect 135996 313284 136048 313336
rect 260932 313284 260984 313336
rect 104164 312604 104216 312656
rect 116032 312604 116084 312656
rect 126888 312604 126940 312656
rect 92480 312536 92532 312588
rect 188344 312536 188396 312588
rect 187700 311924 187752 311976
rect 256884 311924 256936 311976
rect 126336 311856 126388 311908
rect 126888 311856 126940 311908
rect 263876 311856 263928 311908
rect 71044 311176 71096 311228
rect 77484 311176 77536 311228
rect 108212 311176 108264 311228
rect 118700 311176 118752 311228
rect 127624 311176 127676 311228
rect 67732 311108 67784 311160
rect 158720 311108 158772 311160
rect 259552 311108 259604 311160
rect 127624 310496 127676 310548
rect 251916 310496 251968 310548
rect 174728 309748 174780 309800
rect 187700 309748 187752 309800
rect 224868 309748 224920 309800
rect 255320 309748 255372 309800
rect 192484 309544 192536 309596
rect 198832 309544 198884 309596
rect 199384 309544 199436 309596
rect 116584 309136 116636 309188
rect 274916 309136 274968 309188
rect 52276 309068 52328 309120
rect 187700 309068 187752 309120
rect 97264 308388 97316 308440
rect 108212 308388 108264 308440
rect 147588 308388 147640 308440
rect 172520 308388 172572 308440
rect 188896 308388 188948 308440
rect 195244 308388 195296 308440
rect 230480 308388 230532 308440
rect 252744 308388 252796 308440
rect 111800 307776 111852 307828
rect 129096 307776 129148 307828
rect 172520 307776 172572 307828
rect 210056 307776 210108 307828
rect 242808 307776 242860 307828
rect 259460 307776 259512 307828
rect 202144 307708 202196 307760
rect 203984 307708 204036 307760
rect 282920 307708 282972 307760
rect 283104 307708 283156 307760
rect 99196 307096 99248 307148
rect 111800 307096 111852 307148
rect 93124 307028 93176 307080
rect 187792 307028 187844 307080
rect 235908 307028 235960 307080
rect 252560 307028 252612 307080
rect 115204 306416 115256 306468
rect 193864 306416 193916 306468
rect 188068 306348 188120 306400
rect 282920 306348 282972 306400
rect 3424 306280 3476 306332
rect 34428 306280 34480 306332
rect 262864 306144 262916 306196
rect 265072 306144 265124 306196
rect 224224 305668 224276 305720
rect 258080 305668 258132 305720
rect 76288 305600 76340 305652
rect 84844 305600 84896 305652
rect 92388 305600 92440 305652
rect 104164 305600 104216 305652
rect 104716 305600 104768 305652
rect 114652 305600 114704 305652
rect 195428 305600 195480 305652
rect 230388 305600 230440 305652
rect 242440 305600 242492 305652
rect 260104 305600 260156 305652
rect 276296 305600 276348 305652
rect 197360 305192 197412 305244
rect 198372 305192 198424 305244
rect 144736 305056 144788 305108
rect 197360 305056 197412 305108
rect 34428 304988 34480 305040
rect 35164 304988 35216 305040
rect 101496 304988 101548 305040
rect 102048 304988 102100 305040
rect 186320 304988 186372 305040
rect 187516 304988 187568 305040
rect 194416 304988 194468 305040
rect 227628 304716 227680 304768
rect 229192 304716 229244 304768
rect 246304 304648 246356 304700
rect 250168 304648 250220 304700
rect 230388 304308 230440 304360
rect 246580 304308 246632 304360
rect 97172 304240 97224 304292
rect 160192 304240 160244 304292
rect 213184 304240 213236 304292
rect 232780 304240 232832 304292
rect 249156 304240 249208 304292
rect 258172 304240 258224 304292
rect 259460 304240 259512 304292
rect 277584 304240 277636 304292
rect 290004 304240 290056 304292
rect 244740 304036 244792 304088
rect 246948 304036 247000 304088
rect 213828 303832 213880 303884
rect 222016 303832 222068 303884
rect 189816 303696 189868 303748
rect 195612 303696 195664 303748
rect 198740 303696 198792 303748
rect 201040 303696 201092 303748
rect 151084 303628 151136 303680
rect 212080 303628 212132 303680
rect 213920 303628 213972 303680
rect 214564 303628 214616 303680
rect 219440 303628 219492 303680
rect 219900 303628 219952 303680
rect 224960 303628 225012 303680
rect 225236 303628 225288 303680
rect 232228 303628 232280 303680
rect 233148 303628 233200 303680
rect 233884 303628 233936 303680
rect 234620 303628 234672 303680
rect 239404 303628 239456 303680
rect 242808 303628 242860 303680
rect 242900 303628 242952 303680
rect 243820 303628 243872 303680
rect 248420 303628 248472 303680
rect 249616 303628 249668 303680
rect 250812 303628 250864 303680
rect 262496 303628 262548 303680
rect 195980 303560 196032 303612
rect 196716 303560 196768 303612
rect 201500 303560 201552 303612
rect 201868 303560 201920 303612
rect 72700 302880 72752 302932
rect 175188 302880 175240 302932
rect 220820 302880 220872 302932
rect 232504 302880 232556 302932
rect 187700 302268 187752 302320
rect 218428 302268 218480 302320
rect 219348 302268 219400 302320
rect 240600 302268 240652 302320
rect 241428 302268 241480 302320
rect 268016 302268 268068 302320
rect 171784 302200 171836 302252
rect 172244 302200 172296 302252
rect 227444 302200 227496 302252
rect 240048 302200 240100 302252
rect 271972 302200 272024 302252
rect 186320 302132 186372 302184
rect 191472 302132 191524 302184
rect 228456 302132 228508 302184
rect 231032 302132 231084 302184
rect 92296 301520 92348 301572
rect 96620 301520 96672 301572
rect 250444 301520 250496 301572
rect 256792 301520 256844 301572
rect 94596 301452 94648 301504
rect 135996 301452 136048 301504
rect 193128 300908 193180 300960
rect 197636 300908 197688 300960
rect 175648 300840 175700 300892
rect 237380 300908 237432 300960
rect 238668 300908 238720 300960
rect 252376 300840 252428 300892
rect 252836 300840 252888 300892
rect 255596 300840 255648 300892
rect 255964 300840 256016 300892
rect 288624 300840 288676 300892
rect 170404 300772 170456 300824
rect 172244 300772 172296 300824
rect 183468 300772 183520 300824
rect 186964 300772 187016 300824
rect 259276 300160 259328 300212
rect 281540 300160 281592 300212
rect 169208 300092 169260 300144
rect 187700 300092 187752 300144
rect 262128 300092 262180 300144
rect 287060 300092 287112 300144
rect 303620 300092 303672 300144
rect 255504 300024 255556 300076
rect 259276 300024 259328 300076
rect 188344 299616 188396 299668
rect 193680 299616 193732 299668
rect 162216 299412 162268 299464
rect 185676 299412 185728 299464
rect 255504 299412 255556 299464
rect 262128 299412 262180 299464
rect 129188 298800 129240 298852
rect 159364 298800 159416 298852
rect 148324 298732 148376 298784
rect 187792 298732 187844 298784
rect 187608 298120 187660 298172
rect 191472 298120 191524 298172
rect 255504 298120 255556 298172
rect 271144 298120 271196 298172
rect 118700 297372 118752 297424
rect 175648 297372 175700 297424
rect 265624 297372 265676 297424
rect 296812 297372 296864 297424
rect 255504 296760 255556 296812
rect 263784 296760 263836 296812
rect 171140 296692 171192 296744
rect 191472 296692 191524 296744
rect 256056 296692 256108 296744
rect 276204 296692 276256 296744
rect 255504 296556 255556 296608
rect 259828 296556 259880 296608
rect 260748 296556 260800 296608
rect 86960 296012 87012 296064
rect 116676 296012 116728 296064
rect 117228 296012 117280 296064
rect 175924 296012 175976 296064
rect 67272 295944 67324 295996
rect 166448 295944 166500 295996
rect 174544 295944 174596 295996
rect 190000 295944 190052 295996
rect 253940 295604 253992 295656
rect 259460 295604 259512 295656
rect 260748 295332 260800 295384
rect 288440 295332 288492 295384
rect 255320 295264 255372 295316
rect 272156 295264 272208 295316
rect 156604 294652 156656 294704
rect 184848 294652 184900 294704
rect 186228 294652 186280 294704
rect 191472 294652 191524 294704
rect 65892 294584 65944 294636
rect 160100 294584 160152 294636
rect 163596 294584 163648 294636
rect 272156 294584 272208 294636
rect 285956 294584 286008 294636
rect 176200 293972 176252 294024
rect 178868 293972 178920 294024
rect 184848 293972 184900 294024
rect 186228 293972 186280 294024
rect 255412 293972 255464 294024
rect 298100 293972 298152 294024
rect 92572 293904 92624 293956
rect 93768 293904 93820 293956
rect 133788 293904 133840 293956
rect 133788 293224 133840 293276
rect 159364 293224 159416 293276
rect 171140 293292 171192 293344
rect 256700 293292 256752 293344
rect 289912 293292 289964 293344
rect 171784 293224 171836 293276
rect 187608 293224 187660 293276
rect 255412 293224 255464 293276
rect 259368 293224 259420 293276
rect 299480 293224 299532 293276
rect 3424 292544 3476 292596
rect 14464 292544 14516 292596
rect 82176 292544 82228 292596
rect 82636 292544 82688 292596
rect 113824 292544 113876 292596
rect 157248 292476 157300 292528
rect 164056 292476 164108 292528
rect 191472 292544 191524 292596
rect 176108 292408 176160 292460
rect 180064 292408 180116 292460
rect 191472 292408 191524 292460
rect 256608 291864 256660 291916
rect 263600 291864 263652 291916
rect 262864 291796 262916 291848
rect 280252 291796 280304 291848
rect 86224 291592 86276 291644
rect 93124 291592 93176 291644
rect 98276 291184 98328 291236
rect 99288 291184 99340 291236
rect 157248 291184 157300 291236
rect 67548 291116 67600 291168
rect 68560 291116 68612 291168
rect 131120 291116 131172 291168
rect 256516 291048 256568 291100
rect 260840 291048 260892 291100
rect 131120 290436 131172 290488
rect 132408 290436 132460 290488
rect 163688 290436 163740 290488
rect 261484 290436 261536 290488
rect 265072 290436 265124 290488
rect 186044 289960 186096 290012
rect 190828 289960 190880 290012
rect 170496 289892 170548 289944
rect 191472 289892 191524 289944
rect 84568 289824 84620 289876
rect 177396 289824 177448 289876
rect 256516 289824 256568 289876
rect 582564 289824 582616 289876
rect 256608 289756 256660 289808
rect 267740 289756 267792 289808
rect 71596 289144 71648 289196
rect 117228 289144 117280 289196
rect 164976 289144 165028 289196
rect 187608 289144 187660 289196
rect 78956 289076 79008 289128
rect 79968 289076 80020 289128
rect 159456 289076 159508 289128
rect 160008 289076 160060 289128
rect 191472 289076 191524 289128
rect 256516 289076 256568 289128
rect 259460 289076 259512 289128
rect 269304 289076 269356 289128
rect 56416 288396 56468 288448
rect 72516 288396 72568 288448
rect 72792 288396 72844 288448
rect 80060 288328 80112 288380
rect 80704 288328 80756 288380
rect 255872 288328 255924 288380
rect 277400 288328 277452 288380
rect 85856 287920 85908 287972
rect 86776 287920 86828 287972
rect 92480 287716 92532 287768
rect 92940 287716 92992 287768
rect 104624 287716 104676 287768
rect 115204 287716 115256 287768
rect 115296 287716 115348 287768
rect 169668 287716 169720 287768
rect 184756 287716 184808 287768
rect 191472 287716 191524 287768
rect 255964 287716 256016 287768
rect 259552 287716 259604 287768
rect 43444 287648 43496 287700
rect 70492 287648 70544 287700
rect 78588 287648 78640 287700
rect 184204 287648 184256 287700
rect 271144 287648 271196 287700
rect 284944 287648 284996 287700
rect 302240 287648 302292 287700
rect 73896 287036 73948 287088
rect 80060 287036 80112 287088
rect 86776 287036 86828 287088
rect 102140 287036 102192 287088
rect 91928 286968 91980 287020
rect 92388 286968 92440 287020
rect 142896 286968 142948 287020
rect 185584 286968 185636 287020
rect 255872 286968 255924 287020
rect 294052 286968 294104 287020
rect 95332 286696 95384 286748
rect 97264 286696 97316 286748
rect 52092 286288 52144 286340
rect 60648 286288 60700 286340
rect 74724 286356 74776 286408
rect 75736 286288 75788 286340
rect 142896 286288 142948 286340
rect 173624 286288 173676 286340
rect 186320 286288 186372 286340
rect 191472 286288 191524 286340
rect 82360 286220 82412 286272
rect 83464 286220 83516 286272
rect 91376 285880 91428 285932
rect 94596 285880 94648 285932
rect 187608 285880 187660 285932
rect 191380 285880 191432 285932
rect 60372 285676 60424 285728
rect 80980 285744 81032 285796
rect 80888 285676 80940 285728
rect 82176 285676 82228 285728
rect 84292 285676 84344 285728
rect 90364 285676 90416 285728
rect 163504 285676 163556 285728
rect 170588 285676 170640 285728
rect 256516 285676 256568 285728
rect 259736 285676 259788 285728
rect 263600 285676 263652 285728
rect 171048 285608 171100 285660
rect 189908 285608 189960 285660
rect 256608 285608 256660 285660
rect 263876 285608 263928 285660
rect 135996 284928 136048 284980
rect 148508 284928 148560 284980
rect 262220 284928 262272 284980
rect 291476 284928 291528 284980
rect 50988 284384 51040 284436
rect 69020 284384 69072 284436
rect 78220 284384 78272 284436
rect 100024 284384 100076 284436
rect 70308 284316 70360 284368
rect 99104 284316 99156 284368
rect 166356 284316 166408 284368
rect 191472 284316 191524 284368
rect 125600 284248 125652 284300
rect 156604 284248 156656 284300
rect 167644 284248 167696 284300
rect 193128 284248 193180 284300
rect 256424 284248 256476 284300
rect 266544 284248 266596 284300
rect 255780 283840 255832 283892
rect 258172 283840 258224 283892
rect 76150 283704 76202 283756
rect 76656 283704 76708 283756
rect 100944 283568 100996 283620
rect 125600 283568 125652 283620
rect 126428 283568 126480 283620
rect 137284 283568 137336 283620
rect 140136 283568 140188 283620
rect 148692 283568 148744 283620
rect 259276 283568 259328 283620
rect 273536 283568 273588 283620
rect 68836 283024 68888 283076
rect 69204 283024 69256 283076
rect 58992 282956 59044 283008
rect 70768 282956 70820 283008
rect 98736 282956 98788 283008
rect 99380 282888 99432 282940
rect 175924 282888 175976 282940
rect 178684 282888 178736 282940
rect 255504 282820 255556 282872
rect 271880 282820 271932 282872
rect 255412 282752 255464 282804
rect 264980 282752 265032 282804
rect 271880 282412 271932 282464
rect 273352 282412 273404 282464
rect 100760 281596 100812 281648
rect 115204 281596 115256 281648
rect 160836 281596 160888 281648
rect 191472 281596 191524 281648
rect 100852 281528 100904 281580
rect 189908 281528 189960 281580
rect 99380 281460 99432 281512
rect 140596 281460 140648 281512
rect 182824 281460 182876 281512
rect 255412 281460 255464 281512
rect 292580 281460 292632 281512
rect 255504 281392 255556 281444
rect 281724 281392 281776 281444
rect 126244 280848 126296 280900
rect 137468 280848 137520 280900
rect 137284 280780 137336 280832
rect 162124 280780 162176 280832
rect 163688 280780 163740 280832
rect 173808 280780 173860 280832
rect 176016 280780 176068 280832
rect 179236 280780 179288 280832
rect 191472 280780 191524 280832
rect 184296 280236 184348 280288
rect 191472 280236 191524 280288
rect 43444 280168 43496 280220
rect 67272 280168 67324 280220
rect 98736 280100 98788 280152
rect 176200 280100 176252 280152
rect 263968 280100 264020 280152
rect 264980 280100 265032 280152
rect 100760 280032 100812 280084
rect 155316 280032 155368 280084
rect 163596 280032 163648 280084
rect 164056 280032 164108 280084
rect 4068 279420 4120 279472
rect 52460 279420 52512 279472
rect 164056 279420 164108 279472
rect 191472 279420 191524 279472
rect 255412 279420 255464 279472
rect 259276 279420 259328 279472
rect 52460 278740 52512 278792
rect 53564 278740 53616 278792
rect 66812 278740 66864 278792
rect 53472 278672 53524 278724
rect 67548 278672 67600 278724
rect 255504 278672 255556 278724
rect 280160 278672 280212 278724
rect 258356 278604 258408 278656
rect 262404 278604 262456 278656
rect 100852 278060 100904 278112
rect 127716 278060 127768 278112
rect 105636 277992 105688 278044
rect 156052 277992 156104 278044
rect 183468 277992 183520 278044
rect 255412 277992 255464 278044
rect 258356 277992 258408 278044
rect 262864 277992 262916 278044
rect 291384 277992 291436 278044
rect 580172 277992 580224 278044
rect 67272 277924 67324 277976
rect 67548 277924 67600 277976
rect 183468 277380 183520 277432
rect 191472 277380 191524 277432
rect 52276 277312 52328 277364
rect 66904 277312 66956 277364
rect 100852 277312 100904 277364
rect 154028 277312 154080 277364
rect 255412 277312 255464 277364
rect 278872 277312 278924 277364
rect 100208 277244 100260 277296
rect 150532 277244 150584 277296
rect 151268 277244 151320 277296
rect 155316 276632 155368 276684
rect 177488 276632 177540 276684
rect 272340 276632 272392 276684
rect 281816 276632 281868 276684
rect 66168 276020 66220 276072
rect 67824 276020 67876 276072
rect 155500 276020 155552 276072
rect 190644 276020 190696 276072
rect 255504 276020 255556 276072
rect 271880 276020 271932 276072
rect 272340 276020 272392 276072
rect 255412 275952 255464 276004
rect 277676 275952 277728 276004
rect 255504 275612 255556 275664
rect 258080 275612 258132 275664
rect 155776 275340 155828 275392
rect 177396 275340 177448 275392
rect 56232 275272 56284 275324
rect 65708 275272 65760 275324
rect 66444 275272 66496 275324
rect 136548 275272 136600 275324
rect 184204 275272 184256 275324
rect 188436 275000 188488 275052
rect 191564 275000 191616 275052
rect 100944 274660 100996 274712
rect 152832 274660 152884 274712
rect 100852 274592 100904 274644
rect 120724 274592 120776 274644
rect 255504 274592 255556 274644
rect 281632 274592 281684 274644
rect 156604 273980 156656 274032
rect 188896 273980 188948 274032
rect 190828 273980 190880 274032
rect 100116 273912 100168 273964
rect 120172 273912 120224 273964
rect 124956 273912 125008 273964
rect 171784 273912 171836 273964
rect 255412 273912 255464 273964
rect 260932 273912 260984 273964
rect 56508 273300 56560 273352
rect 61108 273300 61160 273352
rect 64696 273232 64748 273284
rect 66628 273232 66680 273284
rect 172336 273164 172388 273216
rect 191564 273164 191616 273216
rect 255504 273164 255556 273216
rect 261484 273164 261536 273216
rect 157984 272552 158036 272604
rect 172336 272552 172388 272604
rect 48228 272484 48280 272536
rect 59084 272484 59136 272536
rect 100852 272484 100904 272536
rect 118056 272484 118108 272536
rect 174728 272484 174780 272536
rect 272064 272484 272116 272536
rect 281632 272484 281684 272536
rect 113180 271872 113232 271924
rect 180156 271804 180208 271856
rect 262404 271804 262456 271856
rect 267832 271804 267884 271856
rect 49516 271124 49568 271176
rect 65800 271124 65852 271176
rect 66536 271124 66588 271176
rect 147036 271124 147088 271176
rect 180800 271124 180852 271176
rect 181720 271124 181772 271176
rect 255412 270784 255464 270836
rect 259368 270784 259420 270836
rect 181720 270512 181772 270564
rect 191564 270512 191616 270564
rect 57612 270444 57664 270496
rect 57888 270444 57940 270496
rect 66812 270444 66864 270496
rect 100852 270444 100904 270496
rect 114560 270444 114612 270496
rect 119344 270444 119396 270496
rect 255412 270444 255464 270496
rect 280344 270444 280396 270496
rect 154028 269832 154080 269884
rect 169116 269832 169168 269884
rect 43996 269764 44048 269816
rect 57888 269764 57940 269816
rect 98828 269764 98880 269816
rect 165068 269764 165120 269816
rect 259368 269764 259420 269816
rect 280344 269764 280396 269816
rect 184204 269356 184256 269408
rect 191564 269356 191616 269408
rect 181996 269016 182048 269068
rect 191564 269016 191616 269068
rect 141424 268404 141476 268456
rect 181996 268404 182048 268456
rect 57796 268336 57848 268388
rect 59268 268336 59320 268388
rect 66812 268336 66864 268388
rect 104164 268336 104216 268388
rect 163504 268336 163556 268388
rect 168288 268336 168340 268388
rect 176660 268336 176712 268388
rect 269028 268336 269080 268388
rect 280436 268336 280488 268388
rect 104808 268200 104860 268252
rect 105544 268200 105596 268252
rect 255412 267792 255464 267844
rect 268108 267792 268160 267844
rect 269028 267792 269080 267844
rect 100852 267724 100904 267776
rect 104808 267724 104860 267776
rect 255504 267724 255556 267776
rect 269396 267724 269448 267776
rect 100024 267656 100076 267708
rect 135168 267656 135220 267708
rect 255412 267656 255464 267708
rect 267924 267656 267976 267708
rect 282920 267112 282972 267164
rect 284484 267112 284536 267164
rect 54944 267044 54996 267096
rect 65984 267044 66036 267096
rect 135168 267044 135220 267096
rect 169116 267044 169168 267096
rect 44088 266976 44140 267028
rect 58348 266976 58400 267028
rect 101404 266976 101456 267028
rect 141700 266976 141752 267028
rect 166448 266976 166500 267028
rect 174636 266976 174688 267028
rect 186136 266976 186188 267028
rect 192576 266976 192628 267028
rect 259368 266364 259420 266416
rect 282920 266364 282972 266416
rect 111800 266296 111852 266348
rect 113088 266296 113140 266348
rect 160836 266296 160888 266348
rect 168196 266296 168248 266348
rect 191656 266296 191708 266348
rect 255412 266160 255464 266212
rect 260104 266160 260156 266212
rect 101128 265616 101180 265668
rect 111800 265616 111852 265668
rect 153936 265616 153988 265668
rect 184940 265616 184992 265668
rect 190644 265616 190696 265668
rect 63132 264936 63184 264988
rect 66812 264936 66864 264988
rect 100852 264936 100904 264988
rect 133236 264936 133288 264988
rect 164976 264936 165028 264988
rect 168196 264936 168248 264988
rect 255320 264936 255372 264988
rect 295432 264936 295484 264988
rect 137468 264256 137520 264308
rect 169208 264256 169260 264308
rect 98736 264188 98788 264240
rect 153936 264188 153988 264240
rect 276020 264188 276072 264240
rect 285772 264188 285824 264240
rect 255412 264120 255464 264172
rect 259368 264120 259420 264172
rect 255504 263712 255556 263764
rect 259736 263712 259788 263764
rect 59268 263576 59320 263628
rect 63224 263576 63276 263628
rect 66628 263576 66680 263628
rect 100944 263576 100996 263628
rect 120724 263576 120776 263628
rect 160836 263576 160888 263628
rect 192024 263576 192076 263628
rect 260748 263576 260800 263628
rect 287244 263576 287296 263628
rect 100852 263508 100904 263560
rect 141608 263508 141660 263560
rect 142896 262964 142948 263016
rect 152740 262964 152792 263016
rect 152556 262896 152608 262948
rect 172520 262896 172572 262948
rect 54852 262828 54904 262880
rect 66260 262828 66312 262880
rect 141516 262828 141568 262880
rect 179420 262828 179472 262880
rect 255504 262284 255556 262336
rect 263876 262284 263928 262336
rect 22744 262216 22796 262268
rect 63224 262216 63276 262268
rect 66904 262216 66956 262268
rect 179420 262216 179472 262268
rect 191656 262216 191708 262268
rect 255412 262216 255464 262268
rect 267832 262216 267884 262268
rect 268292 262216 268344 262268
rect 164148 262148 164200 262200
rect 168380 262148 168432 262200
rect 104808 262080 104860 262132
rect 111064 262080 111116 262132
rect 7564 261468 7616 261520
rect 67088 261468 67140 261520
rect 100852 261468 100904 261520
rect 104624 261468 104676 261520
rect 134616 261468 134668 261520
rect 141516 261468 141568 261520
rect 167092 261468 167144 261520
rect 255504 261468 255556 261520
rect 276020 261468 276072 261520
rect 255412 261332 255464 261384
rect 259368 261332 259420 261384
rect 168380 260856 168432 260908
rect 191656 260856 191708 260908
rect 255412 260448 255464 260500
rect 260748 260448 260800 260500
rect 169300 260176 169352 260228
rect 191380 260176 191432 260228
rect 55036 260108 55088 260160
rect 66260 260108 66312 260160
rect 129280 260108 129332 260160
rect 170496 260108 170548 260160
rect 259368 260108 259420 260160
rect 278964 260108 279016 260160
rect 48228 259428 48280 259480
rect 67732 259428 67784 259480
rect 100852 259428 100904 259480
rect 149888 259428 149940 259480
rect 176660 259428 176712 259480
rect 191656 259428 191708 259480
rect 285772 259428 285824 259480
rect 287336 259428 287388 259480
rect 64604 259360 64656 259412
rect 66812 259360 66864 259412
rect 255412 259360 255464 259412
rect 265164 259360 265216 259412
rect 273904 259360 273956 259412
rect 274732 259360 274784 259412
rect 186320 259088 186372 259140
rect 187148 259088 187200 259140
rect 52184 258680 52236 258732
rect 61752 258680 61804 258732
rect 66260 258680 66312 258732
rect 98368 258136 98420 258188
rect 113916 258136 113968 258188
rect 171140 258136 171192 258188
rect 190460 258136 190512 258188
rect 108488 258068 108540 258120
rect 187148 258068 187200 258120
rect 66260 258000 66312 258052
rect 68192 258000 68244 258052
rect 255412 258000 255464 258052
rect 261484 258000 261536 258052
rect 39856 257320 39908 257372
rect 52460 257320 52512 257372
rect 101956 257320 102008 257372
rect 112720 257320 112772 257372
rect 169024 257320 169076 257372
rect 185492 257320 185544 257372
rect 255320 257320 255372 257372
rect 256976 257320 257028 257372
rect 259552 257320 259604 257372
rect 580908 257320 580960 257372
rect 185584 257184 185636 257236
rect 190644 257184 190696 257236
rect 52460 256708 52512 256760
rect 53472 256708 53524 256760
rect 66260 256708 66312 256760
rect 125048 256708 125100 256760
rect 187056 256708 187108 256760
rect 100852 256640 100904 256692
rect 143080 256640 143132 256692
rect 180248 256164 180300 256216
rect 182824 256164 182876 256216
rect 166908 256028 166960 256080
rect 173900 256028 173952 256080
rect 50896 255960 50948 256012
rect 56508 255960 56560 256012
rect 147036 255960 147088 256012
rect 170404 255960 170456 256012
rect 175188 255960 175240 256012
rect 191656 255960 191708 256012
rect 255504 255348 255556 255400
rect 265072 255348 265124 255400
rect 100944 255280 100996 255332
rect 148508 255280 148560 255332
rect 255412 255280 255464 255332
rect 274916 255280 274968 255332
rect 3424 255212 3476 255264
rect 43444 255212 43496 255264
rect 100852 255212 100904 255264
rect 108948 255212 109000 255264
rect 177764 255212 177816 255264
rect 191012 255212 191064 255264
rect 114652 255144 114704 255196
rect 272340 254600 272392 254652
rect 283196 254600 283248 254652
rect 48136 254532 48188 254584
rect 66812 254532 66864 254584
rect 120724 254532 120776 254584
rect 184388 254532 184440 254584
rect 255412 254532 255464 254584
rect 285772 254532 285824 254584
rect 108396 253920 108448 253972
rect 109684 253920 109736 253972
rect 109868 253920 109920 253972
rect 112444 253920 112496 253972
rect 255504 253920 255556 253972
rect 272064 253920 272116 253972
rect 272340 253920 272392 253972
rect 111800 253240 111852 253292
rect 147128 253240 147180 253292
rect 35164 253172 35216 253224
rect 66996 253172 67048 253224
rect 67272 253172 67324 253224
rect 116676 253172 116728 253224
rect 176016 253172 176068 253224
rect 188896 252968 188948 253020
rect 189724 252968 189776 253020
rect 279332 252764 279384 252816
rect 284392 252764 284444 252816
rect 255412 252696 255464 252748
rect 258264 252696 258316 252748
rect 100852 252560 100904 252612
rect 109684 252560 109736 252612
rect 163504 252560 163556 252612
rect 188896 252560 188948 252612
rect 255504 252560 255556 252612
rect 283104 252560 283156 252612
rect 186044 252492 186096 252544
rect 191104 252492 191156 252544
rect 166264 251880 166316 251932
rect 191012 251880 191064 251932
rect 54760 251812 54812 251864
rect 63500 251812 63552 251864
rect 132040 251812 132092 251864
rect 166356 251812 166408 251864
rect 255412 251812 255464 251864
rect 278872 251812 278924 251864
rect 279332 251812 279384 251864
rect 291108 251812 291160 251864
rect 299572 251812 299624 251864
rect 104256 251744 104308 251796
rect 104808 251744 104860 251796
rect 63500 251268 63552 251320
rect 64696 251268 64748 251320
rect 66812 251268 66864 251320
rect 257988 251268 258040 251320
rect 259552 251268 259604 251320
rect 104808 251200 104860 251252
rect 131120 251200 131172 251252
rect 132040 251200 132092 251252
rect 255320 251200 255372 251252
rect 291108 251200 291160 251252
rect 98736 251132 98788 251184
rect 103428 251132 103480 251184
rect 128360 251132 128412 251184
rect 129280 251132 129332 251184
rect 262496 251132 262548 251184
rect 262864 251132 262916 251184
rect 269028 251132 269080 251184
rect 582656 251132 582708 251184
rect 100852 251064 100904 251116
rect 107568 251064 107620 251116
rect 111064 251064 111116 251116
rect 58992 250520 59044 250572
rect 66812 250520 66864 250572
rect 146116 250520 146168 250572
rect 158720 250520 158772 250572
rect 186320 250520 186372 250572
rect 191656 250520 191708 250572
rect 255412 250520 255464 250572
rect 262496 250520 262548 250572
rect 115296 250452 115348 250504
rect 174728 250452 174780 250504
rect 255504 250452 255556 250504
rect 267924 250452 267976 250504
rect 269028 250452 269080 250504
rect 187148 249908 187200 249960
rect 192668 249908 192720 249960
rect 100852 249704 100904 249756
rect 109868 249704 109920 249756
rect 254216 249364 254268 249416
rect 257988 249364 258040 249416
rect 259552 249364 259604 249416
rect 53656 249024 53708 249076
rect 60648 249024 60700 249076
rect 66444 249024 66496 249076
rect 109868 249024 109920 249076
rect 130568 249024 130620 249076
rect 155500 249024 155552 249076
rect 166356 249024 166408 249076
rect 176108 249024 176160 249076
rect 187148 248412 187200 248464
rect 191012 248412 191064 248464
rect 255412 248412 255464 248464
rect 278044 248412 278096 248464
rect 112536 247732 112588 247784
rect 171784 247732 171836 247784
rect 107016 247664 107068 247716
rect 179512 247664 179564 247716
rect 255412 247664 255464 247716
rect 265072 247664 265124 247716
rect 187608 247460 187660 247512
rect 190460 247460 190512 247512
rect 62028 247052 62080 247104
rect 66812 247052 66864 247104
rect 179512 247052 179564 247104
rect 182916 247052 182968 247104
rect 186964 247052 187016 247104
rect 191748 247052 191800 247104
rect 255504 247052 255556 247104
rect 265716 247052 265768 247104
rect 269212 247052 269264 247104
rect 100668 246984 100720 247036
rect 124956 246984 125008 247036
rect 190368 246372 190420 246424
rect 193404 246372 193456 246424
rect 99380 246304 99432 246356
rect 191196 246304 191248 246356
rect 281448 246304 281500 246356
rect 298284 246304 298336 246356
rect 98644 245624 98696 245676
rect 99380 245624 99432 245676
rect 125140 245624 125192 245676
rect 161480 245624 161532 245676
rect 162676 245624 162728 245676
rect 255504 245624 255556 245676
rect 280804 245624 280856 245676
rect 281448 245624 281500 245676
rect 101036 245556 101088 245608
rect 155960 245556 156012 245608
rect 255412 245556 255464 245608
rect 289820 245556 289872 245608
rect 100852 245488 100904 245540
rect 108396 245488 108448 245540
rect 138848 245488 138900 245540
rect 187700 245488 187752 245540
rect 155960 244876 156012 244928
rect 193496 244876 193548 244928
rect 255412 244264 255464 244316
rect 270408 244264 270460 244316
rect 289820 244264 289872 244316
rect 293960 244264 294012 244316
rect 255872 244196 255924 244248
rect 285680 244196 285732 244248
rect 111156 243516 111208 243568
rect 151176 243516 151228 243568
rect 183468 243516 183520 243568
rect 192484 243516 192536 243568
rect 255504 243516 255556 243568
rect 277492 243516 277544 243568
rect 157340 243312 157392 243364
rect 158168 243312 158220 243364
rect 100852 242972 100904 243024
rect 102784 242972 102836 243024
rect 52368 242904 52420 242956
rect 66720 242904 66772 242956
rect 67640 242904 67692 242956
rect 68468 242904 68520 242956
rect 102876 242904 102928 242956
rect 157340 242904 157392 242956
rect 182088 242904 182140 242956
rect 184296 242904 184348 242956
rect 3424 242156 3476 242208
rect 22744 242156 22796 242208
rect 109776 242156 109828 242208
rect 178868 242156 178920 242208
rect 100852 242088 100904 242140
rect 103612 242088 103664 242140
rect 261024 242156 261076 242208
rect 249156 242020 249208 242072
rect 249800 242020 249852 242072
rect 253020 242020 253072 242072
rect 162308 241952 162360 242004
rect 162768 241952 162820 242004
rect 186320 241544 186372 241596
rect 191748 241544 191800 241596
rect 191840 241544 191892 241596
rect 213276 241544 213328 241596
rect 53748 241476 53800 241528
rect 66812 241476 66864 241528
rect 98414 241476 98466 241528
rect 103428 241476 103480 241528
rect 106280 241476 106332 241528
rect 162308 241476 162360 241528
rect 197176 241476 197228 241528
rect 14464 241408 14516 241460
rect 93124 241408 93176 241460
rect 93446 241408 93498 241460
rect 95654 241408 95706 241460
rect 110420 241408 110472 241460
rect 174728 241408 174780 241460
rect 259460 241408 259512 241460
rect 73528 241340 73580 241392
rect 105636 241340 105688 241392
rect 269764 241000 269816 241052
rect 273444 241000 273496 241052
rect 152832 240728 152884 240780
rect 180248 240728 180300 240780
rect 192668 240728 192720 240780
rect 209044 240728 209096 240780
rect 244924 240728 244976 240780
rect 263784 240728 263836 240780
rect 69480 240252 69532 240304
rect 74540 240116 74592 240168
rect 74908 240116 74960 240168
rect 82820 240116 82872 240168
rect 83740 240116 83792 240168
rect 84200 240116 84252 240168
rect 84844 240116 84896 240168
rect 86960 240116 87012 240168
rect 87604 240116 87656 240168
rect 165712 240048 165764 240100
rect 169024 240048 169076 240100
rect 69020 239980 69072 240032
rect 69940 239980 69992 240032
rect 70492 239980 70544 240032
rect 71320 239980 71372 240032
rect 95148 239980 95200 240032
rect 98736 239980 98788 240032
rect 103428 239980 103480 240032
rect 183376 240048 183428 240100
rect 195244 240048 195296 240100
rect 213276 240048 213328 240100
rect 230756 240048 230808 240100
rect 237656 240048 237708 240100
rect 251824 240048 251876 240100
rect 252284 240048 252336 240100
rect 283012 240048 283064 240100
rect 222200 239980 222252 240032
rect 223488 239980 223540 240032
rect 80060 239776 80112 239828
rect 80980 239776 81032 239828
rect 224868 239572 224920 239624
rect 225972 239572 226024 239624
rect 89352 239436 89404 239488
rect 91928 239436 91980 239488
rect 56416 239368 56468 239420
rect 71044 239368 71096 239420
rect 169024 239368 169076 239420
rect 209136 239368 209188 239420
rect 237380 239368 237432 239420
rect 256884 239368 256936 239420
rect 258816 239368 258868 239420
rect 270776 239368 270828 239420
rect 247040 238756 247092 238808
rect 252468 238756 252520 238808
rect 67824 238688 67876 238740
rect 102876 238688 102928 238740
rect 180064 238688 180116 238740
rect 213920 238688 213972 238740
rect 221096 238688 221148 238740
rect 273904 238688 273956 238740
rect 193588 238620 193640 238672
rect 215300 238620 215352 238672
rect 242716 238620 242768 238672
rect 274640 238620 274692 238672
rect 215300 238348 215352 238400
rect 216312 238348 216364 238400
rect 106280 238076 106332 238128
rect 173256 238076 173308 238128
rect 96896 238008 96948 238060
rect 108396 238008 108448 238060
rect 110420 238008 110472 238060
rect 180800 238008 180852 238060
rect 213920 237396 213972 237448
rect 214656 237396 214708 237448
rect 242256 237396 242308 237448
rect 242716 237396 242768 237448
rect 92572 237328 92624 237380
rect 125048 237328 125100 237380
rect 169760 237328 169812 237380
rect 189724 237328 189776 237380
rect 193680 237328 193732 237380
rect 237932 237328 237984 237380
rect 177396 237260 177448 237312
rect 201500 237260 201552 237312
rect 201960 237260 202012 237312
rect 74448 236648 74500 236700
rect 77300 236648 77352 236700
rect 207664 236648 207716 236700
rect 221096 236648 221148 236700
rect 242164 236648 242216 236700
rect 266452 236648 266504 236700
rect 89628 236444 89680 236496
rect 91100 236444 91152 236496
rect 91100 236308 91152 236360
rect 94780 236308 94832 236360
rect 77668 236172 77720 236224
rect 83556 236172 83608 236224
rect 91192 235968 91244 236020
rect 94688 235968 94740 236020
rect 95240 235968 95292 236020
rect 237472 235968 237524 236020
rect 237932 235968 237984 236020
rect 124312 235900 124364 235952
rect 192576 235900 192628 235952
rect 205732 235900 205784 235952
rect 205732 235424 205784 235476
rect 206744 235424 206796 235476
rect 193128 235288 193180 235340
rect 220820 235288 220872 235340
rect 222844 235288 222896 235340
rect 252744 235288 252796 235340
rect 213184 235220 213236 235272
rect 255504 235220 255556 235272
rect 582656 235220 582708 235272
rect 82084 234540 82136 234592
rect 108488 234540 108540 234592
rect 185584 234540 185636 234592
rect 256976 234540 257028 234592
rect 67732 233996 67784 234048
rect 71780 233996 71832 234048
rect 97908 233860 97960 233912
rect 99472 233860 99524 233912
rect 177396 233860 177448 233912
rect 259736 233860 259788 233912
rect 290464 233656 290516 233708
rect 291108 233656 291160 233708
rect 291108 233248 291160 233300
rect 580264 233248 580316 233300
rect 80336 233180 80388 233232
rect 161480 233180 161532 233232
rect 162308 233180 162360 233232
rect 174636 233180 174688 233232
rect 175188 233180 175240 233232
rect 259644 233180 259696 233232
rect 278044 233180 278096 233232
rect 281816 233180 281868 233232
rect 117964 233112 118016 233164
rect 121644 233112 121696 233164
rect 267004 232568 267056 232620
rect 276296 232568 276348 232620
rect 88340 232500 88392 232552
rect 117964 232500 118016 232552
rect 133236 232500 133288 232552
rect 210424 232500 210476 232552
rect 239404 232500 239456 232552
rect 274916 232500 274968 232552
rect 281816 231820 281868 231872
rect 580172 231820 580224 231872
rect 79968 231140 80020 231192
rect 87604 231140 87656 231192
rect 89720 231140 89772 231192
rect 124128 231140 124180 231192
rect 130660 231140 130712 231192
rect 153936 231140 153988 231192
rect 215944 231140 215996 231192
rect 60372 231072 60424 231124
rect 79324 231072 79376 231124
rect 84200 231072 84252 231124
rect 114744 231072 114796 231124
rect 182548 231072 182600 231124
rect 235264 231072 235316 231124
rect 255688 231072 255740 231124
rect 257344 231072 257396 231124
rect 278964 231072 279016 231124
rect 179236 230392 179288 230444
rect 215392 230392 215444 230444
rect 63224 229712 63276 229764
rect 75920 229712 75972 229764
rect 184756 229712 184808 229764
rect 203524 229712 203576 229764
rect 3424 229168 3476 229220
rect 96988 229168 97040 229220
rect 75920 229100 75972 229152
rect 175924 229100 175976 229152
rect 107568 229032 107620 229084
rect 280344 229032 280396 229084
rect 191196 228964 191248 229016
rect 253204 228964 253256 229016
rect 106924 228692 106976 228744
rect 107568 228692 107620 228744
rect 80060 228352 80112 228404
rect 106372 228352 106424 228404
rect 111156 228352 111208 228404
rect 96528 227740 96580 227792
rect 100852 227740 100904 227792
rect 252744 227740 252796 227792
rect 253204 227740 253256 227792
rect 149888 227672 149940 227724
rect 262404 227672 262456 227724
rect 158168 227604 158220 227656
rect 204352 227604 204404 227656
rect 78588 226992 78640 227044
rect 111156 226992 111208 227044
rect 118056 226992 118108 227044
rect 158168 226312 158220 226364
rect 158628 226312 158680 226364
rect 108304 225632 108356 225684
rect 122104 225632 122156 225684
rect 184388 225632 184440 225684
rect 244280 225632 244332 225684
rect 109684 225564 109736 225616
rect 245660 225564 245712 225616
rect 265072 225564 265124 225616
rect 244280 224884 244332 224936
rect 245016 224884 245068 224936
rect 272064 224884 272116 224936
rect 91376 224272 91428 224324
rect 182916 224272 182968 224324
rect 178868 224204 178920 224256
rect 219440 224204 219492 224256
rect 281724 224204 281776 224256
rect 196716 223524 196768 223576
rect 197268 223524 197320 223576
rect 269304 223524 269356 223576
rect 102784 222844 102836 222896
rect 204904 222844 204956 222896
rect 214564 222844 214616 222896
rect 255596 222844 255648 222896
rect 87052 222096 87104 222148
rect 116032 222096 116084 222148
rect 116584 222096 116636 222148
rect 112628 221416 112680 221468
rect 270592 221416 270644 221468
rect 98000 220736 98052 220788
rect 98920 220736 98972 220788
rect 215944 220736 215996 220788
rect 292672 220736 292724 220788
rect 59176 220124 59228 220176
rect 159548 220124 159600 220176
rect 98920 219988 98972 220040
rect 266360 220056 266412 220108
rect 159548 219376 159600 219428
rect 258816 219376 258868 219428
rect 213276 219308 213328 219360
rect 285956 219308 286008 219360
rect 285680 218764 285732 218816
rect 285956 218764 286008 218816
rect 82820 218696 82872 218748
rect 180064 218696 180116 218748
rect 213184 218696 213236 218748
rect 182916 217948 182968 218000
rect 246304 217948 246356 218000
rect 155408 217268 155460 217320
rect 247040 217268 247092 217320
rect 285128 217268 285180 217320
rect 295524 217268 295576 217320
rect 74540 217132 74592 217184
rect 75644 217132 75696 217184
rect 75644 216656 75696 216708
rect 172336 216656 172388 216708
rect 137560 215976 137612 216028
rect 220084 215976 220136 216028
rect 256056 215976 256108 216028
rect 268016 215976 268068 216028
rect 86960 215908 87012 215960
rect 88248 215908 88300 215960
rect 262220 215908 262272 215960
rect 156696 215228 156748 215280
rect 281816 215228 281868 215280
rect 3516 214888 3568 214940
rect 7564 214888 7616 214940
rect 169760 214548 169812 214600
rect 257344 214548 257396 214600
rect 93124 213868 93176 213920
rect 95700 213868 95752 213920
rect 149796 213868 149848 213920
rect 169760 213868 169812 213920
rect 182824 213868 182876 213920
rect 183468 213868 183520 213920
rect 239404 213868 239456 213920
rect 95240 212508 95292 212560
rect 95700 212508 95752 212560
rect 273352 212508 273404 212560
rect 103612 212440 103664 212492
rect 264980 212440 265032 212492
rect 108396 211760 108448 211812
rect 270500 211760 270552 211812
rect 98828 211148 98880 211200
rect 103612 211148 103664 211200
rect 50896 211080 50948 211132
rect 167000 211080 167052 211132
rect 249800 211080 249852 211132
rect 138020 211012 138072 211064
rect 138756 211012 138808 211064
rect 177396 211012 177448 211064
rect 59176 209040 59228 209092
rect 69020 209040 69072 209092
rect 176568 208292 176620 208344
rect 290464 208292 290516 208344
rect 176016 207816 176068 207868
rect 176568 207816 176620 207868
rect 97264 207000 97316 207052
rect 102232 207000 102284 207052
rect 263692 207000 263744 207052
rect 265072 206932 265124 206984
rect 265716 206932 265768 206984
rect 579804 206932 579856 206984
rect 93860 206320 93912 206372
rect 104992 206320 105044 206372
rect 105728 206320 105780 206372
rect 95884 206252 95936 206304
rect 256700 206252 256752 206304
rect 95332 205980 95384 206032
rect 95884 205980 95936 206032
rect 105728 205640 105780 205692
rect 258080 205640 258132 205692
rect 258356 205640 258408 205692
rect 96620 204892 96672 204944
rect 111892 204892 111944 204944
rect 274640 204688 274692 204740
rect 274824 204688 274876 204740
rect 111892 204280 111944 204332
rect 274640 204280 274692 204332
rect 191104 204212 191156 204264
rect 193312 204212 193364 204264
rect 188988 203532 189040 203584
rect 195980 203532 196032 203584
rect 98000 202784 98052 202836
rect 98920 202784 98972 202836
rect 180156 202172 180208 202224
rect 196624 202172 196676 202224
rect 3516 202104 3568 202156
rect 98000 202104 98052 202156
rect 195888 202104 195940 202156
rect 253940 202104 253992 202156
rect 260196 200812 260248 200864
rect 271972 200812 272024 200864
rect 44088 200744 44140 200796
rect 134708 200744 134760 200796
rect 149796 200744 149848 200796
rect 188344 200744 188396 200796
rect 200028 200744 200080 200796
rect 582472 200744 582524 200796
rect 53472 200064 53524 200116
rect 291384 200064 291436 200116
rect 53472 198704 53524 198756
rect 53656 198704 53708 198756
rect 31760 197956 31812 198008
rect 186964 197956 187016 198008
rect 255228 197956 255280 198008
rect 280252 197956 280304 198008
rect 37280 196596 37332 196648
rect 152648 196596 152700 196648
rect 123484 195304 123536 195356
rect 140044 195304 140096 195356
rect 261484 195304 261536 195356
rect 276204 195304 276256 195356
rect 97816 195236 97868 195288
rect 123576 195236 123628 195288
rect 197360 195236 197412 195288
rect 283104 195236 283156 195288
rect 108304 193808 108356 193860
rect 129188 193808 129240 193860
rect 131764 193808 131816 193860
rect 147036 193808 147088 193860
rect 148508 193808 148560 193860
rect 162216 193808 162268 193860
rect 251916 192516 251968 192568
rect 277584 192516 277636 192568
rect 187608 192448 187660 192500
rect 228364 192448 228416 192500
rect 255964 192448 256016 192500
rect 256608 192448 256660 192500
rect 580172 192448 580224 192500
rect 222936 191088 222988 191140
rect 260932 191088 260984 191140
rect 80704 189728 80756 189780
rect 145564 189728 145616 189780
rect 195244 189728 195296 189780
rect 226616 189728 226668 189780
rect 61752 188300 61804 188352
rect 71780 188300 71832 188352
rect 81348 188300 81400 188352
rect 103520 188300 103572 188352
rect 114560 188300 114612 188352
rect 131856 188300 131908 188352
rect 137376 188300 137428 188352
rect 148416 188300 148468 188352
rect 175924 188300 175976 188352
rect 185676 188300 185728 188352
rect 195796 188300 195848 188352
rect 298100 188300 298152 188352
rect 145564 188096 145616 188148
rect 154028 188096 154080 188148
rect 193128 187008 193180 187060
rect 234620 187008 234672 187060
rect 9680 186940 9732 186992
rect 186320 186940 186372 186992
rect 228364 186940 228416 186992
rect 278872 186940 278924 186992
rect 202144 185580 202196 185632
rect 243544 185580 243596 185632
rect 79324 184900 79376 184952
rect 204260 184900 204312 184952
rect 73160 184220 73212 184272
rect 91744 184220 91796 184272
rect 118792 184220 118844 184272
rect 137468 184220 137520 184272
rect 89628 184152 89680 184204
rect 126520 184152 126572 184204
rect 180156 184152 180208 184204
rect 190460 184152 190512 184204
rect 196716 184152 196768 184204
rect 218704 184152 218756 184204
rect 33784 182792 33836 182844
rect 140136 182792 140188 182844
rect 86868 181500 86920 181552
rect 117320 181500 117372 181552
rect 140044 181500 140096 181552
rect 145656 181500 145708 181552
rect 63132 181432 63184 181484
rect 180156 181432 180208 181484
rect 207756 181432 207808 181484
rect 288532 181432 288584 181484
rect 88432 180072 88484 180124
rect 116124 180072 116176 180124
rect 203524 180072 203576 180124
rect 240232 180072 240284 180124
rect 52184 179392 52236 179444
rect 167736 179392 167788 179444
rect 172428 179392 172480 179444
rect 202880 179392 202932 179444
rect 87604 178644 87656 178696
rect 105084 178644 105136 178696
rect 106924 178644 106976 178696
rect 142988 178644 143040 178696
rect 182824 178644 182876 178696
rect 227720 178644 227772 178696
rect 247684 178644 247736 178696
rect 248328 178644 248380 178696
rect 580172 178644 580224 178696
rect 243544 178304 243596 178356
rect 249892 178304 249944 178356
rect 190368 177284 190420 177336
rect 274732 177284 274784 177336
rect 195980 175312 196032 175364
rect 213184 175312 213236 175364
rect 113824 175244 113876 175296
rect 204904 175244 204956 175296
rect 248972 175244 249024 175296
rect 583024 175244 583076 175296
rect 150532 175176 150584 175228
rect 195980 175176 196032 175228
rect 88340 174496 88392 174548
rect 150532 174496 150584 174548
rect 154028 173884 154080 173936
rect 220820 173884 220872 173936
rect 221464 173884 221516 173936
rect 222292 173816 222344 173868
rect 222936 173816 222988 173868
rect 57704 173136 57756 173188
rect 201592 173136 201644 173188
rect 202144 173136 202196 173188
rect 227996 173136 228048 173188
rect 251824 173136 251876 173188
rect 341524 173136 341576 173188
rect 87144 172524 87196 172576
rect 222292 172524 222344 172576
rect 205824 172456 205876 172508
rect 303620 172456 303672 172508
rect 304080 172456 304132 172508
rect 304080 171776 304132 171828
rect 320180 171776 320232 171828
rect 92664 171096 92716 171148
rect 222844 171096 222896 171148
rect 91192 170348 91244 170400
rect 154028 170348 154080 170400
rect 154396 169804 154448 169856
rect 86224 169736 86276 169788
rect 213920 169736 213972 169788
rect 214564 169736 214616 169788
rect 216864 169736 216916 169788
rect 217968 169736 218020 169788
rect 582748 169736 582800 169788
rect 134708 168444 134760 168496
rect 227996 168444 228048 168496
rect 73344 168376 73396 168428
rect 200304 168308 200356 168360
rect 254032 168308 254084 168360
rect 67732 167016 67784 167068
rect 68928 167016 68980 167068
rect 192576 167084 192628 167136
rect 101404 167016 101456 167068
rect 101588 167016 101640 167068
rect 233240 167016 233292 167068
rect 63224 166268 63276 166320
rect 164056 166268 164108 166320
rect 190460 166268 190512 166320
rect 198740 166268 198792 166320
rect 263600 166268 263652 166320
rect 90364 165588 90416 165640
rect 208400 165588 208452 165640
rect 154488 164908 154540 164960
rect 195796 164908 195848 164960
rect 197544 164908 197596 164960
rect 60464 164840 60516 164892
rect 83464 164840 83516 164892
rect 193864 164840 193916 164892
rect 262588 164840 262640 164892
rect 210424 164160 210476 164212
rect 293960 164160 294012 164212
rect 294420 164160 294472 164212
rect 82912 163548 82964 163600
rect 154396 163548 154448 163600
rect 88984 163480 89036 163532
rect 169760 163480 169812 163532
rect 196808 163480 196860 163532
rect 294420 163480 294472 163532
rect 582932 163480 582984 163532
rect 208400 162800 208452 162852
rect 270684 162800 270736 162852
rect 222200 161848 222252 161900
rect 222936 161848 222988 161900
rect 152648 161508 152700 161560
rect 222200 161508 222252 161560
rect 73068 161440 73120 161492
rect 198740 161440 198792 161492
rect 234620 160692 234672 160744
rect 259552 160692 259604 160744
rect 156788 160148 156840 160200
rect 157248 160148 157300 160200
rect 224224 160148 224276 160200
rect 64604 160080 64656 160132
rect 165068 160080 165120 160132
rect 194600 160080 194652 160132
rect 195888 160080 195940 160132
rect 276664 160080 276716 160132
rect 242900 159468 242952 159520
rect 243544 159468 243596 159520
rect 119344 159332 119396 159384
rect 242900 159332 242952 159384
rect 249064 159332 249116 159384
rect 261208 159332 261260 159384
rect 91836 158720 91888 158772
rect 92388 158720 92440 158772
rect 220820 158720 220872 158772
rect 65984 157972 66036 158024
rect 182824 157972 182876 158024
rect 202788 157972 202840 158024
rect 267740 157972 267792 158024
rect 105544 157360 105596 157412
rect 225052 157360 225104 157412
rect 53564 156612 53616 156664
rect 67824 156612 67876 156664
rect 68652 156612 68704 156664
rect 196624 156612 196676 156664
rect 205732 156612 205784 156664
rect 97264 156408 97316 156460
rect 97908 156408 97960 156460
rect 247040 156408 247092 156460
rect 247684 156408 247736 156460
rect 68652 156000 68704 156052
rect 189908 156000 189960 156052
rect 207112 156000 207164 156052
rect 247040 156000 247092 156052
rect 97908 155932 97960 155984
rect 226432 155932 226484 155984
rect 56232 155864 56284 155916
rect 56508 155864 56560 155916
rect 215392 155184 215444 155236
rect 222292 155184 222344 155236
rect 263600 155184 263652 155236
rect 299480 155184 299532 155236
rect 204352 154912 204404 154964
rect 204904 154912 204956 154964
rect 56508 154640 56560 154692
rect 137468 154640 137520 154692
rect 91928 154572 91980 154624
rect 201684 154572 201736 154624
rect 202788 154572 202840 154624
rect 204904 154572 204956 154624
rect 263600 154572 263652 154624
rect 222200 154504 222252 154556
rect 282920 154504 282972 154556
rect 189172 153824 189224 153876
rect 201500 153824 201552 153876
rect 237380 153824 237432 153876
rect 265624 153824 265676 153876
rect 342260 153824 342312 153876
rect 67272 153280 67324 153332
rect 112444 153280 112496 153332
rect 129096 153280 129148 153332
rect 223580 153280 223632 153332
rect 49516 153212 49568 153264
rect 186228 153212 186280 153264
rect 211160 153144 211212 153196
rect 271880 153144 271932 153196
rect 192576 153076 192628 153128
rect 237380 153076 237432 153128
rect 92756 152532 92808 152584
rect 154488 152532 154540 152584
rect 133236 152464 133288 152516
rect 207112 152464 207164 152516
rect 54944 151784 54996 151836
rect 127716 151784 127768 151836
rect 80060 151104 80112 151156
rect 90364 151104 90416 151156
rect 57796 151036 57848 151088
rect 189172 151036 189224 151088
rect 170496 150492 170548 150544
rect 224960 150492 225012 150544
rect 189172 150424 189224 150476
rect 189816 150424 189868 150476
rect 218244 150424 218296 150476
rect 323584 150424 323636 150476
rect 197360 149948 197412 150000
rect 197636 149948 197688 150000
rect 191104 149812 191156 149864
rect 224868 149812 224920 149864
rect 81992 149744 82044 149796
rect 102140 149744 102192 149796
rect 218336 149744 218388 149796
rect 268108 149744 268160 149796
rect 70308 149676 70360 149728
rect 77944 149676 77996 149728
rect 86868 149676 86920 149728
rect 126336 149676 126388 149728
rect 216680 149676 216732 149728
rect 224868 149676 224920 149728
rect 305644 149676 305696 149728
rect 82820 149472 82872 149524
rect 86316 149472 86368 149524
rect 230020 148996 230072 149048
rect 276020 148996 276072 149048
rect 52460 148316 52512 148368
rect 80704 148316 80756 148368
rect 91008 148316 91060 148368
rect 127624 148316 127676 148368
rect 220912 148384 220964 148436
rect 186228 148316 186280 148368
rect 188804 148316 188856 148368
rect 196716 148316 196768 148368
rect 213920 148316 213972 148368
rect 317420 148316 317472 148368
rect 57888 147636 57940 147688
rect 184296 147636 184348 147688
rect 211896 147636 211948 147688
rect 213920 147636 213972 147688
rect 97816 147092 97868 147144
rect 101404 147092 101456 147144
rect 215392 146956 215444 147008
rect 216220 146956 216272 147008
rect 4252 146888 4304 146940
rect 97448 146888 97500 146940
rect 255320 146752 255372 146804
rect 256056 146752 256108 146804
rect 113916 146344 113968 146396
rect 227812 146344 227864 146396
rect 80520 146276 80572 146328
rect 208492 146276 208544 146328
rect 214564 146276 214616 146328
rect 255320 146276 255372 146328
rect 3424 146208 3476 146260
rect 86868 146208 86920 146260
rect 213184 146208 213236 146260
rect 216772 146208 216824 146260
rect 94320 145596 94372 145648
rect 129096 145596 129148 145648
rect 252836 145596 252888 145648
rect 327080 145596 327132 145648
rect 71780 145528 71832 145580
rect 107568 145528 107620 145580
rect 198004 145528 198056 145580
rect 198832 145528 198884 145580
rect 287244 145528 287296 145580
rect 86868 144916 86920 144968
rect 87696 144916 87748 144968
rect 177304 144916 177356 144968
rect 209872 144916 209924 144968
rect 222936 144848 222988 144900
rect 226524 144848 226576 144900
rect 200212 144440 200264 144492
rect 207756 144440 207808 144492
rect 78680 144372 78732 144424
rect 82176 144372 82228 144424
rect 102324 144168 102376 144220
rect 184204 144168 184256 144220
rect 188436 144168 188488 144220
rect 196532 144168 196584 144220
rect 206836 144168 206888 144220
rect 284944 144168 284996 144220
rect 298744 144168 298796 144220
rect 53656 143556 53708 143608
rect 153936 143556 153988 143608
rect 169668 143556 169720 143608
rect 202052 143624 202104 143676
rect 196808 143556 196860 143608
rect 201316 143556 201368 143608
rect 214012 143488 214064 143540
rect 216864 143488 216916 143540
rect 219532 143488 219584 143540
rect 220084 143488 220136 143540
rect 82912 142808 82964 142860
rect 83556 142808 83608 142860
rect 88432 142264 88484 142316
rect 213276 142264 213328 142316
rect 189080 142196 189132 142248
rect 206836 142196 206888 142248
rect 215300 142196 215352 142248
rect 221464 142196 221516 142248
rect 223212 142196 223264 142248
rect 211804 142128 211856 142180
rect 212816 142128 212868 142180
rect 219992 142128 220044 142180
rect 225604 142128 225656 142180
rect 240784 142128 240836 142180
rect 76288 141380 76340 141432
rect 159456 141380 159508 141432
rect 203156 141380 203208 141432
rect 218796 141380 218848 141432
rect 227904 141380 227956 141432
rect 223580 141176 223632 141228
rect 224500 141176 224552 141228
rect 65892 140836 65944 140888
rect 70492 140836 70544 140888
rect 58992 140768 59044 140820
rect 59268 140768 59320 140820
rect 105636 140768 105688 140820
rect 186320 140768 186372 140820
rect 193220 140768 193272 140820
rect 214380 140836 214432 140888
rect 280896 140836 280948 140888
rect 288624 140836 288676 140888
rect 203432 140768 203484 140820
rect 287704 140768 287756 140820
rect 80428 140700 80480 140752
rect 83464 140700 83516 140752
rect 193312 140700 193364 140752
rect 221464 140700 221516 140752
rect 251916 140700 251968 140752
rect 210056 140496 210108 140548
rect 193036 140428 193088 140480
rect 197360 140428 197412 140480
rect 63132 140088 63184 140140
rect 76012 140088 76064 140140
rect 46848 140020 46900 140072
rect 71412 140020 71464 140072
rect 75828 140020 75880 140072
rect 91928 140020 91980 140072
rect 86868 139408 86920 139460
rect 215392 140428 215444 140480
rect 224592 140428 224644 140480
rect 225696 140428 225748 140480
rect 289084 140020 289136 140072
rect 251180 139408 251232 139460
rect 251916 139408 251968 139460
rect 134616 139340 134668 139392
rect 188528 139340 188580 139392
rect 226340 139340 226392 139392
rect 236092 139340 236144 139392
rect 78036 138728 78088 138780
rect 113824 138728 113876 138780
rect 52092 138660 52144 138712
rect 72332 138660 72384 138712
rect 81900 138660 81952 138712
rect 177304 138660 177356 138712
rect 75920 138048 75972 138100
rect 76380 138048 76432 138100
rect 2872 137912 2924 137964
rect 73068 137912 73120 137964
rect 86132 137912 86184 137964
rect 193312 137912 193364 137964
rect 226708 137912 226760 137964
rect 240140 137912 240192 137964
rect 241428 137912 241480 137964
rect 67180 137300 67232 137352
rect 67548 137300 67600 137352
rect 64788 137232 64840 137284
rect 69204 137232 69256 137284
rect 79600 137232 79652 137284
rect 189080 137232 189132 137284
rect 241428 137232 241480 137284
rect 282184 137232 282236 137284
rect 75552 136688 75604 136740
rect 78772 136688 78824 136740
rect 78496 136620 78548 136672
rect 79324 136620 79376 136672
rect 85488 136620 85540 136672
rect 86224 136620 86276 136672
rect 173808 136552 173860 136604
rect 191748 136552 191800 136604
rect 226708 136280 226760 136332
rect 229836 136280 229888 136332
rect 91744 136144 91796 136196
rect 95976 136144 96028 136196
rect 91008 135872 91060 135924
rect 126612 135872 126664 135924
rect 240048 135872 240100 135924
rect 333980 135872 334032 135924
rect 91192 135532 91244 135584
rect 91836 135532 91888 135584
rect 4804 135260 4856 135312
rect 91192 135260 91244 135312
rect 184204 135260 184256 135312
rect 191748 135260 191800 135312
rect 97448 135192 97500 135244
rect 182916 135192 182968 135244
rect 188988 135192 189040 135244
rect 189724 135192 189776 135244
rect 226340 135192 226392 135244
rect 258724 135192 258776 135244
rect 70308 134988 70360 135040
rect 72424 134988 72476 135040
rect 3424 134512 3476 134564
rect 75920 134580 75972 134632
rect 94412 134580 94464 134632
rect 95148 134580 95200 134632
rect 95148 133968 95200 134020
rect 156788 133968 156840 134020
rect 188896 133968 188948 134020
rect 190460 133968 190512 134020
rect 226708 133900 226760 133952
rect 302884 133900 302936 133952
rect 64604 133832 64656 133884
rect 66812 133832 66864 133884
rect 96712 133832 96764 133884
rect 114008 133832 114060 133884
rect 165068 133832 165120 133884
rect 186320 133832 186372 133884
rect 226340 133832 226392 133884
rect 269120 133832 269172 133884
rect 226708 133764 226760 133816
rect 233884 133764 233936 133816
rect 226432 133492 226484 133544
rect 226708 133492 226760 133544
rect 113824 133152 113876 133204
rect 126428 133152 126480 133204
rect 134616 133152 134668 133204
rect 148508 133152 148560 133204
rect 148692 133152 148744 133204
rect 184388 133152 184440 133204
rect 50988 132404 51040 132456
rect 66812 132404 66864 132456
rect 105636 132404 105688 132456
rect 57704 132336 57756 132388
rect 66260 132336 66312 132388
rect 96712 132336 96764 132388
rect 148600 132336 148652 132388
rect 188344 132404 188396 132456
rect 191656 132404 191708 132456
rect 226340 132404 226392 132456
rect 231952 132404 232004 132456
rect 191104 132336 191156 132388
rect 41328 131724 41380 131776
rect 48320 131724 48372 131776
rect 231216 131724 231268 131776
rect 276020 131724 276072 131776
rect 148416 131112 148468 131164
rect 153844 131112 153896 131164
rect 176016 131044 176068 131096
rect 190000 131044 190052 131096
rect 226708 131044 226760 131096
rect 230480 131044 230532 131096
rect 273260 131044 273312 131096
rect 226800 130976 226852 131028
rect 240324 130976 240376 131028
rect 96804 130364 96856 130416
rect 170496 130364 170548 130416
rect 176016 130364 176068 130416
rect 176568 130364 176620 130416
rect 96712 130160 96764 130212
rect 102968 130160 103020 130212
rect 94780 129684 94832 129736
rect 95884 129684 95936 129736
rect 94964 129616 95016 129668
rect 187516 129684 187568 129736
rect 191748 129684 191800 129736
rect 229744 129684 229796 129736
rect 259460 129684 259512 129736
rect 226524 129004 226576 129056
rect 226708 129004 226760 129056
rect 299480 129004 299532 129056
rect 63224 128256 63276 128308
rect 66812 128256 66864 128308
rect 97632 128256 97684 128308
rect 142988 128256 143040 128308
rect 226708 127644 226760 127696
rect 226892 127644 226944 127696
rect 260104 127644 260156 127696
rect 126336 127576 126388 127628
rect 135996 127576 136048 127628
rect 227996 127576 228048 127628
rect 267924 127576 267976 127628
rect 268384 127576 268436 127628
rect 295340 127576 295392 127628
rect 97264 126896 97316 126948
rect 111248 126896 111300 126948
rect 158076 126896 158128 126948
rect 192300 126964 192352 127016
rect 192852 126964 192904 127016
rect 226340 126896 226392 126948
rect 242900 126896 242952 126948
rect 243360 126896 243412 126948
rect 295340 126896 295392 126948
rect 302332 126896 302384 126948
rect 182824 126828 182876 126880
rect 192392 126828 192444 126880
rect 108488 126216 108540 126268
rect 187516 126216 187568 126268
rect 243360 126216 243412 126268
rect 351920 126216 351972 126268
rect 187516 125672 187568 125724
rect 190368 125672 190420 125724
rect 52184 125536 52236 125588
rect 66904 125536 66956 125588
rect 97540 125536 97592 125588
rect 148692 125536 148744 125588
rect 167736 125536 167788 125588
rect 190276 125536 190328 125588
rect 56508 124856 56560 124908
rect 66812 124856 66864 124908
rect 96620 124856 96672 124908
rect 175924 124856 175976 124908
rect 232504 124856 232556 124908
rect 295432 124856 295484 124908
rect 188804 124788 188856 124840
rect 192944 124788 192996 124840
rect 226524 124720 226576 124772
rect 229744 124720 229796 124772
rect 61936 124108 61988 124160
rect 66260 124108 66312 124160
rect 97908 124108 97960 124160
rect 152648 124108 152700 124160
rect 226340 124108 226392 124160
rect 229100 124108 229152 124160
rect 280804 124108 280856 124160
rect 582840 124108 582892 124160
rect 228364 123428 228416 123480
rect 255964 123428 256016 123480
rect 59084 122748 59136 122800
rect 66352 122748 66404 122800
rect 97540 122748 97592 122800
rect 119344 122748 119396 122800
rect 155868 122748 155920 122800
rect 191748 122816 191800 122868
rect 226340 122748 226392 122800
rect 247040 122748 247092 122800
rect 189816 122340 189868 122392
rect 190368 122340 190420 122392
rect 112444 122068 112496 122120
rect 188344 122068 188396 122120
rect 225696 122068 225748 122120
rect 313280 122068 313332 122120
rect 61844 121388 61896 121440
rect 66812 121388 66864 121440
rect 97724 121388 97776 121440
rect 151176 121388 151228 121440
rect 159548 121388 159600 121440
rect 191196 121388 191248 121440
rect 226432 121388 226484 121440
rect 244372 121388 244424 121440
rect 240876 120708 240928 120760
rect 274640 120708 274692 120760
rect 184756 120640 184808 120692
rect 191748 120640 191800 120692
rect 97540 120096 97592 120148
rect 105544 120096 105596 120148
rect 49516 120028 49568 120080
rect 66812 120028 66864 120080
rect 97724 120028 97776 120080
rect 122104 120028 122156 120080
rect 184296 120028 184348 120080
rect 191748 120028 191800 120080
rect 284944 119348 284996 119400
rect 289912 119348 289964 119400
rect 57796 118600 57848 118652
rect 66904 118600 66956 118652
rect 97908 118600 97960 118652
rect 133236 118600 133288 118652
rect 64512 118532 64564 118584
rect 66812 118532 66864 118584
rect 97816 117920 97868 117972
rect 100024 117920 100076 117972
rect 173256 117920 173308 117972
rect 180156 117920 180208 117972
rect 187700 117920 187752 117972
rect 187700 117376 187752 117428
rect 188988 117376 189040 117428
rect 191748 117376 191800 117428
rect 226524 117376 226576 117428
rect 233884 117376 233936 117428
rect 226708 117308 226760 117360
rect 244280 117308 244332 117360
rect 97356 117240 97408 117292
rect 145656 117240 145708 117292
rect 185676 117240 185728 117292
rect 191748 117240 191800 117292
rect 54944 117172 54996 117224
rect 66812 117172 66864 117224
rect 97908 117172 97960 117224
rect 136088 117172 136140 117224
rect 231768 116560 231820 116612
rect 262404 116560 262456 116612
rect 291660 116560 291712 116612
rect 304264 116560 304316 116612
rect 185768 116016 185820 116068
rect 191288 116016 191340 116068
rect 226708 115948 226760 116000
rect 230480 115948 230532 116000
rect 231768 115948 231820 116000
rect 57888 115880 57940 115932
rect 66812 115880 66864 115932
rect 175188 115880 175240 115932
rect 191012 115880 191064 115932
rect 63316 115268 63368 115320
rect 66812 115268 66864 115320
rect 233332 115200 233384 115252
rect 280160 115200 280212 115252
rect 97540 114588 97592 114640
rect 112444 114588 112496 114640
rect 97908 114520 97960 114572
rect 170496 114520 170548 114572
rect 226340 114520 226392 114572
rect 233332 114520 233384 114572
rect 58992 114452 59044 114504
rect 66812 114452 66864 114504
rect 7564 113772 7616 113824
rect 65984 113772 66036 113824
rect 96712 113772 96764 113824
rect 134800 113772 134852 113824
rect 160928 113772 160980 113824
rect 183376 113772 183428 113824
rect 188252 113228 188304 113280
rect 191196 113228 191248 113280
rect 183376 113160 183428 113212
rect 191748 113160 191800 113212
rect 63132 113092 63184 113144
rect 66812 113092 66864 113144
rect 226708 113092 226760 113144
rect 233240 113092 233292 113144
rect 60556 113024 60608 113076
rect 66904 113024 66956 113076
rect 225604 112480 225656 112532
rect 253020 112480 253072 112532
rect 104256 112412 104308 112464
rect 191564 112412 191616 112464
rect 233240 112412 233292 112464
rect 324412 112412 324464 112464
rect 98092 111936 98144 111988
rect 101588 111936 101640 111988
rect 96896 111868 96948 111920
rect 98644 111868 98696 111920
rect 97908 111800 97960 111852
rect 160744 111800 160796 111852
rect 55128 111732 55180 111784
rect 66812 111732 66864 111784
rect 97356 111732 97408 111784
rect 113916 111732 113968 111784
rect 153936 111732 153988 111784
rect 191380 111732 191432 111784
rect 252652 111732 252704 111784
rect 253020 111732 253072 111784
rect 260196 111732 260248 111784
rect 226340 111120 226392 111172
rect 229100 111120 229152 111172
rect 236000 111120 236052 111172
rect 159364 111052 159416 111104
rect 185768 111052 185820 111104
rect 226524 111052 226576 111104
rect 291200 111052 291252 111104
rect 2872 110780 2924 110832
rect 4804 110780 4856 110832
rect 291200 110440 291252 110492
rect 291844 110440 291896 110492
rect 59268 110372 59320 110424
rect 66812 110372 66864 110424
rect 226984 109760 227036 109812
rect 267832 109760 267884 109812
rect 104256 109692 104308 109744
rect 149796 109692 149848 109744
rect 153844 109692 153896 109744
rect 188252 109692 188304 109744
rect 225604 109692 225656 109744
rect 252560 109692 252612 109744
rect 345664 109692 345716 109744
rect 48228 109012 48280 109064
rect 52552 109012 52604 109064
rect 66904 109012 66956 109064
rect 53656 108944 53708 108996
rect 66720 108944 66772 108996
rect 97908 108944 97960 108996
rect 114652 108944 114704 108996
rect 115848 108944 115900 108996
rect 166448 108944 166500 108996
rect 190276 108944 190328 108996
rect 226524 108944 226576 108996
rect 245660 108944 245712 108996
rect 64788 108876 64840 108928
rect 66444 108876 66496 108928
rect 183468 108876 183520 108928
rect 191196 108876 191248 108928
rect 104900 108332 104952 108384
rect 144184 108332 144236 108384
rect 115848 108264 115900 108316
rect 180156 108264 180208 108316
rect 227076 108264 227128 108316
rect 227720 108264 227772 108316
rect 270592 108264 270644 108316
rect 189080 107720 189132 107772
rect 191196 107720 191248 107772
rect 163504 107584 163556 107636
rect 191748 107584 191800 107636
rect 226708 107584 226760 107636
rect 284392 107584 284444 107636
rect 285036 107584 285088 107636
rect 187608 107516 187660 107568
rect 189080 107516 189132 107568
rect 7564 106904 7616 106956
rect 66996 106904 67048 106956
rect 97816 106904 97868 106956
rect 169116 106904 169168 106956
rect 284392 106904 284444 106956
rect 349160 106904 349212 106956
rect 96988 106632 97040 106684
rect 100024 106632 100076 106684
rect 97540 106020 97592 106072
rect 101496 106020 101548 106072
rect 96896 105884 96948 105936
rect 98736 105884 98788 105936
rect 188344 105884 188396 105936
rect 191748 105884 191800 105936
rect 48136 105544 48188 105596
rect 64788 105544 64840 105596
rect 66536 105544 66588 105596
rect 56416 104796 56468 104848
rect 66352 104796 66404 104848
rect 97724 104796 97776 104848
rect 111064 104864 111116 104916
rect 177304 104864 177356 104916
rect 186228 104864 186280 104916
rect 191748 104864 191800 104916
rect 226708 104864 226760 104916
rect 278044 104796 278096 104848
rect 285680 104796 285732 104848
rect 96528 103504 96580 103556
rect 178776 103504 178828 103556
rect 226524 103504 226576 103556
rect 231952 103504 232004 103556
rect 280804 103504 280856 103556
rect 64696 103436 64748 103488
rect 66628 103436 66680 103488
rect 97908 103028 97960 103080
rect 99564 103028 99616 103080
rect 99564 102756 99616 102808
rect 188344 102756 188396 102808
rect 226708 102756 226760 102808
rect 227812 102756 227864 102808
rect 281540 102756 281592 102808
rect 309784 102756 309836 102808
rect 63408 102212 63460 102264
rect 66076 102212 66128 102264
rect 66536 102212 66588 102264
rect 67364 102144 67416 102196
rect 67640 102144 67692 102196
rect 100668 102144 100720 102196
rect 184296 102144 184348 102196
rect 186964 102144 187016 102196
rect 191656 102144 191708 102196
rect 226708 102144 226760 102196
rect 237564 102144 237616 102196
rect 226340 102076 226392 102128
rect 266360 102076 266412 102128
rect 97908 102008 97960 102060
rect 130568 102008 130620 102060
rect 130568 101464 130620 101516
rect 148508 101464 148560 101516
rect 113916 101396 113968 101448
rect 158628 101396 158680 101448
rect 181996 101396 182048 101448
rect 61936 100852 61988 100904
rect 66812 100852 66864 100904
rect 181996 100716 182048 100768
rect 191656 100716 191708 100768
rect 97908 100648 97960 100700
rect 100668 100648 100720 100700
rect 185584 100648 185636 100700
rect 190644 100648 190696 100700
rect 60648 99628 60700 99680
rect 63408 99628 63460 99680
rect 66812 99628 66864 99680
rect 97540 99356 97592 99408
rect 131028 99356 131080 99408
rect 226432 99356 226484 99408
rect 229192 99356 229244 99408
rect 322204 99356 322256 99408
rect 62028 99288 62080 99340
rect 66812 99288 66864 99340
rect 237380 98676 237432 98728
rect 250536 98676 250588 98728
rect 226524 98608 226576 98660
rect 264980 98608 265032 98660
rect 96896 98336 96948 98388
rect 98920 98336 98972 98388
rect 100116 98064 100168 98116
rect 164148 98064 164200 98116
rect 164884 98064 164936 98116
rect 184388 98064 184440 98116
rect 191656 98064 191708 98116
rect 97356 97996 97408 98048
rect 189816 97996 189868 98048
rect 181536 97928 181588 97980
rect 190644 97928 190696 97980
rect 96896 96840 96948 96892
rect 98828 96840 98880 96892
rect 3056 96636 3108 96688
rect 62764 96636 62816 96688
rect 97908 96636 97960 96688
rect 188436 96636 188488 96688
rect 226524 95956 226576 96008
rect 228364 95956 228416 96008
rect 95424 95208 95476 95260
rect 193128 95208 193180 95260
rect 52368 95140 52420 95192
rect 66812 95140 66864 95192
rect 95976 95140 96028 95192
rect 182088 95140 182140 95192
rect 96988 94460 97040 94512
rect 102232 94460 102284 94512
rect 182088 94460 182140 94512
rect 193404 94460 193456 94512
rect 227628 94460 227680 94512
rect 263692 94460 263744 94512
rect 226616 94392 226668 94444
rect 228364 94392 228416 94444
rect 53748 93780 53800 93832
rect 68008 93780 68060 93832
rect 97908 93780 97960 93832
rect 108396 93780 108448 93832
rect 171048 93100 171100 93152
rect 183560 93100 183612 93152
rect 191748 93100 191800 93152
rect 231308 93100 231360 93152
rect 249156 93100 249208 93152
rect 250536 93100 250588 93152
rect 331220 93100 331272 93152
rect 69020 92896 69072 92948
rect 67364 92828 67416 92880
rect 68468 92828 68520 92880
rect 70262 92692 70314 92744
rect 91790 92692 91842 92744
rect 95240 92692 95292 92744
rect 88662 92624 88714 92676
rect 89628 92624 89680 92676
rect 90134 92624 90186 92676
rect 74632 92556 74684 92608
rect 75782 92556 75834 92608
rect 80152 92556 80204 92608
rect 80934 92556 80986 92608
rect 50896 92352 50948 92404
rect 72792 92352 72844 92404
rect 126520 92488 126572 92540
rect 218796 92488 218848 92540
rect 221924 92488 221976 92540
rect 232504 92488 232556 92540
rect 184296 92420 184348 92472
rect 229192 92420 229244 92472
rect 213184 92352 213236 92404
rect 242256 92352 242308 92404
rect 67456 92284 67508 92336
rect 184388 92284 184440 92336
rect 193128 91740 193180 91792
rect 202144 91740 202196 91792
rect 65892 90992 65944 91044
rect 71136 90992 71188 91044
rect 84660 90992 84712 91044
rect 116124 90992 116176 91044
rect 212448 90992 212500 91044
rect 221372 90992 221424 91044
rect 258080 90992 258132 91044
rect 85212 90312 85264 90364
rect 94504 90312 94556 90364
rect 213460 90312 213512 90364
rect 235264 90312 235316 90364
rect 68928 90244 68980 90296
rect 71044 90244 71096 90296
rect 223764 90244 223816 90296
rect 224868 90244 224920 90296
rect 105544 89700 105596 89752
rect 106372 89700 106424 89752
rect 127624 89700 127676 89752
rect 128360 89700 128412 89752
rect 245660 89700 245712 89752
rect 246304 89700 246356 89752
rect 580264 89700 580316 89752
rect 49608 89632 49660 89684
rect 79416 89632 79468 89684
rect 85580 89632 85632 89684
rect 117320 89632 117372 89684
rect 117780 89632 117832 89684
rect 124128 89632 124180 89684
rect 217692 89632 217744 89684
rect 220636 89632 220688 89684
rect 273352 89632 273404 89684
rect 84108 89564 84160 89616
rect 98736 89564 98788 89616
rect 193404 89564 193456 89616
rect 199384 89564 199436 89616
rect 203708 89564 203760 89616
rect 284300 89564 284352 89616
rect 123576 89224 123628 89276
rect 124128 89224 124180 89276
rect 284300 88952 284352 89004
rect 582840 88952 582892 89004
rect 67272 88272 67324 88324
rect 113916 88272 113968 88324
rect 117780 88272 117832 88324
rect 213460 88272 213512 88324
rect 214564 88272 214616 88324
rect 262220 88272 262272 88324
rect 60464 88204 60516 88256
rect 82636 88204 82688 88256
rect 83464 88204 83516 88256
rect 86684 88204 86736 88256
rect 100760 88204 100812 88256
rect 188528 88204 188580 88256
rect 196072 88204 196124 88256
rect 206376 88204 206428 88256
rect 207388 88204 207440 88256
rect 215852 88204 215904 88256
rect 216036 88204 216088 88256
rect 242164 88204 242216 88256
rect 89812 86912 89864 86964
rect 124312 86912 124364 86964
rect 218244 86912 218296 86964
rect 219532 86912 219584 86964
rect 220084 86912 220136 86964
rect 245660 86912 245712 86964
rect 73804 86844 73856 86896
rect 185124 86844 185176 86896
rect 227720 86844 227772 86896
rect 95976 86776 96028 86828
rect 228364 86232 228416 86284
rect 241520 86232 241572 86284
rect 197360 85552 197412 85604
rect 198004 85552 198056 85604
rect 52368 85484 52420 85536
rect 52552 85484 52604 85536
rect 87236 85484 87288 85536
rect 117964 85484 118016 85536
rect 215392 85484 215444 85536
rect 65984 85416 66036 85468
rect 159364 85416 159416 85468
rect 238484 84872 238536 84924
rect 307024 84872 307076 84924
rect 191748 84804 191800 84856
rect 270592 84804 270644 84856
rect 3332 84192 3384 84244
rect 52368 84192 52420 84244
rect 69020 84124 69072 84176
rect 169024 84124 169076 84176
rect 193312 84124 193364 84176
rect 216680 84124 216732 84176
rect 261484 84124 261536 84176
rect 116032 84056 116084 84108
rect 213920 84056 213972 84108
rect 222292 83036 222344 83088
rect 222844 83036 222896 83088
rect 193312 82832 193364 82884
rect 193956 82832 194008 82884
rect 216680 82832 216732 82884
rect 217324 82832 217376 82884
rect 222844 82832 222896 82884
rect 339500 82832 339552 82884
rect 88340 82764 88392 82816
rect 123576 82764 123628 82816
rect 188344 82764 188396 82816
rect 227812 82764 227864 82816
rect 80244 82696 80296 82748
rect 105544 82696 105596 82748
rect 178040 82696 178092 82748
rect 179328 82696 179380 82748
rect 200120 82696 200172 82748
rect 201408 82696 201460 82748
rect 201408 82084 201460 82136
rect 245660 82084 245712 82136
rect 52368 81336 52420 81388
rect 153844 81336 153896 81388
rect 178776 81336 178828 81388
rect 231952 81336 232004 81388
rect 71872 81268 71924 81320
rect 172520 81268 172572 81320
rect 173808 81268 173860 81320
rect 164148 81200 164200 81252
rect 195980 81200 196032 81252
rect 210516 80656 210568 80708
rect 582932 80656 582984 80708
rect 195980 80044 196032 80096
rect 196624 80044 196676 80096
rect 80060 79976 80112 80028
rect 161480 79976 161532 80028
rect 177304 79976 177356 80028
rect 224960 79976 225012 80028
rect 62764 79908 62816 79960
rect 96620 79908 96672 79960
rect 205640 79908 205692 79960
rect 205640 79500 205692 79552
rect 206284 79500 206336 79552
rect 98644 79296 98696 79348
rect 113824 79296 113876 79348
rect 75828 78616 75880 78668
rect 178040 78616 178092 78668
rect 180156 78616 180208 78668
rect 225052 78616 225104 78668
rect 173808 78548 173860 78600
rect 197452 78548 197504 78600
rect 198004 78548 198056 78600
rect 198740 77936 198792 77988
rect 240140 77936 240192 77988
rect 288348 77936 288400 77988
rect 345020 77936 345072 77988
rect 92480 77188 92532 77240
rect 127624 77188 127676 77240
rect 148508 77188 148560 77240
rect 237564 77188 237616 77240
rect 238024 77188 238076 77240
rect 173256 77120 173308 77172
rect 244280 77120 244332 77172
rect 70308 76508 70360 76560
rect 166356 76508 166408 76560
rect 280068 76508 280120 76560
rect 292672 76508 292724 76560
rect 244280 76304 244332 76356
rect 245016 76304 245068 76356
rect 169116 75828 169168 75880
rect 229100 75828 229152 75880
rect 193220 75760 193272 75812
rect 193864 75760 193916 75812
rect 244924 75760 244976 75812
rect 74540 75148 74592 75200
rect 167644 75148 167696 75200
rect 255228 74536 255280 74588
rect 318064 74536 318116 74588
rect 61936 74468 61988 74520
rect 186964 74468 187016 74520
rect 201500 74468 201552 74520
rect 166356 74400 166408 74452
rect 194600 74400 194652 74452
rect 85580 73788 85632 73840
rect 160836 73788 160888 73840
rect 61384 73176 61436 73228
rect 61936 73176 61988 73228
rect 194600 73176 194652 73228
rect 195244 73176 195296 73228
rect 80152 73108 80204 73160
rect 103520 73108 103572 73160
rect 207020 73108 207072 73160
rect 197360 73040 197412 73092
rect 249800 73108 249852 73160
rect 583024 73108 583076 73160
rect 88340 72428 88392 72480
rect 184940 72428 184992 72480
rect 207020 72428 207072 72480
rect 269028 72428 269080 72480
rect 269764 72428 269816 72480
rect 3516 71680 3568 71732
rect 95332 71680 95384 71732
rect 131028 71680 131080 71732
rect 226432 71680 226484 71732
rect 92480 71000 92532 71052
rect 164976 71000 165028 71052
rect 192852 71000 192904 71052
rect 281540 71000 281592 71052
rect 226432 70388 226484 70440
rect 226984 70388 227036 70440
rect 66076 70320 66128 70372
rect 185584 70320 185636 70372
rect 160744 70252 160796 70304
rect 233332 70252 233384 70304
rect 94688 68960 94740 69012
rect 222844 68960 222896 69012
rect 170496 68892 170548 68944
rect 233884 68892 233936 68944
rect 93860 68280 93912 68332
rect 106924 68280 106976 68332
rect 109040 68280 109092 68332
rect 126336 68280 126388 68332
rect 235264 68280 235316 68332
rect 287060 68280 287112 68332
rect 74632 67532 74684 67584
rect 201500 67532 201552 67584
rect 112444 67464 112496 67516
rect 230480 67464 230532 67516
rect 87052 66172 87104 66224
rect 215300 66104 215352 66156
rect 215944 66104 215996 66156
rect 188896 65492 188948 65544
rect 220084 65492 220136 65544
rect 97264 64812 97316 64864
rect 241520 64812 241572 64864
rect 108396 64132 108448 64184
rect 124864 64132 124916 64184
rect 202972 63520 203024 63572
rect 322296 63520 322348 63572
rect 71044 63452 71096 63504
rect 193864 63452 193916 63504
rect 86960 63384 87012 63436
rect 121552 63384 121604 63436
rect 190368 62772 190420 62824
rect 249800 62772 249852 62824
rect 215208 62500 215260 62552
rect 216036 62500 216088 62552
rect 127624 62024 127676 62076
rect 222200 62024 222252 62076
rect 240784 61344 240836 61396
rect 269764 61344 269816 61396
rect 222200 60732 222252 60784
rect 222844 60732 222896 60784
rect 89628 60664 89680 60716
rect 217324 60664 217376 60716
rect 181996 59984 182048 60036
rect 233884 59984 233936 60036
rect 94504 59304 94556 59356
rect 213184 59304 213236 59356
rect 193956 58624 194008 58676
rect 264980 58624 265032 58676
rect 77208 57876 77260 57928
rect 202972 57876 203024 57928
rect 199384 57196 199436 57248
rect 244280 57196 244332 57248
rect 83464 56516 83516 56568
rect 210424 56516 210476 56568
rect 105544 56448 105596 56500
rect 206376 56448 206428 56500
rect 46940 54476 46992 54528
rect 135904 54476 135956 54528
rect 184296 54476 184348 54528
rect 320272 54476 320324 54528
rect 87604 53048 87656 53100
rect 140044 53048 140096 53100
rect 192944 53048 192996 53100
rect 270500 53048 270552 53100
rect 75184 51756 75236 51808
rect 108304 51756 108356 51808
rect 97264 51688 97316 51740
rect 143540 51688 143592 51740
rect 239404 51688 239456 51740
rect 259460 51688 259512 51740
rect 2872 50328 2924 50380
rect 146944 50328 146996 50380
rect 202144 50328 202196 50380
rect 286324 50328 286376 50380
rect 71780 48968 71832 49020
rect 138664 48968 138716 49020
rect 189724 48968 189776 49020
rect 580172 48968 580224 49020
rect 53840 47540 53892 47592
rect 149704 47540 149756 47592
rect 187516 47540 187568 47592
rect 298100 47540 298152 47592
rect 3516 46180 3568 46232
rect 61384 46180 61436 46232
rect 217324 46180 217376 46232
rect 291936 46180 291988 46232
rect 291844 45568 291896 45620
rect 296812 45568 296864 45620
rect 64880 44820 64932 44872
rect 142896 44820 142948 44872
rect 193036 44820 193088 44872
rect 309140 44820 309192 44872
rect 99380 43392 99432 43444
rect 141424 43392 141476 43444
rect 210424 43392 210476 43444
rect 322940 43392 322992 43444
rect 66260 42032 66312 42084
rect 123484 42032 123536 42084
rect 213184 40672 213236 40724
rect 334072 40672 334124 40724
rect 75920 39312 75972 39364
rect 155316 39312 155368 39364
rect 98000 37884 98052 37936
rect 148416 37884 148468 37936
rect 204904 37204 204956 37256
rect 296720 37204 296772 37256
rect 298008 37204 298060 37256
rect 45560 36524 45612 36576
rect 166264 36524 166316 36576
rect 298008 36524 298060 36576
rect 343640 36524 343692 36576
rect 42800 35164 42852 35216
rect 170404 35164 170456 35216
rect 195244 35164 195296 35216
rect 311900 35164 311952 35216
rect 23480 33736 23532 33788
rect 173164 33736 173216 33788
rect 3516 33056 3568 33108
rect 57244 33056 57296 33108
rect 117320 32444 117372 32496
rect 156604 32444 156656 32496
rect 55220 32376 55272 32428
rect 134616 32376 134668 32428
rect 208400 32376 208452 32428
rect 278780 32376 278832 32428
rect 113180 31016 113232 31068
rect 157984 31016 158036 31068
rect 215944 31016 215996 31068
rect 266360 31016 266412 31068
rect 81440 29588 81492 29640
rect 179420 29588 179472 29640
rect 183376 29588 183428 29640
rect 263692 29588 263744 29640
rect 67640 28228 67692 28280
rect 171140 28228 171192 28280
rect 226984 28228 227036 28280
rect 277400 28228 277452 28280
rect 82820 26868 82872 26920
rect 151084 26868 151136 26920
rect 193864 25508 193916 25560
rect 291200 25508 291252 25560
rect 96620 24148 96672 24200
rect 130476 24148 130528 24200
rect 59360 24080 59412 24132
rect 131764 24080 131816 24132
rect 78680 22720 78732 22772
rect 145564 22720 145616 22772
rect 57980 21360 58032 21412
rect 137376 21360 137428 21412
rect 3424 20612 3476 20664
rect 90364 20612 90416 20664
rect 95240 19932 95292 19984
rect 162860 19932 162912 19984
rect 205548 19932 205600 19984
rect 288440 19932 288492 19984
rect 63500 18572 63552 18624
rect 178684 18572 178736 18624
rect 215208 18572 215260 18624
rect 284392 18572 284444 18624
rect 322204 18572 322256 18624
rect 332600 18572 332652 18624
rect 309784 17960 309836 18012
rect 316132 17960 316184 18012
rect 233884 17280 233936 17332
rect 251272 17280 251324 17332
rect 49700 17212 49752 17264
rect 162124 17212 162176 17264
rect 206284 17212 206336 17264
rect 233976 17212 234028 17264
rect 260104 17212 260156 17264
rect 336740 17212 336792 17264
rect 91560 15852 91612 15904
rect 129096 15852 129148 15904
rect 245016 15852 245068 15904
rect 256700 15852 256752 15904
rect 302884 15852 302936 15904
rect 314660 15852 314712 15904
rect 112 14492 164 14544
rect 96712 14492 96764 14544
rect 222844 14492 222896 14544
rect 302884 14492 302936 14544
rect 87512 14424 87564 14476
rect 231124 14424 231176 14476
rect 89904 13064 89956 13116
rect 155224 13064 155276 13116
rect 200764 13064 200816 13116
rect 340972 13064 341024 13116
rect 61568 11704 61620 11756
rect 133144 11704 133196 11756
rect 188988 11704 189040 11756
rect 280712 11704 280764 11756
rect 324412 11704 324464 11756
rect 325608 11704 325660 11756
rect 108120 10412 108172 10464
rect 142804 10412 142856 10464
rect 73344 10344 73396 10396
rect 108396 10344 108448 10396
rect 86408 10276 86460 10328
rect 126244 10276 126296 10328
rect 198004 10276 198056 10328
rect 342904 10276 342956 10328
rect 1676 8984 1728 9036
rect 87604 8984 87656 9036
rect 78588 8916 78640 8968
rect 168380 8916 168432 8968
rect 196624 8916 196676 8968
rect 258264 8916 258316 8968
rect 258724 8236 258776 8288
rect 261760 8236 261812 8288
rect 111616 7624 111668 7676
rect 148324 7624 148376 7676
rect 67732 7556 67784 7608
rect 125876 7556 125928 7608
rect 224868 7556 224920 7608
rect 254676 7556 254728 7608
rect 280804 7556 280856 7608
rect 330392 7556 330444 7608
rect 3424 6808 3476 6860
rect 7564 6808 7616 6860
rect 80888 6128 80940 6180
rect 130384 6128 130436 6180
rect 206376 6128 206428 6180
rect 247592 6128 247644 6180
rect 286324 6128 286376 6180
rect 329196 6128 329248 6180
rect 134524 5516 134576 5568
rect 136456 5516 136508 5568
rect 305644 5516 305696 5568
rect 309048 5516 309100 5568
rect 346952 5516 347004 5568
rect 349160 5516 349212 5568
rect 69112 4768 69164 4820
rect 152556 4768 152608 4820
rect 220084 4768 220136 4820
rect 244096 4768 244148 4820
rect 238024 4360 238076 4412
rect 239312 4360 239364 4412
rect 276020 4360 276072 4412
rect 278044 4360 278096 4412
rect 228364 4088 228416 4140
rect 248788 4088 248840 4140
rect 249064 4088 249116 4140
rect 267004 4088 267056 4140
rect 267740 4088 267792 4140
rect 302976 3952 303028 4004
rect 306748 3952 306800 4004
rect 323584 3952 323636 4004
rect 326804 3952 326856 4004
rect 150624 3612 150676 3664
rect 152464 3612 152516 3664
rect 251180 3544 251232 3596
rect 252376 3544 252428 3596
rect 316132 3544 316184 3596
rect 317328 3544 317380 3596
rect 2780 3476 2832 3528
rect 4068 3476 4120 3528
rect 19432 3476 19484 3528
rect 22744 3476 22796 3528
rect 35900 3476 35952 3528
rect 37188 3476 37240 3528
rect 84476 3476 84528 3528
rect 98644 3476 98696 3528
rect 101404 3476 101456 3528
rect 102232 3476 102284 3528
rect 118700 3476 118752 3528
rect 119896 3476 119948 3528
rect 143540 3476 143592 3528
rect 144736 3476 144788 3528
rect 270040 3476 270092 3528
rect 270592 3476 270644 3528
rect 289084 3476 289136 3528
rect 290188 3476 290240 3528
rect 291936 3476 291988 3528
rect 294880 3476 294932 3528
rect 298744 3476 298796 3528
rect 305552 3476 305604 3528
rect 307024 3476 307076 3528
rect 311440 3476 311492 3528
rect 319720 3476 319772 3528
rect 320180 3476 320232 3528
rect 351644 3476 351696 3528
rect 353300 3476 353352 3528
rect 63224 3408 63276 3460
rect 75184 3408 75236 3460
rect 77392 3408 77444 3460
rect 104256 3408 104308 3460
rect 140044 3408 140096 3460
rect 184204 3408 184256 3460
rect 233976 3408 234028 3460
rect 242900 3408 242952 3460
rect 276756 3408 276808 3460
rect 286600 3408 286652 3460
rect 581000 3272 581052 3324
rect 582564 3272 582616 3324
rect 318156 3204 318208 3256
rect 322112 3204 322164 3256
rect 348056 3204 348108 3256
rect 351920 3204 351972 3256
rect 260656 3136 260708 3188
rect 263600 3136 263652 3188
rect 269764 3136 269816 3188
rect 272432 3136 272484 3188
rect 322296 3136 322348 3188
rect 324412 3136 324464 3188
rect 345664 3136 345716 3188
rect 349252 3136 349304 3188
rect 287704 3000 287756 3052
rect 292580 3000 292632 3052
rect 282184 2932 282236 2984
rect 283104 2932 283156 2984
rect 299480 2592 299532 2644
rect 300768 2592 300820 2644
rect 93952 2116 94004 2168
rect 137284 2116 137336 2168
rect 7656 2048 7708 2100
rect 33784 2048 33836 2100
rect 51356 2048 51408 2100
rect 97264 2048 97316 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702574 8156 703520
rect 24320 702642 24348 703520
rect 24308 702636 24360 702642
rect 24308 702578 24360 702584
rect 8116 702568 8168 702574
rect 8116 702510 8168 702516
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 33784 683188 33836 683194
rect 33784 683130 33836 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 15844 670744 15896 670750
rect 15844 670686 15896 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3332 580984 3384 580990
rect 3332 580926 3384 580932
rect 3344 580009 3372 580926
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3436 576842 3464 632023
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618662 3556 619103
rect 3516 618656 3568 618662
rect 3516 618598 3568 618604
rect 7564 618656 7616 618662
rect 7564 618598 7616 618604
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 576836 3476 576842
rect 3424 576778 3476 576784
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 2778 553888 2834 553897
rect 2778 553823 2780 553832
rect 2832 553823 2834 553832
rect 2780 553794 2832 553800
rect 3436 536110 3464 566879
rect 4804 553852 4856 553858
rect 4804 553794 4856 553800
rect 4816 538218 4844 553794
rect 7576 540258 7604 618598
rect 15856 541113 15884 670686
rect 33796 543046 33824 683130
rect 36544 656940 36596 656946
rect 36544 656882 36596 656888
rect 36556 589966 36584 656882
rect 36544 589960 36596 589966
rect 36544 589902 36596 589908
rect 40052 589286 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299584 703582 299980 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 67640 702500 67692 702506
rect 67640 702442 67692 702448
rect 62028 700392 62080 700398
rect 62028 700334 62080 700340
rect 40040 589280 40092 589286
rect 40040 589222 40092 589228
rect 55034 582584 55090 582593
rect 55034 582519 55090 582528
rect 53748 579692 53800 579698
rect 53748 579634 53800 579640
rect 52368 565888 52420 565894
rect 52368 565830 52420 565836
rect 39948 564460 40000 564466
rect 39948 564402 40000 564408
rect 33784 543040 33836 543046
rect 33784 542982 33836 542988
rect 15842 541104 15898 541113
rect 15842 541039 15898 541048
rect 7564 540252 7616 540258
rect 7564 540194 7616 540200
rect 4804 538212 4856 538218
rect 4804 538154 4856 538160
rect 3424 536104 3476 536110
rect 3424 536046 3476 536052
rect 3148 528556 3200 528562
rect 3148 528498 3200 528504
rect 3160 527921 3188 528498
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 3424 522300 3476 522306
rect 3424 522242 3476 522248
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 2780 514762 2832 514768
rect 3436 501809 3464 522242
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 475386 3372 475623
rect 3332 475380 3384 475386
rect 3332 475322 3384 475328
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3436 462466 3464 462567
rect 3424 462460 3476 462466
rect 3424 462402 3476 462408
rect 4816 450566 4844 514762
rect 7564 462460 7616 462466
rect 7564 462402 7616 462408
rect 4804 450560 4856 450566
rect 4804 450502 4856 450508
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3424 434852 3476 434858
rect 3424 434794 3476 434800
rect 3436 423609 3464 434794
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3514 410544 3570 410553
rect 3514 410479 3570 410488
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 377369 3464 397423
rect 3528 389230 3556 410479
rect 4804 397520 4856 397526
rect 4804 397462 4856 397468
rect 3516 389224 3568 389230
rect 3516 389166 3568 389172
rect 3516 383716 3568 383722
rect 3516 383658 3568 383664
rect 3422 377360 3478 377369
rect 3422 377295 3478 377304
rect 3528 371385 3556 383658
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 4816 358494 4844 397462
rect 7576 391921 7604 462402
rect 36544 448588 36596 448594
rect 36544 448530 36596 448536
rect 7562 391912 7618 391921
rect 7562 391847 7618 391856
rect 36556 389298 36584 448530
rect 39856 409148 39908 409154
rect 39856 409090 39908 409096
rect 36544 389292 36596 389298
rect 36544 389234 36596 389240
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 4804 358488 4856 358494
rect 2832 358456 2834 358465
rect 4804 358430 4856 358436
rect 2778 358391 2834 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 19338 342952 19394 342961
rect 19338 342887 19394 342896
rect 8298 336016 8354 336025
rect 8298 335951 8354 335960
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3424 306332 3476 306338
rect 3424 306274 3476 306280
rect 3436 306241 3464 306274
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3422 290456 3478 290465
rect 3422 290391 3478 290400
rect 3436 267209 3464 290391
rect 4080 279478 4108 319223
rect 5538 300112 5594 300121
rect 5538 300047 5594 300056
rect 4158 294536 4214 294545
rect 4158 294471 4214 294480
rect 4068 279472 4120 279478
rect 4068 279414 4120 279420
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3436 254153 3464 255206
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 242208 3476 242214
rect 3424 242150 3476 242156
rect 3436 241097 3464 242150
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3424 229220 3476 229226
rect 3424 229162 3476 229168
rect 2778 215928 2834 215937
rect 2778 215863 2834 215872
rect 112 14544 164 14550
rect 112 14486 164 14492
rect 124 490 152 14486
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 8978
rect 2792 3534 2820 215863
rect 3436 188873 3464 229162
rect 3514 214976 3570 214985
rect 3514 214911 3516 214920
rect 3568 214911 3570 214920
rect 3516 214882 3568 214888
rect 3516 202156 3568 202162
rect 3516 202098 3568 202104
rect 3528 201929 3556 202098
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3436 146266 3464 162823
rect 3424 146260 3476 146266
rect 3424 146202 3476 146208
rect 2872 137964 2924 137970
rect 2872 137906 2924 137912
rect 2884 136785 2912 137906
rect 2870 136776 2926 136785
rect 2870 136711 2926 136720
rect 3424 134564 3476 134570
rect 3424 134506 3476 134512
rect 2872 110832 2924 110838
rect 2872 110774 2924 110780
rect 2884 110673 2912 110774
rect 2870 110664 2926 110673
rect 2870 110599 2926 110608
rect 3054 97608 3110 97617
rect 3054 97543 3110 97552
rect 3068 96694 3096 97543
rect 3056 96688 3108 96694
rect 3056 96630 3108 96636
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 3436 58585 3464 134506
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 2872 50380 2924 50386
rect 2872 50322 2924 50328
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 50322
rect 3516 46232 3568 46238
rect 3516 46174 3568 46180
rect 3528 45529 3556 46174
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 294471
rect 4250 149832 4306 149841
rect 4250 149767 4306 149776
rect 4264 146946 4292 149767
rect 4252 146940 4304 146946
rect 4252 146882 4304 146888
rect 4804 135312 4856 135318
rect 4804 135254 4856 135260
rect 4816 110838 4844 135254
rect 4804 110832 4856 110838
rect 4804 110774 4856 110780
rect 5552 16574 5580 300047
rect 7564 261520 7616 261526
rect 7564 261462 7616 261468
rect 7576 214946 7604 261462
rect 7564 214940 7616 214946
rect 7564 214882 7616 214888
rect 7576 113830 7604 214882
rect 7564 113824 7616 113830
rect 7564 113766 7616 113772
rect 7564 106956 7616 106962
rect 7564 106898 7616 106904
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 480 4108 3470
rect 5276 480 5304 16546
rect 6012 490 6040 16546
rect 7576 6866 7604 106898
rect 8312 16574 8340 335951
rect 12438 334656 12494 334665
rect 12438 334591 12494 334600
rect 11058 298752 11114 298761
rect 11058 298687 11114 298696
rect 9680 186992 9732 186998
rect 9680 186934 9732 186940
rect 9692 16574 9720 186934
rect 8312 16546 8800 16574
rect 9692 16546 9996 16574
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 6288 598 6500 626
rect 6288 490 6316 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 462 6316 490
rect 6472 480 6500 598
rect 7668 480 7696 2042
rect 8772 480 8800 16546
rect 9968 480 9996 16546
rect 11072 6914 11100 298687
rect 11150 25528 11206 25537
rect 11150 25463 11206 25472
rect 11164 16574 11192 25463
rect 12452 16574 12480 334591
rect 16578 330440 16634 330449
rect 16578 330375 16634 330384
rect 15198 320784 15254 320793
rect 15198 320719 15254 320728
rect 14464 292596 14516 292602
rect 14464 292538 14516 292544
rect 14476 241466 14504 292538
rect 14464 241460 14516 241466
rect 14464 241402 14516 241408
rect 13818 236056 13874 236065
rect 13818 235991 13874 236000
rect 13832 16574 13860 235991
rect 15212 16574 15240 320719
rect 16592 16574 16620 330375
rect 17958 302288 18014 302297
rect 17958 302223 18014 302232
rect 17972 16574 18000 302223
rect 19352 16574 19380 342887
rect 33140 338768 33192 338774
rect 33140 338710 33192 338716
rect 30380 333260 30432 333266
rect 30380 333202 30432 333208
rect 20718 331800 20774 331809
rect 20718 331735 20774 331744
rect 20732 16574 20760 331735
rect 22098 327176 22154 327185
rect 22098 327111 22154 327120
rect 22112 16574 22140 327111
rect 26238 323640 26294 323649
rect 26238 323575 26294 323584
rect 24858 291816 24914 291825
rect 24858 291751 24914 291760
rect 22744 262268 22796 262274
rect 22744 262210 22796 262216
rect 22756 242214 22784 262210
rect 22744 242208 22796 242214
rect 22744 242150 22796 242156
rect 22742 235240 22798 235249
rect 22742 235175 22798 235184
rect 11164 16546 11928 16574
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 17972 16546 18276 16574
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 11072 6886 11192 6914
rect 11164 480 11192 6886
rect 11900 490 11928 16546
rect 12176 598 12388 626
rect 12176 490 12204 598
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 11900 462 12204 490
rect 12360 480 12388 598
rect 13556 480 13584 16546
rect 14292 490 14320 16546
rect 14568 598 14780 626
rect 14568 490 14596 598
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 462 14596 490
rect 14752 480 14780 598
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 18248 480 18276 16546
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 480 19472 3470
rect 20180 490 20208 16546
rect 20456 598 20668 626
rect 20456 490 20484 598
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 462 20484 490
rect 20640 480 20668 598
rect 21836 480 21864 16546
rect 22572 490 22600 16546
rect 22756 3534 22784 235175
rect 23480 33788 23532 33794
rect 23480 33730 23532 33736
rect 23492 16574 23520 33730
rect 24872 16574 24900 291751
rect 26252 16574 26280 323575
rect 28998 301472 29054 301481
rect 28998 301407 29054 301416
rect 27618 297392 27674 297401
rect 27618 297327 27674 297336
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 26252 16546 26556 16574
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22848 598 23060 626
rect 22848 490 22876 598
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 462 22876 490
rect 23032 480 23060 598
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 26528 480 26556 16546
rect 27632 6914 27660 297327
rect 27710 152416 27766 152425
rect 27710 152351 27766 152360
rect 27724 16574 27752 152351
rect 29012 16574 29040 301407
rect 30392 16574 30420 333202
rect 31760 198008 31812 198014
rect 31760 197950 31812 197956
rect 31772 16574 31800 197950
rect 33152 16574 33180 338710
rect 34518 328536 34574 328545
rect 34518 328471 34574 328480
rect 34428 316736 34480 316742
rect 34428 316678 34480 316684
rect 34440 306338 34468 316678
rect 34428 306332 34480 306338
rect 34428 306274 34480 306280
rect 34440 305046 34468 306274
rect 34428 305040 34480 305046
rect 34428 304982 34480 304988
rect 33784 182844 33836 182850
rect 33784 182786 33836 182792
rect 27724 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 28460 490 28488 16546
rect 28736 598 28948 626
rect 28736 490 28764 598
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28460 462 28764 490
rect 28920 480 28948 598
rect 30116 480 30144 16546
rect 30852 490 30880 16546
rect 31128 598 31340 626
rect 31128 490 31156 598
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 462 31156 490
rect 31312 480 31340 598
rect 31956 490 31984 16546
rect 32232 598 32444 626
rect 32232 490 32260 598
rect 31270 -960 31382 480
rect 31956 462 32260 490
rect 32416 480 32444 598
rect 33612 480 33640 16546
rect 33796 2106 33824 182786
rect 34532 16574 34560 328471
rect 35900 322380 35952 322386
rect 35900 322322 35952 322328
rect 35164 305040 35216 305046
rect 35164 304982 35216 304988
rect 35176 253230 35204 304982
rect 35164 253224 35216 253230
rect 35164 253166 35216 253172
rect 34532 16546 34836 16574
rect 33784 2100 33836 2106
rect 33784 2042 33836 2048
rect 34808 480 34836 16546
rect 35912 3534 35940 322322
rect 39868 257378 39896 409090
rect 39960 389201 39988 564402
rect 50988 543788 51040 543794
rect 50988 543730 51040 543736
rect 43444 538348 43496 538354
rect 43444 538290 43496 538296
rect 41328 536104 41380 536110
rect 41328 536046 41380 536052
rect 41236 436144 41288 436150
rect 41236 436086 41288 436092
rect 39946 389192 40002 389201
rect 39946 389127 40002 389136
rect 41248 324358 41276 436086
rect 41340 396778 41368 536046
rect 43456 475386 43484 538290
rect 48136 534744 48188 534750
rect 48136 534686 48188 534692
rect 43444 475380 43496 475386
rect 43444 475322 43496 475328
rect 42706 437608 42762 437617
rect 42706 437543 42762 437552
rect 41328 396772 41380 396778
rect 41328 396714 41380 396720
rect 42720 346390 42748 437543
rect 43456 391270 43484 475322
rect 44088 422952 44140 422958
rect 44088 422894 44140 422900
rect 43444 391264 43496 391270
rect 43444 391206 43496 391212
rect 42708 346384 42760 346390
rect 42708 346326 42760 346332
rect 42720 345914 42748 346326
rect 42708 345908 42760 345914
rect 42708 345850 42760 345856
rect 43444 345908 43496 345914
rect 43444 345850 43496 345856
rect 41326 337376 41382 337385
rect 41326 337311 41382 337320
rect 41236 324352 41288 324358
rect 41236 324294 41288 324300
rect 41248 319462 41276 324294
rect 41236 319456 41288 319462
rect 41236 319398 41288 319404
rect 40040 315308 40092 315314
rect 40040 315250 40092 315256
rect 39856 257372 39908 257378
rect 39856 257314 39908 257320
rect 38658 233880 38714 233889
rect 38658 233815 38714 233824
rect 35990 202192 36046 202201
rect 35990 202127 36046 202136
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 202127
rect 37280 196648 37332 196654
rect 37280 196590 37332 196596
rect 37292 16574 37320 196590
rect 38672 16574 38700 233815
rect 40052 16574 40080 315250
rect 41340 131782 41368 337311
rect 41418 325816 41474 325825
rect 41418 325751 41474 325760
rect 41328 131776 41380 131782
rect 41328 131718 41380 131724
rect 41432 16574 41460 325751
rect 43456 287706 43484 345850
rect 43444 287700 43496 287706
rect 43444 287642 43496 287648
rect 43444 280220 43496 280226
rect 43444 280162 43496 280168
rect 43456 255270 43484 280162
rect 43996 269816 44048 269822
rect 43996 269758 44048 269764
rect 43444 255264 43496 255270
rect 43444 255206 43496 255212
rect 44008 149161 44036 269758
rect 44100 267034 44128 422894
rect 48148 407794 48176 534686
rect 51000 513330 51028 543730
rect 50988 513324 51040 513330
rect 50988 513266 51040 513272
rect 51000 439550 51028 513266
rect 52380 456929 52408 565830
rect 52366 456920 52422 456929
rect 52366 456855 52422 456864
rect 50988 439544 51040 439550
rect 50988 439486 51040 439492
rect 52276 436212 52328 436218
rect 52276 436154 52328 436160
rect 48228 429208 48280 429214
rect 48228 429150 48280 429156
rect 48136 407788 48188 407794
rect 48136 407730 48188 407736
rect 48148 380866 48176 407730
rect 48136 380860 48188 380866
rect 48136 380802 48188 380808
rect 44272 318096 44324 318102
rect 44272 318038 44324 318044
rect 44088 267028 44140 267034
rect 44088 266970 44140 266976
rect 44088 200796 44140 200802
rect 44088 200738 44140 200744
rect 43994 149152 44050 149161
rect 43994 149087 44050 149096
rect 44008 120737 44036 149087
rect 43994 120728 44050 120737
rect 43994 120663 44050 120672
rect 42800 35216 42852 35222
rect 42800 35158 42852 35164
rect 42812 16574 42840 35158
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 42812 16546 43116 16574
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 37200 480 37228 3470
rect 38396 480 38424 16546
rect 39132 490 39160 16546
rect 39408 598 39620 626
rect 39408 490 39436 598
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 462 39436 490
rect 39592 480 39620 598
rect 40236 490 40264 16546
rect 40512 598 40724 626
rect 40512 490 40540 598
rect 39550 -960 39662 480
rect 40236 462 40540 490
rect 40696 480 40724 598
rect 41892 480 41920 16546
rect 43088 480 43116 16546
rect 44100 3482 44128 200738
rect 44284 16574 44312 318038
rect 46846 285832 46902 285841
rect 46846 285767 46902 285776
rect 46860 140078 46888 285767
rect 48148 254590 48176 380802
rect 48240 272542 48268 429150
rect 49608 425740 49660 425746
rect 49608 425682 49660 425688
rect 48228 272536 48280 272542
rect 48228 272478 48280 272484
rect 49516 271176 49568 271182
rect 49516 271118 49568 271124
rect 48228 259480 48280 259486
rect 48228 259422 48280 259428
rect 48136 254584 48188 254590
rect 48136 254526 48188 254532
rect 46848 140072 46900 140078
rect 46848 140014 46900 140020
rect 48148 105602 48176 254526
rect 48240 109070 48268 259422
rect 49528 153270 49556 271118
rect 49620 268433 49648 425682
rect 50988 420980 51040 420986
rect 50988 420922 51040 420928
rect 50896 406428 50948 406434
rect 50896 406370 50948 406376
rect 50802 387696 50858 387705
rect 50802 387631 50858 387640
rect 49606 268424 49662 268433
rect 49606 268359 49662 268368
rect 50816 265033 50844 387631
rect 50802 265024 50858 265033
rect 50802 264959 50858 264968
rect 50908 256018 50936 406370
rect 51000 387705 51028 420922
rect 52184 411936 52236 411942
rect 52184 411878 52236 411884
rect 50986 387696 51042 387705
rect 50986 387631 51042 387640
rect 52092 286340 52144 286346
rect 52092 286282 52144 286288
rect 50988 284436 51040 284442
rect 50988 284378 51040 284384
rect 50896 256012 50948 256018
rect 50896 255954 50948 255960
rect 50894 239456 50950 239465
rect 50894 239391 50950 239400
rect 49606 237960 49662 237969
rect 49606 237895 49662 237904
rect 49516 153264 49568 153270
rect 49516 153206 49568 153212
rect 48320 131776 48372 131782
rect 48320 131718 48372 131724
rect 48228 109064 48280 109070
rect 48228 109006 48280 109012
rect 48136 105596 48188 105602
rect 48136 105538 48188 105544
rect 46940 54528 46992 54534
rect 46940 54470 46992 54476
rect 45560 36576 45612 36582
rect 45560 36518 45612 36524
rect 45572 16574 45600 36518
rect 46952 16574 46980 54470
rect 48332 16574 48360 131718
rect 49528 120086 49556 153206
rect 49516 120080 49568 120086
rect 49516 120022 49568 120028
rect 49620 89690 49648 237895
rect 50908 211138 50936 239391
rect 50896 211132 50948 211138
rect 50896 211074 50948 211080
rect 50908 92410 50936 211074
rect 51000 132462 51028 284378
rect 52104 138718 52132 286282
rect 52196 258738 52224 411878
rect 52288 309126 52316 436154
rect 52380 409154 52408 456855
rect 53470 434752 53526 434761
rect 53470 434687 53526 434696
rect 52368 409148 52420 409154
rect 52368 409090 52420 409096
rect 52276 309120 52328 309126
rect 52276 309062 52328 309068
rect 52288 277370 52316 309062
rect 52460 279472 52512 279478
rect 52460 279414 52512 279420
rect 52472 278798 52500 279414
rect 52460 278792 52512 278798
rect 52460 278734 52512 278740
rect 53484 278730 53512 434687
rect 53760 433362 53788 579634
rect 53748 433356 53800 433362
rect 53748 433298 53800 433304
rect 54852 414044 54904 414050
rect 54852 413986 54904 413992
rect 54760 403028 54812 403034
rect 54760 402970 54812 402976
rect 53656 398880 53708 398886
rect 53656 398822 53708 398828
rect 53564 278792 53616 278798
rect 53564 278734 53616 278740
rect 53472 278724 53524 278730
rect 53472 278666 53524 278672
rect 52276 277364 52328 277370
rect 52276 277306 52328 277312
rect 52184 258732 52236 258738
rect 52184 258674 52236 258680
rect 52460 257372 52512 257378
rect 52460 257314 52512 257320
rect 52472 256766 52500 257314
rect 52460 256760 52512 256766
rect 52460 256702 52512 256708
rect 53472 256760 53524 256766
rect 53472 256702 53524 256708
rect 52368 242956 52420 242962
rect 52368 242898 52420 242904
rect 52380 214577 52408 242898
rect 52366 214568 52422 214577
rect 52366 214503 52422 214512
rect 52184 179444 52236 179450
rect 52184 179386 52236 179392
rect 52092 138712 52144 138718
rect 52092 138654 52144 138660
rect 50988 132456 51040 132462
rect 50988 132398 51040 132404
rect 52196 125594 52224 179386
rect 52184 125588 52236 125594
rect 52184 125530 52236 125536
rect 52380 95198 52408 214503
rect 53484 200122 53512 256702
rect 53472 200116 53524 200122
rect 53472 200058 53524 200064
rect 53484 198762 53512 200058
rect 53472 198756 53524 198762
rect 53472 198698 53524 198704
rect 53576 156670 53604 278734
rect 53668 249082 53696 398822
rect 54772 251870 54800 402970
rect 54864 262886 54892 413986
rect 55048 411942 55076 582519
rect 55128 578264 55180 578270
rect 55128 578206 55180 578212
rect 55036 411936 55088 411942
rect 55036 411878 55088 411884
rect 55140 402966 55168 578206
rect 60648 571396 60700 571402
rect 60648 571338 60700 571344
rect 57888 569968 57940 569974
rect 57888 569910 57940 569916
rect 57796 553444 57848 553450
rect 57796 553386 57848 553392
rect 57704 433356 57756 433362
rect 57704 433298 57756 433304
rect 56508 431248 56560 431254
rect 56508 431190 56560 431196
rect 55128 402960 55180 402966
rect 55128 402902 55180 402908
rect 56416 288448 56468 288454
rect 56416 288390 56468 288396
rect 56232 275324 56284 275330
rect 56232 275266 56284 275272
rect 54944 267096 54996 267102
rect 54944 267038 54996 267044
rect 54852 262880 54904 262886
rect 54852 262822 54904 262828
rect 54760 251864 54812 251870
rect 54760 251806 54812 251812
rect 53656 249076 53708 249082
rect 53656 249018 53708 249024
rect 53748 241528 53800 241534
rect 53748 241470 53800 241476
rect 53656 198756 53708 198762
rect 53656 198698 53708 198704
rect 53564 156664 53616 156670
rect 53564 156606 53616 156612
rect 52460 148368 52512 148374
rect 52460 148310 52512 148316
rect 52368 95192 52420 95198
rect 52368 95134 52420 95140
rect 50896 92404 50948 92410
rect 50896 92346 50948 92352
rect 49608 89684 49660 89690
rect 49608 89626 49660 89632
rect 52368 85536 52420 85542
rect 52368 85478 52420 85484
rect 52380 84250 52408 85478
rect 52368 84244 52420 84250
rect 52368 84186 52420 84192
rect 52380 81394 52408 84186
rect 52368 81388 52420 81394
rect 52368 81330 52420 81336
rect 49700 17264 49752 17270
rect 49700 17206 49752 17212
rect 49712 16574 49740 17206
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44100 3454 44312 3482
rect 44284 480 44312 3454
rect 45020 490 45048 16546
rect 45296 598 45508 626
rect 45296 490 45324 598
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 462 45324 490
rect 45480 480 45508 598
rect 46676 480 46704 16546
rect 47412 490 47440 16546
rect 47688 598 47900 626
rect 47688 490 47716 598
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 462 47716 490
rect 47872 480 47900 598
rect 48516 490 48544 16546
rect 48792 598 49004 626
rect 48792 490 48820 598
rect 47830 -960 47942 480
rect 48516 462 48820 490
rect 48976 480 49004 598
rect 50172 480 50200 16546
rect 52472 6914 52500 148310
rect 53668 143614 53696 198698
rect 53656 143608 53708 143614
rect 53656 143550 53708 143556
rect 52552 109064 52604 109070
rect 52552 109006 52604 109012
rect 52564 85542 52592 109006
rect 53668 109002 53696 143550
rect 53656 108996 53708 109002
rect 53656 108938 53708 108944
rect 53760 93838 53788 241470
rect 54956 151842 54984 267038
rect 55036 260160 55088 260166
rect 55036 260102 55088 260108
rect 54944 151836 54996 151842
rect 54944 151778 54996 151784
rect 54956 117230 54984 151778
rect 55048 146985 55076 260102
rect 56244 155922 56272 275266
rect 56322 254144 56378 254153
rect 56322 254079 56378 254088
rect 56336 229094 56364 254079
rect 56428 239426 56456 288390
rect 56520 273358 56548 431190
rect 57610 425640 57666 425649
rect 57610 425575 57666 425584
rect 56508 273352 56560 273358
rect 56508 273294 56560 273300
rect 57624 270502 57652 425575
rect 57716 310457 57744 433298
rect 57808 416838 57836 553386
rect 57900 449206 57928 569910
rect 59084 539640 59136 539646
rect 59084 539582 59136 539588
rect 57888 449200 57940 449206
rect 57888 449142 57940 449148
rect 57900 420238 57928 449142
rect 57888 420232 57940 420238
rect 57888 420174 57940 420180
rect 57796 416832 57848 416838
rect 57796 416774 57848 416780
rect 57980 413296 58032 413302
rect 57980 413238 58032 413244
rect 57992 411942 58020 413238
rect 57980 411936 58032 411942
rect 57980 411878 58032 411884
rect 58992 400240 59044 400246
rect 58992 400182 59044 400188
rect 57702 310448 57758 310457
rect 57702 310383 57758 310392
rect 57716 306374 57744 310383
rect 57716 306346 57836 306374
rect 57702 283112 57758 283121
rect 57702 283047 57758 283056
rect 57612 270496 57664 270502
rect 57612 270438 57664 270444
rect 56508 256012 56560 256018
rect 56508 255954 56560 255960
rect 56520 254153 56548 255954
rect 56506 254144 56562 254153
rect 56506 254079 56562 254088
rect 56416 239420 56468 239426
rect 56416 239362 56468 239368
rect 56336 229066 56456 229094
rect 56428 218657 56456 229066
rect 56414 218648 56470 218657
rect 56414 218583 56470 218592
rect 56232 155916 56284 155922
rect 56232 155858 56284 155864
rect 55034 146976 55090 146985
rect 55034 146911 55090 146920
rect 55048 142154 55076 146911
rect 55048 142126 55168 142154
rect 54944 117224 54996 117230
rect 54944 117166 54996 117172
rect 55140 111790 55168 142126
rect 55128 111784 55180 111790
rect 55128 111726 55180 111732
rect 56428 104854 56456 218583
rect 57716 173194 57744 283047
rect 57808 274825 57836 306346
rect 59004 283014 59032 400182
rect 59096 391513 59124 539582
rect 59176 536852 59228 536858
rect 59176 536794 59228 536800
rect 59082 391504 59138 391513
rect 59082 391439 59138 391448
rect 59188 388482 59216 536794
rect 60660 524414 60688 571338
rect 61936 558952 61988 558958
rect 61936 558894 61988 558900
rect 60648 524408 60700 524414
rect 60648 524350 60700 524356
rect 60554 519480 60610 519489
rect 60554 519415 60610 519424
rect 59268 423700 59320 423706
rect 59268 423642 59320 423648
rect 59176 388476 59228 388482
rect 59176 388418 59228 388424
rect 58992 283008 59044 283014
rect 58992 282950 59044 282956
rect 57794 274816 57850 274825
rect 57794 274751 57850 274760
rect 57888 270496 57940 270502
rect 57888 270438 57940 270444
rect 57900 269822 57928 270438
rect 57888 269816 57940 269822
rect 57888 269758 57940 269764
rect 57796 268388 57848 268394
rect 57796 268330 57848 268336
rect 57704 173188 57756 173194
rect 57704 173130 57756 173136
rect 56508 155916 56560 155922
rect 56508 155858 56560 155864
rect 56520 154698 56548 155858
rect 56508 154692 56560 154698
rect 56508 154634 56560 154640
rect 56520 124914 56548 154634
rect 57242 135960 57298 135969
rect 57242 135895 57298 135904
rect 56508 124908 56560 124914
rect 56508 124850 56560 124856
rect 56416 104848 56468 104854
rect 56416 104790 56468 104796
rect 53748 93832 53800 93838
rect 53748 93774 53800 93780
rect 52552 85536 52604 85542
rect 52552 85478 52604 85484
rect 52550 77888 52606 77897
rect 52550 77823 52606 77832
rect 52564 16574 52592 77823
rect 53840 47592 53892 47598
rect 53840 47534 53892 47540
rect 53852 16574 53880 47534
rect 56598 40624 56654 40633
rect 56598 40559 56654 40568
rect 55220 32428 55272 32434
rect 55220 32370 55272 32376
rect 55232 16574 55260 32370
rect 56612 16574 56640 40559
rect 57256 33114 57284 135895
rect 57716 132394 57744 173130
rect 57808 151094 57836 268330
rect 58348 267028 58400 267034
rect 58348 266970 58400 266976
rect 58360 266529 58388 266970
rect 58346 266520 58402 266529
rect 58346 266455 58402 266464
rect 57886 265024 57942 265033
rect 57886 264959 57942 264968
rect 57796 151088 57848 151094
rect 57796 151030 57848 151036
rect 57704 132388 57756 132394
rect 57704 132330 57756 132336
rect 57808 118658 57836 151030
rect 57900 147694 57928 264959
rect 59004 250578 59032 282950
rect 59084 272536 59136 272542
rect 59084 272478 59136 272484
rect 59096 271969 59124 272478
rect 59082 271960 59138 271969
rect 59082 271895 59138 271904
rect 58992 250572 59044 250578
rect 58992 250514 59044 250520
rect 59096 160721 59124 271895
rect 59280 268394 59308 423642
rect 60004 410576 60056 410582
rect 60004 410518 60056 410524
rect 60016 409154 60044 410518
rect 60004 409148 60056 409154
rect 60004 409090 60056 409096
rect 60568 393378 60596 519415
rect 60646 443048 60702 443057
rect 60646 442983 60702 442992
rect 60556 393372 60608 393378
rect 60556 393314 60608 393320
rect 60556 392012 60608 392018
rect 60556 391954 60608 391960
rect 60568 364334 60596 391954
rect 60476 364306 60596 364334
rect 60372 285728 60424 285734
rect 60372 285670 60424 285676
rect 59268 268388 59320 268394
rect 59268 268330 59320 268336
rect 59174 266520 59230 266529
rect 59174 266455 59230 266464
rect 59188 220182 59216 266455
rect 59268 263628 59320 263634
rect 59268 263570 59320 263576
rect 59176 220176 59228 220182
rect 59176 220118 59228 220124
rect 59176 209092 59228 209098
rect 59176 209034 59228 209040
rect 59082 160712 59138 160721
rect 59082 160647 59138 160656
rect 57888 147688 57940 147694
rect 57888 147630 57940 147636
rect 57796 118652 57848 118658
rect 57796 118594 57848 118600
rect 57900 115938 57928 147630
rect 58992 140820 59044 140826
rect 58992 140762 59044 140768
rect 57888 115932 57940 115938
rect 57888 115874 57940 115880
rect 59004 114510 59032 140762
rect 59096 122806 59124 160647
rect 59084 122800 59136 122806
rect 59084 122742 59136 122748
rect 58992 114504 59044 114510
rect 58992 114446 59044 114452
rect 59188 94489 59216 209034
rect 59280 140826 59308 263570
rect 60384 231130 60412 285670
rect 60476 245585 60504 364306
rect 60568 364274 60596 364306
rect 60556 364268 60608 364274
rect 60556 364210 60608 364216
rect 60660 286346 60688 442983
rect 61844 441720 61896 441726
rect 61844 441662 61896 441668
rect 60740 423632 60792 423638
rect 60740 423574 60792 423580
rect 60752 422958 60780 423574
rect 60740 422952 60792 422958
rect 60740 422894 60792 422900
rect 61856 420918 61884 441662
rect 61844 420912 61896 420918
rect 61844 420854 61896 420860
rect 61844 416764 61896 416770
rect 61844 416706 61896 416712
rect 61856 415478 61884 416706
rect 61844 415472 61896 415478
rect 61844 415414 61896 415420
rect 60740 396772 60792 396778
rect 60740 396714 60792 396720
rect 60752 396098 60780 396714
rect 60740 396092 60792 396098
rect 60740 396034 60792 396040
rect 61856 287054 61884 415414
rect 61948 398818 61976 558894
rect 62040 537538 62068 700334
rect 67548 611380 67600 611386
rect 67548 611322 67600 611328
rect 66166 603120 66222 603129
rect 66166 603055 66222 603064
rect 66076 599004 66128 599010
rect 66076 598946 66128 598952
rect 63408 579760 63460 579766
rect 63408 579702 63460 579708
rect 62028 537532 62080 537538
rect 62028 537474 62080 537480
rect 62040 536858 62068 537474
rect 62028 536852 62080 536858
rect 62028 536794 62080 536800
rect 62028 526448 62080 526454
rect 62028 526390 62080 526396
rect 62040 434790 62068 526390
rect 63420 515438 63448 579702
rect 64604 572756 64656 572762
rect 64604 572698 64656 572704
rect 63408 515432 63460 515438
rect 63408 515374 63460 515380
rect 63408 454708 63460 454714
rect 63408 454650 63460 454656
rect 62028 434784 62080 434790
rect 62028 434726 62080 434732
rect 62040 423638 62068 434726
rect 63316 431996 63368 432002
rect 63316 431938 63368 431944
rect 62028 423632 62080 423638
rect 62028 423574 62080 423580
rect 63328 422294 63356 431938
rect 63236 422266 63356 422294
rect 63236 418334 63264 422266
rect 63224 418328 63276 418334
rect 63224 418270 63276 418276
rect 62028 404388 62080 404394
rect 62028 404330 62080 404336
rect 61936 398812 61988 398818
rect 61936 398754 61988 398760
rect 61936 396092 61988 396098
rect 61936 396034 61988 396040
rect 61948 372570 61976 396034
rect 61936 372564 61988 372570
rect 61936 372506 61988 372512
rect 61764 287026 61884 287054
rect 60648 286340 60700 286346
rect 60648 286282 60700 286288
rect 61764 284889 61792 287026
rect 61750 284880 61806 284889
rect 61750 284815 61806 284824
rect 61108 273352 61160 273358
rect 61106 273320 61108 273329
rect 61160 273320 61162 273329
rect 61106 273255 61162 273264
rect 61764 261089 61792 284815
rect 61934 273320 61990 273329
rect 61934 273255 61990 273264
rect 61842 270736 61898 270745
rect 61842 270671 61898 270680
rect 60554 261080 60610 261089
rect 60554 261015 60610 261024
rect 61750 261080 61806 261089
rect 61750 261015 61806 261024
rect 60462 245576 60518 245585
rect 60462 245511 60518 245520
rect 60372 231124 60424 231130
rect 60372 231066 60424 231072
rect 60464 164892 60516 164898
rect 60464 164834 60516 164840
rect 59268 140820 59320 140826
rect 59268 140762 59320 140768
rect 59266 139496 59322 139505
rect 59266 139431 59322 139440
rect 59280 110430 59308 139431
rect 59268 110424 59320 110430
rect 59268 110366 59320 110372
rect 59174 94480 59230 94489
rect 59174 94415 59230 94424
rect 60476 88262 60504 164834
rect 60568 113082 60596 261015
rect 61752 258732 61804 258738
rect 61752 258674 61804 258680
rect 60648 249076 60700 249082
rect 60648 249018 60700 249024
rect 60556 113076 60608 113082
rect 60556 113018 60608 113024
rect 60660 99686 60688 249018
rect 61764 235929 61792 258674
rect 61750 235920 61806 235929
rect 61750 235855 61806 235864
rect 61752 188352 61804 188358
rect 61752 188294 61804 188300
rect 61764 113174 61792 188294
rect 61856 144945 61884 270671
rect 61842 144936 61898 144945
rect 61842 144871 61898 144880
rect 61856 121446 61884 144871
rect 61948 138145 61976 273255
rect 62040 252770 62068 404330
rect 63132 264988 63184 264994
rect 63132 264930 63184 264936
rect 62118 252784 62174 252793
rect 62040 252742 62118 252770
rect 62118 252719 62174 252728
rect 62028 247104 62080 247110
rect 62028 247046 62080 247052
rect 62040 221513 62068 247046
rect 62026 221504 62082 221513
rect 62026 221439 62082 221448
rect 61934 138136 61990 138145
rect 61934 138071 61990 138080
rect 61948 124166 61976 138071
rect 61936 124160 61988 124166
rect 61936 124102 61988 124108
rect 61844 121440 61896 121446
rect 61844 121382 61896 121388
rect 61764 113146 61976 113174
rect 61948 100910 61976 113146
rect 61936 100904 61988 100910
rect 61936 100846 61988 100852
rect 60648 99680 60700 99686
rect 60648 99622 60700 99628
rect 60464 88256 60516 88262
rect 60464 88198 60516 88204
rect 61948 74526 61976 100846
rect 62040 99346 62068 221439
rect 63144 181490 63172 264930
rect 63236 263634 63264 418270
rect 63420 418130 63448 454650
rect 63408 418124 63460 418130
rect 63408 418066 63460 418072
rect 63316 408536 63368 408542
rect 63316 408478 63368 408484
rect 63328 289785 63356 408478
rect 64616 406434 64644 572698
rect 64696 563100 64748 563106
rect 64696 563042 64748 563048
rect 64708 531282 64736 563042
rect 65798 548312 65854 548321
rect 65798 548247 65854 548256
rect 64696 531276 64748 531282
rect 64696 531218 64748 531224
rect 65812 517206 65840 548247
rect 65890 546816 65946 546825
rect 65890 546751 65946 546760
rect 65904 534721 65932 546751
rect 66088 546417 66116 598946
rect 66180 561649 66208 603055
rect 67364 585200 67416 585206
rect 67364 585142 67416 585148
rect 66626 580000 66682 580009
rect 66626 579935 66682 579944
rect 66640 579766 66668 579935
rect 66628 579760 66680 579766
rect 66628 579702 66680 579708
rect 66442 578640 66498 578649
rect 66442 578575 66498 578584
rect 66456 578270 66484 578575
rect 66444 578264 66496 578270
rect 66444 578206 66496 578212
rect 67178 577416 67234 577425
rect 67178 577351 67234 577360
rect 66626 573200 66682 573209
rect 66626 573135 66682 573144
rect 66640 572762 66668 573135
rect 66628 572756 66680 572762
rect 66628 572698 66680 572704
rect 66626 571840 66682 571849
rect 66626 571775 66682 571784
rect 66640 571402 66668 571775
rect 66628 571396 66680 571402
rect 66628 571338 66680 571344
rect 66626 570208 66682 570217
rect 66626 570143 66682 570152
rect 66640 569974 66668 570143
rect 66628 569968 66680 569974
rect 66628 569910 66680 569916
rect 66810 564768 66866 564777
rect 66810 564703 66866 564712
rect 66824 564466 66852 564703
rect 66812 564460 66864 564466
rect 66812 564402 66864 564408
rect 66718 563408 66774 563417
rect 66718 563343 66774 563352
rect 66732 563106 66760 563343
rect 66720 563100 66772 563106
rect 66720 563042 66772 563048
rect 66166 561640 66222 561649
rect 66166 561575 66222 561584
rect 66810 559328 66866 559337
rect 66810 559263 66866 559272
rect 66824 558958 66852 559263
rect 66812 558952 66864 558958
rect 66812 558894 66864 558900
rect 66166 558104 66222 558113
rect 66166 558039 66222 558048
rect 66074 546408 66130 546417
rect 66074 546343 66130 546352
rect 65984 543040 66036 543046
rect 65984 542982 66036 542988
rect 65890 534712 65946 534721
rect 65890 534647 65946 534656
rect 65996 525065 66024 542982
rect 65982 525056 66038 525065
rect 65982 524991 66038 525000
rect 65800 517200 65852 517206
rect 65800 517142 65852 517148
rect 66180 460222 66208 558039
rect 66718 553616 66774 553625
rect 66718 553551 66774 553560
rect 66732 553450 66760 553551
rect 66720 553444 66772 553450
rect 66720 553386 66772 553392
rect 66810 544096 66866 544105
rect 66810 544031 66866 544040
rect 66824 543794 66852 544031
rect 66812 543788 66864 543794
rect 66812 543730 66864 543736
rect 66534 543144 66590 543153
rect 66534 543079 66590 543088
rect 66548 543046 66576 543079
rect 66536 543040 66588 543046
rect 66536 542982 66588 542988
rect 66626 540016 66682 540025
rect 66626 539951 66682 539960
rect 66640 539646 66668 539951
rect 66628 539640 66680 539646
rect 66628 539582 66680 539588
rect 66168 460216 66220 460222
rect 66168 460158 66220 460164
rect 66076 448588 66128 448594
rect 66076 448530 66128 448536
rect 66088 434625 66116 448530
rect 66168 447840 66220 447846
rect 66168 447782 66220 447788
rect 66074 434616 66130 434625
rect 66074 434551 66130 434560
rect 66180 432585 66208 447782
rect 67192 446486 67220 577351
rect 67376 575385 67404 585142
rect 67456 581120 67508 581126
rect 67456 581062 67508 581068
rect 67362 575376 67418 575385
rect 67362 575311 67418 575320
rect 67468 569945 67496 581062
rect 67560 576842 67588 611322
rect 67548 576836 67600 576842
rect 67548 576778 67600 576784
rect 67560 576473 67588 576778
rect 67546 576464 67602 576473
rect 67546 576399 67602 576408
rect 67560 575550 67588 576399
rect 67548 575544 67600 575550
rect 67548 575486 67600 575492
rect 67454 569936 67510 569945
rect 67454 569871 67510 569880
rect 67454 567624 67510 567633
rect 67454 567559 67510 567568
rect 67362 555248 67418 555257
rect 67362 555183 67418 555192
rect 67270 552256 67326 552265
rect 67270 552191 67326 552200
rect 67284 539850 67312 552191
rect 67272 539844 67324 539850
rect 67272 539786 67324 539792
rect 67376 534070 67404 555183
rect 67364 534064 67416 534070
rect 67364 534006 67416 534012
rect 67468 529242 67496 567559
rect 67652 566681 67680 702442
rect 72988 700398 73016 703520
rect 85580 702636 85632 702642
rect 85580 702578 85632 702584
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 84108 700392 84160 700398
rect 84108 700334 84160 700340
rect 71688 700324 71740 700330
rect 71688 700266 71740 700272
rect 69848 593428 69900 593434
rect 69848 593370 69900 593376
rect 69860 581074 69888 593370
rect 71700 585818 71728 700266
rect 71780 612808 71832 612814
rect 71780 612750 71832 612756
rect 71688 585812 71740 585818
rect 71688 585754 71740 585760
rect 71700 585206 71728 585754
rect 71688 585200 71740 585206
rect 71688 585142 71740 585148
rect 71792 581074 71820 612750
rect 79322 599448 79378 599457
rect 79322 599383 79378 599392
rect 77392 590028 77444 590034
rect 77392 589970 77444 589976
rect 74632 589960 74684 589966
rect 74632 589902 74684 589908
rect 73528 583840 73580 583846
rect 73528 583782 73580 583788
rect 73540 581074 73568 583782
rect 74262 581224 74318 581233
rect 74262 581159 74318 581168
rect 74276 581074 74304 581159
rect 69860 581046 70288 581074
rect 71792 581046 72128 581074
rect 73232 581046 73568 581074
rect 74152 581046 74304 581074
rect 74644 581074 74672 589902
rect 77208 582820 77260 582826
rect 77208 582762 77260 582768
rect 76288 582480 76340 582486
rect 76288 582422 76340 582428
rect 75366 581088 75422 581097
rect 74644 581046 75366 581074
rect 76300 581074 76328 582422
rect 77220 581074 77248 582762
rect 75992 581046 76328 581074
rect 76912 581046 77248 581074
rect 77404 581074 77432 589970
rect 79048 583772 79100 583778
rect 79048 583714 79100 583720
rect 79060 581074 79088 583714
rect 79336 582826 79364 599383
rect 84120 590034 84148 700334
rect 85592 596174 85620 702578
rect 89180 700398 89208 703520
rect 96620 702568 96672 702574
rect 96620 702510 96672 702516
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 94688 605872 94740 605878
rect 94688 605814 94740 605820
rect 88982 601896 89038 601905
rect 88982 601831 89038 601840
rect 86960 596216 87012 596222
rect 85592 596146 85896 596174
rect 86960 596158 87012 596164
rect 84108 590028 84160 590034
rect 84108 589970 84160 589976
rect 85488 587920 85540 587926
rect 85488 587862 85540 587868
rect 81808 587172 81860 587178
rect 81808 587114 81860 587120
rect 79324 582820 79376 582826
rect 79324 582762 79376 582768
rect 79966 581224 80022 581233
rect 79966 581159 80022 581168
rect 79980 581074 80008 581159
rect 81820 581074 81848 587114
rect 82726 582720 82782 582729
rect 82726 582655 82782 582664
rect 82740 581074 82768 582655
rect 83002 582584 83058 582593
rect 83002 582519 83058 582528
rect 77404 581046 77832 581074
rect 78752 581046 79088 581074
rect 79672 581046 80008 581074
rect 80256 581058 80928 581074
rect 80244 581052 80928 581058
rect 75366 581023 75422 581032
rect 80296 581046 80928 581052
rect 81512 581046 81848 581074
rect 82432 581046 82768 581074
rect 83016 581074 83044 582519
rect 85500 581074 85528 587862
rect 83016 581046 83352 581074
rect 85376 581046 85528 581074
rect 80244 580994 80296 581000
rect 80900 580825 80928 581046
rect 71502 580816 71558 580825
rect 69032 580774 69368 580802
rect 71208 580774 71502 580802
rect 69032 580718 69060 580774
rect 71502 580751 71558 580760
rect 80886 580816 80942 580825
rect 80886 580751 80942 580760
rect 84198 580816 84254 580825
rect 85868 580802 85896 596146
rect 86972 581074 87000 596158
rect 88996 583438 89024 601831
rect 92480 595468 92532 595474
rect 92480 595410 92532 595416
rect 89720 592068 89772 592074
rect 89720 592010 89772 592016
rect 88248 583432 88300 583438
rect 88248 583374 88300 583380
rect 88984 583432 89036 583438
rect 88984 583374 89036 583380
rect 88260 581074 88288 583374
rect 86972 581046 87216 581074
rect 88136 581046 88288 581074
rect 89732 581074 89760 592010
rect 92112 585200 92164 585206
rect 92112 585142 92164 585148
rect 92124 581074 92152 585142
rect 89732 581046 89976 581074
rect 91816 581046 92152 581074
rect 92492 581074 92520 595410
rect 94412 583432 94464 583438
rect 94412 583374 94464 583380
rect 93768 582412 93820 582418
rect 93768 582354 93820 582360
rect 92492 581046 92736 581074
rect 93780 580938 93808 582354
rect 93656 580910 93808 580938
rect 89258 580816 89314 580825
rect 84254 580774 84456 580802
rect 85868 580774 86632 580802
rect 89056 580774 89258 580802
rect 84198 580751 84254 580760
rect 86604 580718 86632 580774
rect 94424 580802 94452 583374
rect 90896 580774 91048 580802
rect 94424 580774 94576 580802
rect 89258 580751 89314 580760
rect 91020 580718 91048 580774
rect 69020 580712 69072 580718
rect 69020 580654 69072 580660
rect 86592 580712 86644 580718
rect 86592 580654 86644 580660
rect 91008 580712 91060 580718
rect 91008 580654 91060 580660
rect 94700 576094 94728 605814
rect 95148 591320 95200 591326
rect 95148 591262 95200 591268
rect 95160 589286 95188 591262
rect 95148 589280 95200 589286
rect 95148 589222 95200 589228
rect 95160 588962 95188 589222
rect 95160 588934 95372 588962
rect 95148 582480 95200 582486
rect 95148 582422 95200 582428
rect 95160 578950 95188 582422
rect 95148 578944 95200 578950
rect 95148 578886 95200 578892
rect 94688 576088 94740 576094
rect 94688 576030 94740 576036
rect 67824 575544 67876 575550
rect 67824 575486 67876 575492
rect 67638 566672 67694 566681
rect 67638 566607 67694 566616
rect 67652 565894 67680 566607
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67730 562048 67786 562057
rect 67730 561983 67786 561992
rect 67638 556608 67694 556617
rect 67638 556543 67694 556552
rect 67456 529236 67508 529242
rect 67456 529178 67508 529184
rect 67652 461650 67680 556543
rect 67744 469849 67772 561983
rect 67836 527785 67864 575486
rect 95238 563680 95294 563689
rect 95238 563615 95294 563624
rect 94686 558648 94742 558657
rect 94686 558583 94742 558592
rect 73160 539912 73212 539918
rect 73160 539854 73212 539860
rect 94318 539880 94374 539889
rect 71780 539844 71832 539850
rect 71780 539786 71832 539792
rect 68816 539158 68968 539186
rect 68940 536586 68968 539158
rect 69400 539158 69736 539186
rect 70656 539158 70992 539186
rect 68928 536580 68980 536586
rect 68928 536522 68980 536528
rect 69400 536110 69428 539158
rect 70964 538218 70992 539158
rect 71148 539158 71576 539186
rect 70952 538212 71004 538218
rect 70952 538154 71004 538160
rect 70964 536110 70992 538154
rect 69388 536104 69440 536110
rect 69388 536046 69440 536052
rect 70952 536104 71004 536110
rect 70952 536046 71004 536052
rect 71148 528554 71176 539158
rect 70504 528526 71176 528554
rect 67822 527776 67878 527785
rect 67822 527711 67878 527720
rect 68926 525056 68982 525065
rect 68926 524991 68982 525000
rect 67730 469840 67786 469849
rect 67730 469775 67786 469784
rect 68940 466478 68968 524991
rect 69664 517200 69716 517206
rect 69664 517142 69716 517148
rect 68928 466472 68980 466478
rect 68928 466414 68980 466420
rect 67640 461644 67692 461650
rect 67640 461586 67692 461592
rect 67180 446480 67232 446486
rect 67180 446422 67232 446428
rect 67192 441614 67220 446422
rect 68940 443698 68968 466414
rect 69676 448497 69704 517142
rect 70504 448594 70532 528526
rect 70492 448588 70544 448594
rect 70492 448530 70544 448536
rect 69662 448488 69718 448497
rect 69662 448423 69718 448432
rect 68928 443692 68980 443698
rect 68928 443634 68980 443640
rect 68284 441652 68336 441658
rect 67192 441586 67496 441614
rect 68284 441594 68336 441600
rect 69676 441614 69704 448423
rect 71136 443012 71188 443018
rect 71136 442954 71188 442960
rect 67364 438184 67416 438190
rect 67364 438126 67416 438132
rect 67272 433832 67324 433838
rect 67272 433774 67324 433780
rect 66810 433392 66866 433401
rect 66810 433327 66812 433336
rect 66864 433327 66866 433336
rect 66812 433298 66864 433304
rect 66166 432576 66222 432585
rect 65708 432540 65760 432546
rect 66166 432511 66168 432520
rect 65708 432482 65760 432488
rect 66220 432511 66222 432520
rect 66168 432482 66220 432488
rect 64696 429412 64748 429418
rect 64696 429354 64748 429360
rect 64604 406428 64656 406434
rect 64604 406370 64656 406376
rect 64604 397520 64656 397526
rect 64604 397462 64656 397468
rect 64616 375329 64644 397462
rect 64602 375320 64658 375329
rect 64602 375255 64658 375264
rect 63314 289776 63370 289785
rect 63314 289711 63370 289720
rect 63328 267734 63356 289711
rect 64602 287736 64658 287745
rect 64602 287671 64658 287680
rect 63328 267706 63448 267734
rect 63224 263628 63276 263634
rect 63224 263570 63276 263576
rect 63224 262268 63276 262274
rect 63224 262210 63276 262216
rect 63236 229770 63264 262210
rect 63420 255377 63448 267706
rect 64616 259418 64644 287671
rect 64708 273290 64736 429354
rect 64788 411324 64840 411330
rect 64788 411266 64840 411272
rect 64800 287745 64828 411266
rect 64786 287736 64842 287745
rect 64786 287671 64842 287680
rect 64786 283384 64842 283393
rect 64786 283319 64842 283328
rect 64696 273284 64748 273290
rect 64696 273226 64748 273232
rect 64604 259412 64656 259418
rect 64604 259354 64656 259360
rect 63406 255368 63462 255377
rect 63406 255303 63462 255312
rect 63406 252784 63462 252793
rect 63406 252719 63462 252728
rect 63224 229764 63276 229770
rect 63224 229706 63276 229712
rect 63132 181484 63184 181490
rect 63132 181426 63184 181432
rect 63144 180794 63172 181426
rect 63144 180766 63356 180794
rect 63224 166320 63276 166326
rect 63224 166262 63276 166268
rect 63132 140140 63184 140146
rect 63132 140082 63184 140088
rect 63144 113150 63172 140082
rect 63236 128314 63264 166262
rect 63224 128308 63276 128314
rect 63224 128250 63276 128256
rect 63328 115326 63356 180766
rect 63316 115320 63368 115326
rect 63316 115262 63368 115268
rect 63132 113144 63184 113150
rect 63132 113086 63184 113092
rect 63420 102270 63448 252719
rect 63500 251864 63552 251870
rect 63500 251806 63552 251812
rect 63512 251326 63540 251806
rect 63500 251320 63552 251326
rect 63500 251262 63552 251268
rect 64696 251320 64748 251326
rect 64696 251262 64748 251268
rect 64604 160132 64656 160138
rect 64604 160074 64656 160080
rect 64510 135280 64566 135289
rect 64510 135215 64566 135224
rect 64524 118590 64552 135215
rect 64616 133890 64644 160074
rect 64708 136921 64736 251262
rect 64800 137290 64828 283319
rect 65720 275330 65748 432482
rect 66180 432451 66208 432482
rect 66810 430400 66866 430409
rect 66810 430335 66866 430344
rect 66824 429214 66852 430335
rect 67284 429418 67312 433774
rect 67376 431497 67404 438126
rect 67362 431488 67418 431497
rect 67362 431423 67418 431432
rect 67376 431254 67404 431423
rect 67364 431248 67416 431254
rect 67364 431190 67416 431196
rect 67362 429448 67418 429457
rect 67272 429412 67324 429418
rect 67362 429383 67418 429392
rect 67272 429354 67324 429360
rect 67284 429321 67312 429354
rect 67270 429312 67326 429321
rect 67270 429247 67326 429256
rect 66812 429208 66864 429214
rect 66812 429150 66864 429156
rect 65800 427372 65852 427378
rect 65800 427314 65852 427320
rect 65708 275324 65760 275330
rect 65708 275266 65760 275272
rect 65812 271182 65840 427314
rect 67376 426329 67404 429383
rect 67362 426320 67418 426329
rect 67362 426255 67418 426264
rect 66996 425740 67048 425746
rect 66996 425682 67048 425688
rect 67008 425241 67036 425682
rect 67376 425649 67404 426255
rect 67362 425640 67418 425649
rect 67362 425575 67418 425584
rect 66994 425232 67050 425241
rect 66994 425167 67050 425176
rect 66718 424144 66774 424153
rect 66718 424079 66774 424088
rect 66732 423706 66760 424079
rect 66720 423700 66772 423706
rect 66720 423642 66772 423648
rect 66812 423632 66864 423638
rect 66812 423574 66864 423580
rect 66824 423337 66852 423574
rect 66810 423328 66866 423337
rect 66810 423263 66866 423272
rect 66810 421152 66866 421161
rect 66810 421087 66866 421096
rect 65984 421048 66036 421054
rect 65984 420990 66036 420996
rect 65892 294636 65944 294642
rect 65892 294578 65944 294584
rect 65904 279721 65932 294578
rect 65890 279712 65946 279721
rect 65890 279647 65946 279656
rect 65800 271176 65852 271182
rect 65800 271118 65852 271124
rect 65890 268560 65946 268569
rect 65890 268495 65946 268504
rect 65904 240825 65932 268495
rect 65996 267102 66024 420990
rect 66824 420986 66852 421087
rect 66812 420980 66864 420986
rect 66812 420922 66864 420928
rect 66904 420912 66956 420918
rect 66904 420854 66956 420860
rect 66812 420232 66864 420238
rect 66812 420174 66864 420180
rect 66442 418976 66498 418985
rect 66442 418911 66498 418920
rect 66456 418334 66484 418911
rect 66444 418328 66496 418334
rect 66444 418270 66496 418276
rect 66442 418160 66498 418169
rect 66442 418095 66444 418104
rect 66496 418095 66498 418104
rect 66444 418066 66496 418072
rect 66824 417081 66852 420174
rect 66916 420073 66944 420854
rect 66902 420064 66958 420073
rect 66902 419999 66958 420008
rect 66810 417072 66866 417081
rect 66810 417007 66866 417016
rect 66902 415984 66958 415993
rect 66902 415919 66958 415928
rect 66916 415478 66944 415919
rect 66904 415472 66956 415478
rect 66904 415414 66956 415420
rect 66810 414896 66866 414905
rect 66810 414831 66866 414840
rect 66824 414050 66852 414831
rect 67362 414080 67418 414089
rect 66812 414044 66864 414050
rect 67362 414015 67418 414024
rect 66812 413986 66864 413992
rect 66628 413296 66680 413302
rect 66628 413238 66680 413244
rect 66640 413001 66668 413238
rect 66626 412992 66682 413001
rect 66626 412927 66682 412936
rect 66902 411904 66958 411913
rect 66902 411839 66958 411848
rect 66916 411330 66944 411839
rect 66904 411324 66956 411330
rect 66904 411266 66956 411272
rect 66810 410816 66866 410825
rect 66810 410751 66866 410760
rect 66824 410582 66852 410751
rect 66812 410576 66864 410582
rect 66812 410518 66864 410524
rect 66442 408912 66498 408921
rect 66442 408847 66498 408856
rect 66456 408542 66484 408847
rect 66444 408536 66496 408542
rect 66444 408478 66496 408484
rect 66810 407824 66866 407833
rect 66810 407759 66812 407768
rect 66864 407759 66866 407768
rect 66812 407730 66864 407736
rect 66442 406736 66498 406745
rect 66442 406671 66498 406680
rect 66456 406434 66484 406671
rect 66444 406428 66496 406434
rect 66444 406370 66496 406376
rect 66902 404560 66958 404569
rect 66902 404495 66958 404504
rect 66916 404394 66944 404495
rect 66904 404388 66956 404394
rect 66904 404330 66956 404336
rect 66442 403744 66498 403753
rect 66442 403679 66498 403688
rect 66456 403034 66484 403679
rect 66444 403028 66496 403034
rect 66444 402970 66496 402976
rect 66442 401568 66498 401577
rect 66442 401503 66498 401512
rect 66456 400246 66484 401503
rect 67270 400480 67326 400489
rect 67270 400415 67326 400424
rect 66444 400240 66496 400246
rect 66444 400182 66496 400188
rect 66810 399664 66866 399673
rect 66810 399599 66866 399608
rect 66824 398886 66852 399599
rect 66812 398880 66864 398886
rect 66812 398822 66864 398828
rect 67088 398812 67140 398818
rect 67088 398754 67140 398760
rect 67100 398585 67128 398754
rect 67086 398576 67142 398585
rect 67086 398511 67142 398520
rect 66812 397520 66864 397526
rect 66810 397488 66812 397497
rect 66864 397488 66866 397497
rect 66810 397423 66866 397432
rect 66258 396400 66314 396409
rect 66258 396335 66314 396344
rect 66272 396098 66300 396335
rect 66260 396092 66312 396098
rect 66260 396034 66312 396040
rect 66626 392320 66682 392329
rect 66626 392255 66682 392264
rect 66640 392018 66668 392255
rect 66628 392012 66680 392018
rect 66628 391954 66680 391960
rect 67284 379506 67312 400415
rect 67376 382226 67404 414015
rect 67468 405657 67496 441586
rect 68192 434036 68244 434042
rect 68192 433978 68244 433984
rect 67732 433288 67784 433294
rect 67732 433230 67784 433236
rect 67548 433220 67600 433226
rect 67548 433162 67600 433168
rect 67560 428233 67588 433162
rect 67546 428224 67602 428233
rect 67546 428159 67602 428168
rect 67546 427408 67602 427417
rect 67546 427343 67548 427352
rect 67600 427343 67602 427352
rect 67548 427314 67600 427320
rect 67548 426420 67600 426426
rect 67548 426362 67600 426368
rect 67560 422249 67588 426362
rect 67546 422240 67602 422249
rect 67546 422175 67602 422184
rect 67560 421054 67588 422175
rect 67548 421048 67600 421054
rect 67548 420990 67600 420996
rect 67546 418160 67602 418169
rect 67546 418095 67602 418104
rect 67454 405648 67510 405657
rect 67454 405583 67510 405592
rect 67454 398576 67510 398585
rect 67454 398511 67510 398520
rect 67364 382220 67416 382226
rect 67364 382162 67416 382168
rect 67272 379500 67324 379506
rect 67272 379442 67324 379448
rect 67468 365673 67496 398511
rect 67454 365664 67510 365673
rect 67454 365599 67510 365608
rect 67560 339522 67588 418095
rect 67744 412634 67772 433230
rect 68204 426426 68232 433978
rect 68296 433226 68324 441594
rect 69676 441586 69888 441614
rect 69756 440904 69808 440910
rect 69756 440846 69808 440852
rect 68926 438152 68982 438161
rect 68926 438087 68982 438096
rect 68940 436286 68968 438087
rect 68928 436280 68980 436286
rect 68928 436222 68980 436228
rect 68652 436144 68704 436150
rect 68652 436086 68704 436092
rect 68284 433220 68336 433226
rect 68284 433162 68336 433168
rect 68192 426420 68244 426426
rect 68192 426362 68244 426368
rect 67652 412606 67772 412634
rect 67652 409737 67680 412606
rect 67638 409728 67694 409737
rect 67638 409663 67694 409672
rect 67640 402960 67692 402966
rect 67640 402902 67692 402908
rect 67652 402665 67680 402902
rect 67638 402656 67694 402665
rect 67638 402591 67694 402600
rect 67652 376553 67680 402591
rect 67744 393417 67772 393443
rect 67730 393408 67786 393417
rect 67730 393343 67732 393352
rect 67784 393343 67786 393352
rect 67732 393314 67784 393320
rect 67638 376544 67694 376553
rect 67638 376479 67694 376488
rect 67744 367062 67772 393314
rect 68560 391944 68612 391950
rect 68560 391886 68612 391892
rect 68572 391241 68600 391886
rect 68558 391232 68614 391241
rect 68558 391167 68614 391176
rect 68664 390538 68692 436086
rect 68940 434330 68968 436222
rect 68816 434302 68968 434330
rect 69202 434344 69258 434353
rect 69768 434330 69796 440846
rect 69860 434761 69888 441586
rect 70490 436248 70546 436257
rect 70490 436183 70492 436192
rect 70544 436183 70546 436192
rect 70858 436248 70914 436257
rect 70858 436183 70914 436192
rect 70492 436154 70544 436160
rect 69846 434752 69902 434761
rect 69846 434687 69902 434696
rect 69258 434302 69796 434330
rect 69860 434330 69888 434687
rect 69860 434302 70288 434330
rect 69202 434279 69258 434288
rect 70872 434058 70900 436183
rect 70872 434030 71024 434058
rect 71148 433838 71176 442954
rect 71792 436218 71820 539786
rect 73172 539730 73200 539854
rect 94318 539815 94374 539824
rect 89718 539744 89774 539753
rect 73172 539716 73416 539730
rect 73172 539702 73430 539716
rect 71884 539158 72496 539186
rect 71884 529310 71912 539158
rect 73402 539050 73430 539702
rect 89718 539679 89774 539688
rect 89732 539594 89760 539679
rect 89240 539566 89760 539594
rect 91744 539640 91796 539646
rect 91744 539582 91796 539588
rect 73632 539158 74336 539186
rect 74552 539158 75256 539186
rect 76024 539158 76176 539186
rect 76760 539158 77096 539186
rect 77312 539158 78016 539186
rect 78936 539158 79272 539186
rect 80040 539158 80192 539186
rect 73402 539022 73476 539050
rect 73160 537532 73212 537538
rect 73160 537474 73212 537480
rect 73172 536790 73200 537474
rect 73160 536784 73212 536790
rect 73160 536726 73212 536732
rect 72424 536580 72476 536586
rect 72424 536522 72476 536528
rect 71872 529304 71924 529310
rect 71872 529246 71924 529252
rect 72436 518226 72464 536522
rect 73448 532030 73476 539022
rect 73436 532024 73488 532030
rect 73436 531966 73488 531972
rect 73632 528554 73660 539158
rect 73172 528526 73660 528554
rect 72424 518220 72476 518226
rect 72424 518162 72476 518168
rect 73172 455394 73200 528526
rect 73160 455388 73212 455394
rect 73160 455330 73212 455336
rect 74552 454714 74580 539158
rect 75828 532092 75880 532098
rect 75828 532034 75880 532040
rect 75840 458250 75868 532034
rect 76024 509250 76052 539158
rect 76760 536790 76788 539158
rect 76748 536784 76800 536790
rect 76748 536726 76800 536732
rect 76012 509244 76064 509250
rect 76012 509186 76064 509192
rect 76024 508366 76052 509186
rect 76012 508360 76064 508366
rect 76012 508302 76064 508308
rect 76564 508360 76616 508366
rect 76564 508302 76616 508308
rect 75184 458244 75236 458250
rect 75184 458186 75236 458192
rect 75828 458244 75880 458250
rect 75828 458186 75880 458192
rect 74540 454708 74592 454714
rect 74540 454650 74592 454656
rect 74446 452704 74502 452713
rect 74446 452639 74502 452648
rect 72424 444440 72476 444446
rect 72424 444382 72476 444388
rect 71780 436212 71832 436218
rect 71780 436154 71832 436160
rect 72436 436150 72464 444382
rect 73896 438252 73948 438258
rect 73896 438194 73948 438200
rect 72700 436212 72752 436218
rect 72700 436154 72752 436160
rect 71688 436144 71740 436150
rect 71688 436086 71740 436092
rect 72424 436144 72476 436150
rect 72424 436086 72476 436092
rect 71700 434330 71728 436086
rect 72606 434888 72662 434897
rect 72606 434823 72662 434832
rect 72620 434330 72648 434823
rect 71576 434302 71728 434330
rect 72312 434302 72648 434330
rect 72712 434330 72740 436154
rect 73908 434330 73936 438194
rect 72712 434302 73048 434330
rect 73784 434302 73936 434330
rect 71136 433832 71188 433838
rect 71136 433774 71188 433780
rect 70676 433696 70728 433702
rect 70674 433664 70676 433673
rect 70728 433664 70730 433673
rect 70674 433599 70730 433608
rect 74078 433664 74134 433673
rect 74460 433650 74488 452639
rect 75196 436257 75224 458186
rect 75828 451920 75880 451926
rect 75828 451862 75880 451868
rect 75840 441614 75868 451862
rect 76576 443057 76604 508302
rect 77312 464370 77340 539158
rect 79244 538218 79272 539158
rect 80164 538393 80192 539158
rect 80256 539158 80960 539186
rect 81880 539158 82216 539186
rect 82800 539158 82860 539186
rect 83720 539158 84056 539186
rect 80150 538384 80206 538393
rect 80150 538319 80206 538328
rect 79232 538212 79284 538218
rect 79232 538154 79284 538160
rect 79244 537062 79272 538154
rect 79232 537056 79284 537062
rect 79232 536998 79284 537004
rect 79968 537056 80020 537062
rect 79968 536998 80020 537004
rect 79980 471306 80008 536998
rect 80256 528554 80284 539158
rect 82188 536722 82216 539158
rect 82176 536716 82228 536722
rect 82176 536658 82228 536664
rect 82728 533384 82780 533390
rect 82728 533326 82780 533332
rect 80072 528526 80284 528554
rect 79968 471300 80020 471306
rect 79968 471242 80020 471248
rect 79324 468512 79376 468518
rect 79324 468454 79376 468460
rect 77300 464364 77352 464370
rect 77300 464306 77352 464312
rect 77944 452668 77996 452674
rect 77944 452610 77996 452616
rect 76656 446412 76708 446418
rect 76656 446354 76708 446360
rect 76562 443048 76618 443057
rect 76562 442983 76618 442992
rect 75472 441586 75868 441614
rect 75472 437474 75500 441586
rect 75380 437446 75500 437474
rect 75182 436248 75238 436257
rect 75182 436183 75238 436192
rect 74134 433622 74488 433650
rect 74814 433664 74870 433673
rect 74078 433599 74134 433608
rect 75380 433650 75408 437446
rect 76576 437442 76604 442983
rect 76668 438190 76696 446354
rect 76840 439612 76892 439618
rect 76840 439554 76892 439560
rect 76656 438184 76708 438190
rect 76656 438126 76708 438132
rect 76564 437436 76616 437442
rect 76564 437378 76616 437384
rect 75458 433800 75514 433809
rect 75514 433758 75808 433786
rect 75458 433735 75514 433744
rect 74870 433622 75408 433650
rect 76194 433664 76250 433673
rect 74814 433599 74870 433608
rect 76852 433650 76880 439554
rect 77956 438258 77984 452610
rect 78680 449948 78732 449954
rect 78680 449890 78732 449896
rect 78692 441614 78720 449890
rect 78692 441586 78904 441614
rect 77944 438252 77996 438258
rect 77944 438194 77996 438200
rect 77390 437608 77446 437617
rect 77390 437543 77446 437552
rect 77404 434330 77432 437543
rect 78588 437504 78640 437510
rect 78588 437446 78640 437452
rect 78600 434602 78628 437446
rect 77280 434302 77432 434330
rect 78554 434574 78628 434602
rect 78554 434316 78582 434574
rect 78876 434330 78904 441586
rect 79336 437617 79364 468454
rect 80072 458833 80100 528526
rect 81346 525872 81402 525881
rect 81346 525807 81402 525816
rect 80058 458824 80114 458833
rect 80058 458759 80114 458768
rect 81360 457473 81388 525807
rect 81346 457464 81402 457473
rect 81346 457399 81402 457408
rect 82740 455462 82768 533326
rect 82832 462330 82860 539158
rect 84028 538121 84056 539158
rect 84304 539158 84640 539186
rect 85560 539158 85896 539186
rect 86480 539158 86724 539186
rect 87400 539158 87736 539186
rect 88320 539158 88380 539186
rect 84014 538112 84070 538121
rect 84014 538047 84070 538056
rect 84304 533361 84332 539158
rect 85868 538286 85896 539158
rect 85856 538280 85908 538286
rect 85856 538222 85908 538228
rect 86224 536104 86276 536110
rect 86224 536046 86276 536052
rect 84290 533352 84346 533361
rect 84290 533287 84346 533296
rect 85488 476808 85540 476814
rect 85488 476750 85540 476756
rect 82820 462324 82872 462330
rect 82820 462266 82872 462272
rect 83464 461644 83516 461650
rect 83464 461586 83516 461592
rect 82084 455456 82136 455462
rect 82084 455398 82136 455404
rect 82728 455456 82780 455462
rect 82728 455398 82780 455404
rect 80060 443692 80112 443698
rect 80060 443634 80112 443640
rect 79322 437608 79378 437617
rect 79322 437543 79378 437552
rect 80072 436257 80100 443634
rect 81440 438184 81492 438190
rect 81440 438126 81492 438132
rect 80242 436384 80298 436393
rect 80242 436319 80298 436328
rect 80058 436248 80114 436257
rect 80058 436183 80114 436192
rect 80072 434602 80100 436183
rect 80026 434574 80100 434602
rect 78876 434302 79304 434330
rect 80026 434316 80054 434574
rect 80256 434330 80284 436319
rect 81452 436098 81480 438126
rect 82096 436121 82124 455398
rect 83476 444514 83504 461586
rect 83464 444508 83516 444514
rect 83464 444450 83516 444456
rect 82912 437436 82964 437442
rect 82912 437378 82964 437384
rect 81360 436070 81480 436098
rect 82082 436112 82138 436121
rect 81360 434602 81388 436070
rect 82082 436047 82138 436056
rect 82096 434602 82124 436047
rect 81314 434574 81388 434602
rect 82050 434574 82124 434602
rect 80978 434344 81034 434353
rect 80256 434302 80592 434330
rect 81314 434330 81342 434574
rect 81034 434316 81342 434330
rect 82050 434316 82078 434574
rect 81034 434302 81328 434316
rect 80978 434279 81034 434288
rect 82924 434194 82952 437378
rect 83476 434602 83504 444450
rect 85500 441614 85528 476750
rect 86236 460222 86264 536046
rect 86696 535974 86724 539158
rect 87708 536761 87736 539158
rect 88248 536852 88300 536858
rect 88248 536794 88300 536800
rect 87694 536752 87750 536761
rect 87694 536687 87750 536696
rect 86684 535968 86736 535974
rect 86684 535910 86736 535916
rect 87604 535968 87656 535974
rect 87604 535910 87656 535916
rect 87616 463010 87644 535910
rect 87604 463004 87656 463010
rect 87604 462946 87656 462952
rect 85672 460216 85724 460222
rect 85672 460158 85724 460164
rect 86224 460216 86276 460222
rect 86224 460158 86276 460164
rect 85224 441586 85528 441614
rect 85684 441614 85712 460158
rect 88260 444378 88288 536794
rect 88352 530777 88380 539158
rect 89732 539158 90160 539186
rect 91204 539158 91264 539186
rect 88338 530768 88394 530777
rect 88338 530703 88394 530712
rect 88982 484392 89038 484401
rect 88982 484327 89038 484336
rect 88996 483041 89024 484327
rect 88982 483032 89038 483041
rect 88982 482967 89038 482976
rect 86960 444372 87012 444378
rect 86960 444314 87012 444320
rect 88248 444372 88300 444378
rect 88248 444314 88300 444320
rect 85684 441586 85896 441614
rect 83740 439544 83792 439550
rect 83740 439486 83792 439492
rect 83476 434574 83550 434602
rect 83522 434316 83550 434574
rect 83752 434489 83780 439486
rect 83738 434480 83794 434489
rect 83738 434415 83794 434424
rect 83752 434330 83780 434415
rect 84566 434344 84622 434353
rect 83752 434302 84088 434330
rect 85224 434330 85252 441586
rect 85868 434353 85896 441586
rect 86972 434602 87000 444314
rect 88260 443766 88288 444314
rect 88248 443760 88300 443766
rect 88248 443702 88300 443708
rect 88996 438190 89024 482967
rect 89732 439618 89760 539158
rect 91008 535492 91060 535498
rect 91008 535434 91060 535440
rect 91020 469305 91048 535434
rect 90362 469296 90418 469305
rect 90362 469231 90418 469240
rect 91006 469296 91062 469305
rect 91006 469231 91062 469240
rect 89720 439612 89772 439618
rect 89720 439554 89772 439560
rect 88984 438184 89036 438190
rect 90376 438161 90404 469231
rect 91204 468518 91232 539158
rect 91756 536722 91784 539582
rect 91848 539158 92184 539186
rect 93104 539158 93440 539186
rect 94024 539158 94084 539186
rect 91744 536716 91796 536722
rect 91744 536658 91796 536664
rect 91848 535498 91876 539158
rect 93412 536790 93440 539158
rect 93400 536784 93452 536790
rect 93400 536726 93452 536732
rect 91836 535492 91888 535498
rect 91836 535434 91888 535440
rect 94056 531214 94084 539158
rect 93124 531208 93176 531214
rect 93124 531150 93176 531156
rect 94044 531208 94096 531214
rect 94044 531150 94096 531156
rect 93136 522306 93164 531150
rect 94332 528554 94360 539815
rect 94594 538928 94650 538937
rect 94594 538863 94650 538872
rect 94608 538354 94636 538863
rect 94596 538348 94648 538354
rect 94596 538290 94648 538296
rect 94700 533390 94728 558583
rect 94778 555520 94834 555529
rect 94778 555455 94834 555464
rect 94688 533384 94740 533390
rect 94688 533326 94740 533332
rect 94148 528526 94360 528554
rect 93124 522300 93176 522306
rect 93124 522242 93176 522248
rect 92572 515432 92624 515438
rect 92572 515374 92624 515380
rect 91192 468512 91244 468518
rect 91192 468454 91244 468460
rect 90640 438184 90692 438190
rect 88984 438126 89036 438132
rect 90362 438152 90418 438161
rect 90640 438126 90692 438132
rect 90362 438087 90418 438096
rect 89350 436792 89406 436801
rect 89350 436727 89406 436736
rect 86972 434574 87046 434602
rect 84622 434302 85252 434330
rect 85854 434344 85910 434353
rect 84566 434279 84622 434288
rect 85910 434302 86296 434330
rect 87018 434316 87046 434574
rect 89364 434330 89392 436727
rect 89056 434302 89392 434330
rect 85854 434279 85910 434288
rect 85868 434219 85896 434279
rect 82800 434166 82952 434194
rect 90652 433945 90680 438126
rect 91098 436112 91154 436121
rect 91098 436047 91154 436056
rect 91112 434602 91140 436047
rect 92584 434602 92612 515374
rect 94148 476814 94176 528526
rect 94792 523705 94820 555455
rect 94778 523696 94834 523705
rect 94778 523631 94834 523640
rect 94504 522300 94556 522306
rect 94504 522242 94556 522248
rect 94136 476808 94188 476814
rect 94136 476750 94188 476756
rect 93952 472660 94004 472666
rect 93952 472602 94004 472608
rect 93860 468512 93912 468518
rect 93860 468454 93912 468460
rect 93872 434602 93900 468454
rect 93964 441614 93992 472602
rect 94516 465594 94544 522242
rect 95252 520985 95280 563615
rect 95344 558929 95372 588934
rect 95422 565856 95478 565865
rect 95422 565791 95478 565800
rect 95330 558920 95386 558929
rect 95330 558855 95386 558864
rect 95330 545728 95386 545737
rect 95330 545663 95386 545672
rect 95238 520976 95294 520985
rect 95238 520911 95294 520920
rect 94594 482216 94650 482225
rect 94594 482151 94650 482160
rect 94608 472666 94636 482151
rect 94596 472660 94648 472666
rect 94596 472602 94648 472608
rect 94504 465588 94556 465594
rect 94504 465530 94556 465536
rect 95148 465588 95200 465594
rect 95148 465530 95200 465536
rect 95160 465118 95188 465530
rect 95148 465112 95200 465118
rect 95148 465054 95200 465060
rect 95160 448594 95188 465054
rect 95240 449268 95292 449274
rect 95240 449210 95292 449216
rect 95148 448588 95200 448594
rect 95148 448530 95200 448536
rect 93964 441586 94176 441614
rect 91066 434574 91140 434602
rect 92538 434574 92612 434602
rect 93826 434574 93900 434602
rect 91066 434316 91094 434574
rect 92538 434194 92566 434574
rect 93826 434316 93854 434574
rect 94148 434330 94176 441586
rect 95252 434602 95280 449210
rect 95344 444961 95372 545663
rect 95436 536858 95464 565791
rect 96632 552129 96660 702510
rect 105464 700330 105492 703520
rect 137848 702642 137876 703520
rect 137836 702636 137888 702642
rect 137836 702578 137888 702584
rect 154132 702574 154160 703520
rect 170324 702778 170352 703520
rect 184296 703044 184348 703050
rect 184296 702986 184348 702992
rect 169760 702772 169812 702778
rect 169760 702714 169812 702720
rect 170312 702772 170364 702778
rect 170312 702714 170364 702720
rect 154120 702568 154172 702574
rect 154120 702510 154172 702516
rect 169772 702506 169800 702714
rect 169760 702500 169812 702506
rect 169760 702442 169812 702448
rect 180064 702500 180116 702506
rect 180064 702442 180116 702448
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 144828 622464 144880 622470
rect 144828 622406 144880 622412
rect 129648 618316 129700 618322
rect 129648 618258 129700 618264
rect 123484 610020 123536 610026
rect 123484 609962 123536 609968
rect 98644 605872 98696 605878
rect 98644 605814 98696 605820
rect 98656 583438 98684 605814
rect 115294 604480 115350 604489
rect 115294 604415 115350 604424
rect 104164 601724 104216 601730
rect 104164 601666 104216 601672
rect 98644 583432 98696 583438
rect 98644 583374 98696 583380
rect 98550 581224 98606 581233
rect 98550 581159 98606 581168
rect 96802 578912 96858 578921
rect 96802 578847 96858 578856
rect 96816 578270 96844 578847
rect 96804 578264 96856 578270
rect 96804 578206 96856 578212
rect 98564 578202 98592 581159
rect 98644 580712 98696 580718
rect 98644 580654 98696 580660
rect 98656 579698 98684 580654
rect 98644 579692 98696 579698
rect 98644 579634 98696 579640
rect 98552 578196 98604 578202
rect 98552 578138 98604 578144
rect 97906 577552 97962 577561
rect 97962 577510 98040 577538
rect 97906 577487 97962 577496
rect 97908 576836 97960 576842
rect 97908 576778 97960 576784
rect 97920 576745 97948 576778
rect 97906 576736 97962 576745
rect 97906 576671 97962 576680
rect 96712 576088 96764 576094
rect 96712 576030 96764 576036
rect 96724 569129 96752 576030
rect 96802 574832 96858 574841
rect 96802 574767 96858 574776
rect 96816 574122 96844 574767
rect 96804 574116 96856 574122
rect 96804 574058 96856 574064
rect 96894 573472 96950 573481
rect 96894 573407 96950 573416
rect 96908 572762 96936 573407
rect 98012 573374 98040 577510
rect 98000 573368 98052 573374
rect 98000 573310 98052 573316
rect 96896 572756 96948 572762
rect 96896 572698 96948 572704
rect 97908 572688 97960 572694
rect 97906 572656 97908 572665
rect 97960 572656 97962 572665
rect 97906 572591 97962 572600
rect 97722 571432 97778 571441
rect 97722 571367 97724 571376
rect 97776 571367 97778 571376
rect 97724 571338 97776 571344
rect 97906 570072 97962 570081
rect 97906 570007 97962 570016
rect 97920 569974 97948 570007
rect 97908 569968 97960 569974
rect 97908 569910 97960 569916
rect 97448 569220 97500 569226
rect 97448 569162 97500 569168
rect 97460 569129 97488 569162
rect 96710 569120 96766 569129
rect 96710 569055 96766 569064
rect 97446 569120 97502 569129
rect 97446 569055 97502 569064
rect 96804 568540 96856 568546
rect 96804 568482 96856 568488
rect 96816 567905 96844 568482
rect 96802 567896 96858 567905
rect 96802 567831 96858 567840
rect 96894 561096 96950 561105
rect 96894 561031 96950 561040
rect 96908 560998 96936 561031
rect 96896 560992 96948 560998
rect 96896 560934 96948 560940
rect 96710 556880 96766 556889
rect 96710 556815 96766 556824
rect 96618 552120 96674 552129
rect 96618 552055 96674 552064
rect 96436 538280 96488 538286
rect 96436 538222 96488 538228
rect 95424 536852 95476 536858
rect 95424 536794 95476 536800
rect 96448 533361 96476 538222
rect 96434 533352 96490 533361
rect 96434 533287 96490 533296
rect 96724 526454 96752 556815
rect 96908 547874 96936 560934
rect 96986 559600 97042 559609
rect 96986 559535 97042 559544
rect 97000 558958 97028 559535
rect 96988 558952 97040 558958
rect 96988 558894 97040 558900
rect 97906 556880 97962 556889
rect 97906 556815 97908 556824
rect 97960 556815 97962 556824
rect 97908 556786 97960 556792
rect 96986 554160 97042 554169
rect 96986 554095 97042 554104
rect 96816 547846 96936 547874
rect 96816 532098 96844 547846
rect 96894 541784 96950 541793
rect 96894 541719 96950 541728
rect 96908 534750 96936 541719
rect 96896 534744 96948 534750
rect 96896 534686 96948 534692
rect 96804 532092 96856 532098
rect 96804 532034 96856 532040
rect 96712 526448 96764 526454
rect 96712 526390 96764 526396
rect 95884 448588 95936 448594
rect 95884 448530 95936 448536
rect 95330 444952 95386 444961
rect 95330 444887 95386 444896
rect 95896 436354 95924 448530
rect 97000 441614 97028 554095
rect 97906 552800 97962 552809
rect 97906 552735 97962 552744
rect 97920 552362 97948 552735
rect 97908 552356 97960 552362
rect 97908 552298 97960 552304
rect 97906 552120 97962 552129
rect 97906 552055 97962 552064
rect 97920 549914 97948 552055
rect 97908 549908 97960 549914
rect 97908 549850 97960 549856
rect 97538 544368 97594 544377
rect 97538 544303 97594 544312
rect 97552 543794 97580 544303
rect 97540 543788 97592 543794
rect 97540 543730 97592 543736
rect 97538 543008 97594 543017
rect 97538 542943 97594 542952
rect 97552 542434 97580 542943
rect 97540 542428 97592 542434
rect 97540 542370 97592 542376
rect 97906 541784 97962 541793
rect 97906 541719 97962 541728
rect 97920 541686 97948 541719
rect 97908 541680 97960 541686
rect 97908 541622 97960 541628
rect 98012 528562 98040 573310
rect 101404 571396 101456 571402
rect 101404 571338 101456 571344
rect 98090 562320 98146 562329
rect 98090 562255 98146 562264
rect 98104 559570 98132 562255
rect 98092 559564 98144 559570
rect 98092 559506 98144 559512
rect 100760 552356 100812 552362
rect 100760 552298 100812 552304
rect 100772 548554 100800 552298
rect 101416 551993 101444 571338
rect 101402 551984 101458 551993
rect 101402 551919 101458 551928
rect 100760 548548 100812 548554
rect 100760 548490 100812 548496
rect 99380 546508 99432 546514
rect 99380 546450 99432 546456
rect 99392 538286 99420 546450
rect 104176 538354 104204 601666
rect 112444 597644 112496 597650
rect 112444 597586 112496 597592
rect 106924 585812 106976 585818
rect 106924 585754 106976 585760
rect 105542 581088 105598 581097
rect 105542 581023 105598 581032
rect 105556 551342 105584 581023
rect 105544 551336 105596 551342
rect 105544 551278 105596 551284
rect 104256 543788 104308 543794
rect 104256 543730 104308 543736
rect 104164 538348 104216 538354
rect 104164 538290 104216 538296
rect 99380 538280 99432 538286
rect 99380 538222 99432 538228
rect 102784 532024 102836 532030
rect 102784 531966 102836 531972
rect 98000 528556 98052 528562
rect 98000 528498 98052 528504
rect 99472 518220 99524 518226
rect 99472 518162 99524 518168
rect 98000 492720 98052 492726
rect 98000 492662 98052 492668
rect 96908 441586 97028 441614
rect 95884 436348 95936 436354
rect 95884 436290 95936 436296
rect 96344 436144 96396 436150
rect 96908 436121 96936 441586
rect 96988 436348 97040 436354
rect 96988 436290 97040 436296
rect 96344 436086 96396 436092
rect 96894 436112 96950 436121
rect 95252 434574 95326 434602
rect 94148 434302 94576 434330
rect 95298 434316 95326 434574
rect 95698 434344 95754 434353
rect 96356 434330 96384 436086
rect 96894 436047 96950 436056
rect 96908 434330 96936 436047
rect 95754 434302 96384 434330
rect 96600 434302 96936 434330
rect 97000 434330 97028 436290
rect 98012 434602 98040 492662
rect 98734 462360 98790 462369
rect 98734 462295 98790 462304
rect 98748 451926 98776 462295
rect 98736 451920 98788 451926
rect 98642 451888 98698 451897
rect 98736 451862 98788 451868
rect 98642 451823 98698 451832
rect 98656 436801 98684 451823
rect 99484 441614 99512 518162
rect 102796 471986 102824 531966
rect 104268 528562 104296 543730
rect 106936 535430 106964 585754
rect 111064 583840 111116 583846
rect 111064 583782 111116 583788
rect 108304 578944 108356 578950
rect 108304 578886 108356 578892
rect 106924 535424 106976 535430
rect 106924 535366 106976 535372
rect 104256 528556 104308 528562
rect 104256 528498 104308 528504
rect 104808 528556 104860 528562
rect 104808 528498 104860 528504
rect 102140 471980 102192 471986
rect 102140 471922 102192 471928
rect 102784 471980 102836 471986
rect 102784 471922 102836 471928
rect 101404 471300 101456 471306
rect 101404 471242 101456 471248
rect 100024 457496 100076 457502
rect 100024 457438 100076 457444
rect 99484 441586 99696 441614
rect 98642 436792 98698 436801
rect 98642 436727 98698 436736
rect 98012 434574 98086 434602
rect 97000 434302 97336 434330
rect 98058 434316 98086 434574
rect 99668 434330 99696 441586
rect 100036 436150 100064 457438
rect 101416 437442 101444 471242
rect 102152 470626 102180 471922
rect 102140 470620 102192 470626
rect 102140 470562 102192 470568
rect 102152 441614 102180 470562
rect 104820 460970 104848 528498
rect 108316 495514 108344 578886
rect 108948 496120 109000 496126
rect 108948 496062 109000 496068
rect 108960 495514 108988 496062
rect 108304 495508 108356 495514
rect 108304 495450 108356 495456
rect 108948 495508 109000 495514
rect 108948 495450 109000 495456
rect 108856 473408 108908 473414
rect 108856 473350 108908 473356
rect 106280 463752 106332 463758
rect 106280 463694 106332 463700
rect 104900 463004 104952 463010
rect 104900 462946 104952 462952
rect 104912 462398 104940 462946
rect 104900 462392 104952 462398
rect 104900 462334 104952 462340
rect 104808 460964 104860 460970
rect 104808 460906 104860 460912
rect 104164 450560 104216 450566
rect 104164 450502 104216 450508
rect 102152 441586 102640 441614
rect 101404 437436 101456 437442
rect 101404 437378 101456 437384
rect 102508 437368 102560 437374
rect 102508 437310 102560 437316
rect 100024 436144 100076 436150
rect 100024 436086 100076 436092
rect 100206 434344 100262 434353
rect 99668 434302 100206 434330
rect 95698 434279 95754 434288
rect 102520 434330 102548 437310
rect 102304 434302 102548 434330
rect 102612 434330 102640 441586
rect 104176 441522 104204 450502
rect 104164 441516 104216 441522
rect 104164 441458 104216 441464
rect 104176 438954 104204 441458
rect 104176 438926 104296 438954
rect 104820 438938 104848 460906
rect 104912 441614 104940 462334
rect 105544 451920 105596 451926
rect 105544 451862 105596 451868
rect 104912 441586 105400 441614
rect 104164 437436 104216 437442
rect 104164 437378 104216 437384
rect 104176 436150 104204 437378
rect 103888 436144 103940 436150
rect 103888 436086 103940 436092
rect 104164 436144 104216 436150
rect 104164 436086 104216 436092
rect 103900 434330 103928 436086
rect 104268 434602 104296 438926
rect 104808 438932 104860 438938
rect 104808 438874 104860 438880
rect 104268 434574 104342 434602
rect 102612 434302 103040 434330
rect 103592 434302 103928 434330
rect 104314 434316 104342 434574
rect 105372 434330 105400 441586
rect 105556 437374 105584 451862
rect 105544 437368 105596 437374
rect 105544 437310 105596 437316
rect 106292 434602 106320 463694
rect 108868 462330 108896 473350
rect 108856 462324 108908 462330
rect 108856 462266 108908 462272
rect 107660 438932 107712 438938
rect 107660 438874 107712 438880
rect 107672 436257 107700 438874
rect 108960 436257 108988 495450
rect 111076 478174 111104 583782
rect 111800 572756 111852 572762
rect 111800 572698 111852 572704
rect 111812 572014 111840 572698
rect 112456 572694 112484 597586
rect 112444 572688 112496 572694
rect 112444 572630 112496 572636
rect 111800 572008 111852 572014
rect 111800 571950 111852 571956
rect 115204 559564 115256 559570
rect 115204 559506 115256 559512
rect 113824 558952 113876 558958
rect 113824 558894 113876 558900
rect 112444 548548 112496 548554
rect 112444 548490 112496 548496
rect 112456 532710 112484 548490
rect 112444 532704 112496 532710
rect 112444 532646 112496 532652
rect 113088 532704 113140 532710
rect 113088 532646 113140 532652
rect 111064 478168 111116 478174
rect 111064 478110 111116 478116
rect 111076 477562 111104 478110
rect 110420 477556 110472 477562
rect 110420 477498 110472 477504
rect 111064 477556 111116 477562
rect 111064 477498 111116 477504
rect 109040 462324 109092 462330
rect 109040 462266 109092 462272
rect 109052 441614 109080 462266
rect 110432 441614 110460 477498
rect 110512 464364 110564 464370
rect 110512 464306 110564 464312
rect 110524 461650 110552 464306
rect 110512 461644 110564 461650
rect 110512 461586 110564 461592
rect 113100 459610 113128 532646
rect 112444 459604 112496 459610
rect 112444 459546 112496 459552
rect 113088 459604 113140 459610
rect 113088 459546 113140 459552
rect 109052 441586 109448 441614
rect 110432 441586 110920 441614
rect 107658 436248 107714 436257
rect 107658 436183 107714 436192
rect 108946 436248 109002 436257
rect 108946 436183 109002 436192
rect 106292 434574 106366 434602
rect 105372 434302 105800 434330
rect 106338 434316 106366 434574
rect 107672 434330 107700 436183
rect 108960 434330 108988 436183
rect 107672 434302 107824 434330
rect 108560 434302 108988 434330
rect 109420 434330 109448 441586
rect 110788 436756 110840 436762
rect 110788 436698 110840 436704
rect 110800 434330 110828 436698
rect 109420 434302 109848 434330
rect 110584 434302 110828 434330
rect 110892 434330 110920 441586
rect 112260 434852 112312 434858
rect 112260 434794 112312 434800
rect 112272 434330 112300 434794
rect 112456 434330 112484 459546
rect 112996 455388 113048 455394
rect 112996 455330 113048 455336
rect 113008 454073 113036 455330
rect 112994 454064 113050 454073
rect 112994 453999 113050 454008
rect 113836 450702 113864 558894
rect 115216 558890 115244 559506
rect 115204 558884 115256 558890
rect 115204 558826 115256 558832
rect 114560 460216 114612 460222
rect 114560 460158 114612 460164
rect 113824 450696 113876 450702
rect 113824 450638 113876 450644
rect 114468 450696 114520 450702
rect 114468 450638 114520 450644
rect 114480 450022 114508 450638
rect 114468 450016 114520 450022
rect 114468 449958 114520 449964
rect 110892 434302 111320 434330
rect 112272 434302 112608 434330
rect 100206 434279 100262 434288
rect 92662 434208 92718 434217
rect 92538 434180 92662 434194
rect 92552 434166 92662 434180
rect 92662 434143 92718 434152
rect 90638 433936 90694 433945
rect 90638 433871 90694 433880
rect 101218 433800 101274 433809
rect 101274 433758 101568 433786
rect 101218 433735 101274 433744
rect 78126 433664 78182 433673
rect 76250 433622 76880 433650
rect 77832 433622 78126 433650
rect 76194 433599 76250 433608
rect 85854 433664 85910 433673
rect 85560 433622 85854 433650
rect 78126 433599 78182 433608
rect 85854 433599 85910 433608
rect 87326 433664 87382 433673
rect 87970 433664 88026 433673
rect 87382 433622 87584 433650
rect 87326 433599 87382 433608
rect 89626 433664 89682 433673
rect 88026 433622 88320 433650
rect 87970 433599 88026 433608
rect 90086 433664 90142 433673
rect 89682 433622 89792 433650
rect 89626 433599 89682 433608
rect 91558 433664 91614 433673
rect 90142 433622 90344 433650
rect 90086 433599 90142 433608
rect 92938 433664 92994 433673
rect 91614 433622 91816 433650
rect 91558 433599 91614 433608
rect 98458 433664 98514 433673
rect 92994 433622 93288 433650
rect 92938 433599 92994 433608
rect 99838 433664 99894 433673
rect 98514 433622 98808 433650
rect 99544 433622 99838 433650
rect 98458 433599 98514 433608
rect 100942 433664 100998 433673
rect 100832 433622 100942 433650
rect 99838 433599 99894 433608
rect 105174 433664 105230 433673
rect 105064 433622 105174 433650
rect 100942 433599 100998 433608
rect 105174 433599 105230 433608
rect 106738 433664 106794 433673
rect 109498 433664 109554 433673
rect 106794 433622 107088 433650
rect 109296 433622 109498 433650
rect 106738 433599 106794 433608
rect 109498 433599 109554 433608
rect 111706 433664 111762 433673
rect 111762 433622 112056 433650
rect 111706 433599 111762 433608
rect 113270 428224 113326 428233
rect 113270 428159 113326 428168
rect 113178 420880 113234 420889
rect 113178 420815 113234 420824
rect 113086 407144 113142 407153
rect 113086 407079 113088 407088
rect 113140 407079 113142 407088
rect 113088 407050 113140 407056
rect 93952 390992 94004 390998
rect 82174 390960 82230 390969
rect 81880 390918 82174 390946
rect 82174 390895 82230 390904
rect 85486 390960 85542 390969
rect 93840 390940 93952 390946
rect 93840 390934 94004 390940
rect 99470 390960 99526 390969
rect 93840 390918 93992 390934
rect 85486 390895 85542 390904
rect 83186 390688 83242 390697
rect 83242 390646 83352 390674
rect 83186 390623 83242 390632
rect 68572 390510 68692 390538
rect 79120 390510 79456 390538
rect 67824 390176 67876 390182
rect 67824 390118 67876 390124
rect 67836 371210 67864 390118
rect 68572 383654 68600 390510
rect 72422 390416 72478 390425
rect 68802 390182 68830 390388
rect 69124 390374 69368 390402
rect 69768 390374 70104 390402
rect 70504 390374 70840 390402
rect 71240 390374 71576 390402
rect 72128 390374 72422 390402
rect 68790 390176 68842 390182
rect 68790 390118 68842 390124
rect 69020 387048 69072 387054
rect 69020 386990 69072 386996
rect 68572 383626 68692 383654
rect 67824 371204 67876 371210
rect 67824 371146 67876 371152
rect 67732 367056 67784 367062
rect 67732 366998 67784 367004
rect 67836 354674 67864 371146
rect 67652 354646 67864 354674
rect 67548 339516 67600 339522
rect 67548 339458 67600 339464
rect 67560 335354 67588 339458
rect 67468 335326 67588 335354
rect 67362 325000 67418 325009
rect 67362 324935 67418 324944
rect 67272 295996 67324 296002
rect 67272 295938 67324 295944
rect 67284 282169 67312 295938
rect 67270 282160 67326 282169
rect 67270 282095 67326 282104
rect 67270 281344 67326 281353
rect 67270 281279 67326 281288
rect 67284 280226 67312 281279
rect 67272 280220 67324 280226
rect 67272 280162 67324 280168
rect 66810 278896 66866 278905
rect 66810 278831 66866 278840
rect 66824 278798 66852 278831
rect 66812 278792 66864 278798
rect 66812 278734 66864 278740
rect 67284 277982 67312 280162
rect 67272 277976 67324 277982
rect 67272 277918 67324 277924
rect 66904 277364 66956 277370
rect 66904 277306 66956 277312
rect 66916 276457 66944 277306
rect 66902 276448 66958 276457
rect 66902 276383 66958 276392
rect 66168 276072 66220 276078
rect 66168 276014 66220 276020
rect 66074 272368 66130 272377
rect 66074 272303 66130 272312
rect 65984 267096 66036 267102
rect 65984 267038 66036 267044
rect 65996 266665 66024 267038
rect 65982 266656 66038 266665
rect 65982 266591 66038 266600
rect 65890 240816 65946 240825
rect 65890 240751 65946 240760
rect 66088 161474 66116 272303
rect 66180 162761 66208 276014
rect 66444 275324 66496 275330
rect 66444 275266 66496 275272
rect 66456 274825 66484 275266
rect 66442 274816 66498 274825
rect 66442 274751 66498 274760
rect 66628 273284 66680 273290
rect 66628 273226 66680 273232
rect 66640 272377 66668 273226
rect 66810 273184 66866 273193
rect 66810 273119 66866 273128
rect 66626 272368 66682 272377
rect 66626 272303 66682 272312
rect 66824 271969 66852 273119
rect 66810 271960 66866 271969
rect 66810 271895 66866 271904
rect 66536 271176 66588 271182
rect 66536 271118 66588 271124
rect 66548 270745 66576 271118
rect 66534 270736 66590 270745
rect 66534 270671 66590 270680
rect 66812 270496 66864 270502
rect 66812 270438 66864 270444
rect 66824 269929 66852 270438
rect 66810 269920 66866 269929
rect 66810 269855 66866 269864
rect 66812 268388 66864 268394
rect 66812 268330 66864 268336
rect 66824 268297 66852 268330
rect 66810 268288 66866 268297
rect 66810 268223 66866 268232
rect 66810 265024 66866 265033
rect 66810 264959 66812 264968
rect 66864 264959 66866 264968
rect 66812 264930 66864 264936
rect 66626 264208 66682 264217
rect 66626 264143 66682 264152
rect 66640 263634 66668 264143
rect 66628 263628 66680 263634
rect 66628 263570 66680 263576
rect 67086 263392 67142 263401
rect 67086 263327 67142 263336
rect 66260 262880 66312 262886
rect 66260 262822 66312 262828
rect 66272 260953 66300 262822
rect 66902 262576 66958 262585
rect 66902 262511 66958 262520
rect 66916 262274 66944 262511
rect 66904 262268 66956 262274
rect 66904 262210 66956 262216
rect 67100 261526 67128 263327
rect 67088 261520 67140 261526
rect 67088 261462 67140 261468
rect 66258 260944 66314 260953
rect 66258 260879 66314 260888
rect 66272 260166 66300 260879
rect 66260 260160 66312 260166
rect 66260 260102 66312 260108
rect 66812 259412 66864 259418
rect 66812 259354 66864 259360
rect 66260 258732 66312 258738
rect 66260 258674 66312 258680
rect 66272 258058 66300 258674
rect 66824 258505 66852 259354
rect 66810 258496 66866 258505
rect 66810 258431 66866 258440
rect 66260 258052 66312 258058
rect 66260 257994 66312 258000
rect 66258 257680 66314 257689
rect 66258 257615 66314 257624
rect 66272 256766 66300 257615
rect 67376 256873 67404 324935
rect 67468 263401 67496 335326
rect 67548 291168 67600 291174
rect 67548 291110 67600 291116
rect 67560 281353 67588 291110
rect 67546 281344 67602 281353
rect 67546 281279 67602 281288
rect 67548 278724 67600 278730
rect 67548 278666 67600 278672
rect 67560 278089 67588 278666
rect 67546 278080 67602 278089
rect 67546 278015 67602 278024
rect 67548 277976 67600 277982
rect 67548 277918 67600 277924
rect 67454 263392 67510 263401
rect 67454 263327 67510 263336
rect 67362 256864 67418 256873
rect 67362 256799 67418 256808
rect 66260 256760 66312 256766
rect 66260 256702 66312 256708
rect 66810 255232 66866 255241
rect 66810 255167 66866 255176
rect 66824 254590 66852 255167
rect 66812 254584 66864 254590
rect 66812 254526 66864 254532
rect 66994 253600 67050 253609
rect 66994 253535 67050 253544
rect 67008 253230 67036 253535
rect 66996 253224 67048 253230
rect 66996 253166 67048 253172
rect 67272 253224 67324 253230
rect 67272 253166 67324 253172
rect 66810 251968 66866 251977
rect 66810 251903 66866 251912
rect 66824 251326 66852 251903
rect 66812 251320 66864 251326
rect 66812 251262 66864 251268
rect 66812 250572 66864 250578
rect 66812 250514 66864 250520
rect 66824 250345 66852 250514
rect 66810 250336 66866 250345
rect 66810 250271 66866 250280
rect 66444 249076 66496 249082
rect 66444 249018 66496 249024
rect 66456 248713 66484 249018
rect 66442 248704 66498 248713
rect 66442 248639 66498 248648
rect 66810 247888 66866 247897
rect 66810 247823 66866 247832
rect 66824 247110 66852 247823
rect 66812 247104 66864 247110
rect 66812 247046 66864 247052
rect 66718 243808 66774 243817
rect 66718 243743 66774 243752
rect 66732 242962 66760 243743
rect 66720 242956 66772 242962
rect 66720 242898 66772 242904
rect 66810 242176 66866 242185
rect 66810 242111 66866 242120
rect 66824 241534 66852 242111
rect 66812 241528 66864 241534
rect 66812 241470 66864 241476
rect 66166 162752 66222 162761
rect 66166 162687 66222 162696
rect 65996 161446 66116 161474
rect 65996 158030 66024 161446
rect 65984 158024 66036 158030
rect 65984 157966 66036 157972
rect 65892 140888 65944 140894
rect 65892 140830 65944 140836
rect 64788 137284 64840 137290
rect 64788 137226 64840 137232
rect 64786 137048 64842 137057
rect 64786 136983 64842 136992
rect 64694 136912 64750 136921
rect 64694 136847 64750 136856
rect 64604 133884 64656 133890
rect 64604 133826 64656 133832
rect 64512 118584 64564 118590
rect 64512 118526 64564 118532
rect 64708 103494 64736 136847
rect 64800 108934 64828 136983
rect 64788 108928 64840 108934
rect 64788 108870 64840 108876
rect 64788 105596 64840 105602
rect 64788 105538 64840 105544
rect 64696 103488 64748 103494
rect 64696 103430 64748 103436
rect 63408 102264 63460 102270
rect 63408 102206 63460 102212
rect 63408 99680 63460 99686
rect 63408 99622 63460 99628
rect 62028 99340 62080 99346
rect 62028 99282 62080 99288
rect 62764 96688 62816 96694
rect 62764 96630 62816 96636
rect 62776 79966 62804 96630
rect 63420 82793 63448 99622
rect 64800 83745 64828 105538
rect 65904 91050 65932 140830
rect 65996 121417 66024 157966
rect 66074 153232 66130 153241
rect 66074 153167 66130 153176
rect 65982 121408 66038 121417
rect 65982 121343 66038 121352
rect 66088 117065 66116 153167
rect 66180 126041 66208 162687
rect 67284 153338 67312 253166
rect 67272 153332 67324 153338
rect 67272 153274 67324 153280
rect 67180 137352 67232 137358
rect 67180 137294 67232 137300
rect 66812 133884 66864 133890
rect 66812 133826 66864 133832
rect 66824 133657 66852 133826
rect 66810 133648 66866 133657
rect 66810 133583 66866 133592
rect 66812 132456 66864 132462
rect 66812 132398 66864 132404
rect 66260 132388 66312 132394
rect 66260 132330 66312 132336
rect 66272 131209 66300 132330
rect 66824 132025 66852 132398
rect 66810 132016 66866 132025
rect 66810 131951 66866 131960
rect 66258 131200 66314 131209
rect 66258 131135 66314 131144
rect 67192 129849 67220 137294
rect 67178 129840 67234 129849
rect 67178 129775 67234 129784
rect 66812 128308 66864 128314
rect 66812 128250 66864 128256
rect 66824 128217 66852 128250
rect 66810 128208 66866 128217
rect 66810 128143 66866 128152
rect 66166 126032 66222 126041
rect 66166 125967 66222 125976
rect 66904 125588 66956 125594
rect 66904 125530 66956 125536
rect 66812 124908 66864 124914
rect 66812 124850 66864 124856
rect 66260 124160 66312 124166
rect 66260 124102 66312 124108
rect 66272 123049 66300 124102
rect 66824 123865 66852 124850
rect 66916 124409 66944 125530
rect 66902 124400 66958 124409
rect 66902 124335 66958 124344
rect 66810 123856 66866 123865
rect 66810 123791 66866 123800
rect 66258 123040 66314 123049
rect 66258 122975 66314 122984
rect 66352 122800 66404 122806
rect 66352 122742 66404 122748
rect 66364 122233 66392 122742
rect 66350 122224 66406 122233
rect 66350 122159 66406 122168
rect 66812 121440 66864 121446
rect 66812 121382 66864 121388
rect 66824 120601 66852 121382
rect 66902 120728 66958 120737
rect 66902 120663 66958 120672
rect 66810 120592 66866 120601
rect 66810 120527 66866 120536
rect 66812 120080 66864 120086
rect 66810 120048 66812 120057
rect 66864 120048 66866 120057
rect 66810 119983 66866 119992
rect 66916 119241 66944 120663
rect 66902 119232 66958 119241
rect 66902 119167 66958 119176
rect 66904 118652 66956 118658
rect 66904 118594 66956 118600
rect 66812 118584 66864 118590
rect 66812 118526 66864 118532
rect 66824 118425 66852 118526
rect 66810 118416 66866 118425
rect 66810 118351 66866 118360
rect 66916 117609 66944 118594
rect 66902 117600 66958 117609
rect 66902 117535 66958 117544
rect 66812 117224 66864 117230
rect 66812 117166 66864 117172
rect 66074 117056 66130 117065
rect 66074 116991 66130 117000
rect 66824 116249 66852 117166
rect 66810 116240 66866 116249
rect 66810 116175 66866 116184
rect 66812 115932 66864 115938
rect 66812 115874 66864 115880
rect 66824 115433 66852 115874
rect 66810 115424 66866 115433
rect 66810 115359 66866 115368
rect 66812 115320 66864 115326
rect 66812 115262 66864 115268
rect 66824 114617 66852 115262
rect 66810 114608 66866 114617
rect 66810 114543 66866 114552
rect 66812 114504 66864 114510
rect 66812 114446 66864 114452
rect 65984 113824 66036 113830
rect 66824 113801 66852 114446
rect 65984 113766 66036 113772
rect 66810 113792 66866 113801
rect 65996 113257 66024 113766
rect 66810 113727 66866 113736
rect 65982 113248 66038 113257
rect 65982 113183 66038 113192
rect 65892 91044 65944 91050
rect 65892 90986 65944 90992
rect 65996 85474 66024 113183
rect 66812 113144 66864 113150
rect 66812 113086 66864 113092
rect 66824 112441 66852 113086
rect 66904 113076 66956 113082
rect 66904 113018 66956 113024
rect 66810 112432 66866 112441
rect 66810 112367 66866 112376
rect 66812 111784 66864 111790
rect 66812 111726 66864 111732
rect 66824 110809 66852 111726
rect 66916 111625 66944 113018
rect 66902 111616 66958 111625
rect 66902 111551 66958 111560
rect 66810 110800 66866 110809
rect 66810 110735 66866 110744
rect 66812 110424 66864 110430
rect 66812 110366 66864 110372
rect 66824 109449 66852 110366
rect 66902 110256 66958 110265
rect 66902 110191 66958 110200
rect 66810 109440 66866 109449
rect 66810 109375 66866 109384
rect 66916 109070 66944 110191
rect 66904 109064 66956 109070
rect 66904 109006 66956 109012
rect 66720 108996 66772 109002
rect 66720 108938 66772 108944
rect 66444 108928 66496 108934
rect 66444 108870 66496 108876
rect 66456 108633 66484 108870
rect 66442 108624 66498 108633
rect 66442 108559 66498 108568
rect 66732 107817 66760 108938
rect 66718 107808 66774 107817
rect 66718 107743 66774 107752
rect 66994 106992 67050 107001
rect 66994 106927 66996 106936
rect 67048 106927 67050 106936
rect 66996 106898 67048 106904
rect 66534 105632 66590 105641
rect 66534 105567 66536 105576
rect 66588 105567 66590 105576
rect 66536 105538 66588 105544
rect 66352 104848 66404 104854
rect 66350 104816 66352 104825
rect 66404 104816 66406 104825
rect 66350 104751 66406 104760
rect 67284 104009 67312 153274
rect 67376 150657 67404 256799
rect 67454 246256 67510 246265
rect 67454 246191 67510 246200
rect 67468 233209 67496 246191
rect 67454 233200 67510 233209
rect 67454 233135 67510 233144
rect 67362 150648 67418 150657
rect 67362 150583 67418 150592
rect 67376 107001 67404 150583
rect 67362 106992 67418 107001
rect 67362 106927 67418 106936
rect 67270 104000 67326 104009
rect 67270 103935 67326 103944
rect 66628 103488 66680 103494
rect 66628 103430 66680 103436
rect 66534 103184 66590 103193
rect 66534 103119 66590 103128
rect 66548 102270 66576 103119
rect 66640 102649 66668 103430
rect 66626 102640 66682 102649
rect 66626 102575 66682 102584
rect 66076 102264 66128 102270
rect 66076 102206 66128 102212
rect 66536 102264 66588 102270
rect 66536 102206 66588 102212
rect 65984 85468 66036 85474
rect 65984 85410 66036 85416
rect 64786 83736 64842 83745
rect 64786 83671 64842 83680
rect 63406 82784 63462 82793
rect 63406 82719 63462 82728
rect 62764 79960 62816 79966
rect 62764 79902 62816 79908
rect 61936 74520 61988 74526
rect 61936 74462 61988 74468
rect 61948 73234 61976 74462
rect 61384 73228 61436 73234
rect 61384 73170 61436 73176
rect 61936 73228 61988 73234
rect 61936 73170 61988 73176
rect 61396 46238 61424 73170
rect 66088 70378 66116 102206
rect 67364 102196 67416 102202
rect 67364 102138 67416 102144
rect 66810 101824 66866 101833
rect 66810 101759 66866 101768
rect 66824 100910 66852 101759
rect 66812 100904 66864 100910
rect 66812 100846 66864 100852
rect 67270 100192 67326 100201
rect 67270 100127 67326 100136
rect 66812 99680 66864 99686
rect 66810 99648 66812 99657
rect 66864 99648 66866 99657
rect 66810 99583 66866 99592
rect 66812 99340 66864 99346
rect 66812 99282 66864 99288
rect 66824 98841 66852 99282
rect 66810 98832 66866 98841
rect 66810 98767 66866 98776
rect 66812 95192 66864 95198
rect 66812 95134 66864 95140
rect 66824 95033 66852 95134
rect 66810 95024 66866 95033
rect 66810 94959 66866 94968
rect 67284 88330 67312 100127
rect 67376 92886 67404 102138
rect 67468 97209 67496 233135
rect 67560 137358 67588 277918
rect 67652 242962 67680 354646
rect 67732 311160 67784 311166
rect 67732 311102 67784 311108
rect 67744 260137 67772 311102
rect 68664 296714 68692 383626
rect 69032 358766 69060 386990
rect 69124 368422 69152 390374
rect 69768 387054 69796 390374
rect 69756 387048 69808 387054
rect 69756 386990 69808 386996
rect 70400 387048 70452 387054
rect 70400 386990 70452 386996
rect 69112 368416 69164 368422
rect 69112 368358 69164 368364
rect 70412 362273 70440 386990
rect 70504 383489 70532 390374
rect 71240 387054 71268 390374
rect 72344 388482 72372 390374
rect 77206 390416 77262 390425
rect 72422 390351 72478 390360
rect 72528 390374 72864 390402
rect 73600 390374 73844 390402
rect 72422 389328 72478 389337
rect 72422 389263 72478 389272
rect 71688 388476 71740 388482
rect 71688 388418 71740 388424
rect 72332 388476 72384 388482
rect 72332 388418 72384 388424
rect 71700 387870 71728 388418
rect 71688 387864 71740 387870
rect 71688 387806 71740 387812
rect 71228 387048 71280 387054
rect 71228 386990 71280 386996
rect 71700 383625 71728 387806
rect 71686 383616 71742 383625
rect 71686 383551 71742 383560
rect 70490 383480 70546 383489
rect 70490 383415 70546 383424
rect 70398 362264 70454 362273
rect 70398 362199 70454 362208
rect 69020 358760 69072 358766
rect 69020 358702 69072 358708
rect 69664 358760 69716 358766
rect 69664 358702 69716 358708
rect 68572 296686 68692 296714
rect 68572 291174 68600 296686
rect 68560 291168 68612 291174
rect 69676 291145 69704 358702
rect 71044 311228 71096 311234
rect 71044 311170 71096 311176
rect 70306 307864 70362 307873
rect 70306 307799 70362 307808
rect 68560 291110 68612 291116
rect 69662 291136 69718 291145
rect 69662 291071 69718 291080
rect 69018 288552 69074 288561
rect 69018 288487 69074 288496
rect 69032 284442 69060 288487
rect 69846 287192 69902 287201
rect 69846 287127 69902 287136
rect 69020 284436 69072 284442
rect 69020 284378 69072 284384
rect 69032 283778 69060 284378
rect 68986 283750 69060 283778
rect 68986 283492 69014 283750
rect 67822 283248 67878 283257
rect 67822 283183 67878 283192
rect 67836 277273 67864 283183
rect 69860 283098 69888 287127
rect 70320 284374 70348 307799
rect 70492 287700 70544 287706
rect 70492 287642 70544 287648
rect 70308 284368 70360 284374
rect 70308 284310 70360 284316
rect 70320 283506 70348 284310
rect 70104 283478 70348 283506
rect 70504 283370 70532 287642
rect 71056 283506 71084 311170
rect 71596 289196 71648 289202
rect 71596 289138 71648 289144
rect 71608 283529 71636 289138
rect 72436 283665 72464 389263
rect 72528 387870 72556 390374
rect 72516 387864 72568 387870
rect 72516 387806 72568 387812
rect 73066 387016 73122 387025
rect 73066 386951 73122 386960
rect 73080 345778 73108 386951
rect 73816 384334 73844 390374
rect 73908 390374 74336 390402
rect 74644 390374 75072 390402
rect 75288 390374 75624 390402
rect 75932 390374 76360 390402
rect 77096 390374 77206 390402
rect 73804 384328 73856 384334
rect 73804 384270 73856 384276
rect 73908 383654 73936 390374
rect 74540 387048 74592 387054
rect 74540 386990 74592 386996
rect 73172 383626 73936 383654
rect 73172 371249 73200 383626
rect 73802 382936 73858 382945
rect 73802 382871 73858 382880
rect 73158 371240 73214 371249
rect 73158 371175 73214 371184
rect 72516 345772 72568 345778
rect 72516 345714 72568 345720
rect 73068 345772 73120 345778
rect 73068 345714 73120 345720
rect 72528 345098 72556 345714
rect 72516 345092 72568 345098
rect 72516 345034 72568 345040
rect 72528 288454 72556 345034
rect 72700 302932 72752 302938
rect 72700 302874 72752 302880
rect 72516 288448 72568 288454
rect 72516 288390 72568 288396
rect 71870 283656 71926 283665
rect 71870 283591 71926 283600
rect 72422 283656 72478 283665
rect 72422 283591 72478 283600
rect 71594 283520 71650 283529
rect 71056 283478 71208 283506
rect 70504 283356 70656 283370
rect 70504 283342 70670 283356
rect 69216 283082 69888 283098
rect 68836 283076 68888 283082
rect 68836 283018 68888 283024
rect 69204 283076 69888 283082
rect 69256 283070 69888 283076
rect 69204 283018 69256 283024
rect 68848 277394 68876 283018
rect 70642 282962 70670 283342
rect 70768 283008 70820 283014
rect 70642 282956 70768 282962
rect 70642 282950 70820 282956
rect 70858 282976 70914 282985
rect 70642 282948 70808 282950
rect 70656 282934 70808 282948
rect 71056 282962 71084 283478
rect 71594 283455 71650 283464
rect 71608 283234 71636 283455
rect 71884 283257 71912 283591
rect 71962 283520 72018 283529
rect 72712 283506 72740 302874
rect 72792 288448 72844 288454
rect 72792 288390 72844 288396
rect 72804 283778 72832 288390
rect 73816 285841 73844 382871
rect 74552 353258 74580 386990
rect 74644 361486 74672 390374
rect 75288 387054 75316 390374
rect 75276 387048 75328 387054
rect 75276 386990 75328 386996
rect 74632 361480 74684 361486
rect 74632 361422 74684 361428
rect 75932 356046 75960 390374
rect 77206 390351 77262 390360
rect 77312 390374 77832 390402
rect 78048 390374 78384 390402
rect 77220 388793 77248 390351
rect 77206 388784 77262 388793
rect 77206 388719 77262 388728
rect 77208 385824 77260 385830
rect 77208 385766 77260 385772
rect 77220 369209 77248 385766
rect 77312 380798 77340 390374
rect 77482 388512 77538 388521
rect 77482 388447 77538 388456
rect 77300 380792 77352 380798
rect 77300 380734 77352 380740
rect 77206 369200 77262 369209
rect 77206 369135 77262 369144
rect 75920 356040 75972 356046
rect 75920 355982 75972 355988
rect 76564 356040 76616 356046
rect 76564 355982 76616 355988
rect 74540 353252 74592 353258
rect 74540 353194 74592 353200
rect 76288 305652 76340 305658
rect 76288 305594 76340 305600
rect 74630 288688 74686 288697
rect 74630 288623 74686 288632
rect 73896 287088 73948 287094
rect 73896 287030 73948 287036
rect 73802 285832 73858 285841
rect 73802 285767 73858 285776
rect 72804 283750 72878 283778
rect 72018 283478 72740 283506
rect 72850 283492 72878 283750
rect 73250 283520 73306 283529
rect 71962 283455 72018 283464
rect 73816 283506 73844 285767
rect 73908 284209 73936 287030
rect 73894 284200 73950 284209
rect 73894 284135 73950 284144
rect 74644 283506 74672 288623
rect 74724 286408 74776 286414
rect 74724 286350 74776 286356
rect 73306 283478 73416 283506
rect 73816 283478 73968 283506
rect 74520 283478 74672 283506
rect 74736 283506 74764 286350
rect 75736 286340 75788 286346
rect 75736 286282 75788 286288
rect 75748 283506 75776 286282
rect 76150 283756 76202 283762
rect 76150 283698 76202 283704
rect 74736 283478 75072 283506
rect 75624 283478 75776 283506
rect 75826 283520 75882 283529
rect 73250 283455 73306 283464
rect 76162 283506 76190 283698
rect 75882 283492 76190 283506
rect 76300 283506 76328 305594
rect 76576 284209 76604 355982
rect 77496 311234 77524 388447
rect 78048 385830 78076 390374
rect 78680 387048 78732 387054
rect 78680 386990 78732 386996
rect 78036 385824 78088 385830
rect 78036 385766 78088 385772
rect 78586 385112 78642 385121
rect 78586 385047 78642 385056
rect 77484 311228 77536 311234
rect 77484 311170 77536 311176
rect 76654 309088 76710 309097
rect 76654 309023 76710 309032
rect 76562 284200 76618 284209
rect 76562 284135 76618 284144
rect 76668 283762 76696 309023
rect 77298 306504 77354 306513
rect 77298 306439 77354 306448
rect 77312 283778 77340 306439
rect 78600 296714 78628 385047
rect 78508 296686 78628 296714
rect 78508 292574 78536 296686
rect 78232 292546 78536 292574
rect 78232 284442 78260 292546
rect 78588 287700 78640 287706
rect 78588 287642 78640 287648
rect 78220 284436 78272 284442
rect 78220 284378 78272 284384
rect 76656 283756 76708 283762
rect 76656 283698 76708 283704
rect 77266 283750 77340 283778
rect 75882 283478 76176 283492
rect 76300 283478 76728 283506
rect 77266 283492 77294 283750
rect 78232 283506 78260 284378
rect 78600 283506 78628 287642
rect 78692 284209 78720 386990
rect 78770 386880 78826 386889
rect 78770 386815 78826 386824
rect 78784 306374 78812 386815
rect 79428 384985 79456 390510
rect 79520 390374 79856 390402
rect 80592 390374 80928 390402
rect 79520 387054 79548 390374
rect 80058 390144 80114 390153
rect 80058 390079 80114 390088
rect 79508 387048 79560 387054
rect 79508 386990 79560 386996
rect 79414 384976 79470 384985
rect 79414 384911 79470 384920
rect 78784 306346 79088 306374
rect 78956 289128 79008 289134
rect 78956 289070 79008 289076
rect 78678 284200 78734 284209
rect 78678 284135 78734 284144
rect 78968 283778 78996 289070
rect 77832 283478 78260 283506
rect 78384 283478 78628 283506
rect 78922 283750 78996 283778
rect 78922 283492 78950 283750
rect 79060 283529 79088 306346
rect 79966 293176 80022 293185
rect 79966 293111 80022 293120
rect 79980 289134 80008 293111
rect 80072 291145 80100 390079
rect 80900 385801 80928 390374
rect 81314 390153 81342 390388
rect 82004 390374 82616 390402
rect 81300 390144 81356 390153
rect 81300 390079 81356 390088
rect 80886 385792 80942 385801
rect 80886 385727 80942 385736
rect 80702 378720 80758 378729
rect 80702 378655 80758 378664
rect 80058 291136 80114 291145
rect 80058 291071 80114 291080
rect 79968 289128 80020 289134
rect 79968 289070 80020 289076
rect 80716 288386 80744 378655
rect 82004 376417 82032 390374
rect 82726 387560 82782 387569
rect 82726 387495 82782 387504
rect 81990 376408 82046 376417
rect 81990 376343 82046 376352
rect 82004 373994 82032 376343
rect 82004 373966 82124 373994
rect 80794 311128 80850 311137
rect 80794 311063 80850 311072
rect 80808 306374 80836 311063
rect 80808 306346 81020 306374
rect 80060 288380 80112 288386
rect 80060 288322 80112 288328
rect 80704 288380 80756 288386
rect 80704 288322 80756 288328
rect 80072 287094 80100 288322
rect 80060 287088 80112 287094
rect 80060 287030 80112 287036
rect 80072 283778 80100 287030
rect 80992 285802 81020 306346
rect 82096 291145 82124 373966
rect 82634 304192 82690 304201
rect 82634 304127 82690 304136
rect 82648 292602 82676 304127
rect 82176 292596 82228 292602
rect 82176 292538 82228 292544
rect 82636 292596 82688 292602
rect 82636 292538 82688 292544
rect 82082 291136 82138 291145
rect 82082 291071 82138 291080
rect 80980 285796 81032 285802
rect 80980 285738 81032 285744
rect 80888 285728 80940 285734
rect 80888 285670 80940 285676
rect 80026 283750 80100 283778
rect 79046 283520 79102 283529
rect 75826 283455 75882 283464
rect 79102 283478 79488 283506
rect 80026 283492 80054 283750
rect 80900 283506 80928 285670
rect 80592 283478 80928 283506
rect 80992 283506 81020 285738
rect 82188 285734 82216 292538
rect 82740 287054 82768 387495
rect 83200 386986 83228 390623
rect 83476 390374 84088 390402
rect 84824 390374 85160 390402
rect 83188 386980 83240 386986
rect 83188 386922 83240 386928
rect 82820 373994 82872 373998
rect 83476 373994 83504 390374
rect 84108 386980 84160 386986
rect 84108 386922 84160 386928
rect 82820 373992 83504 373994
rect 82872 373966 83504 373992
rect 82820 373934 82872 373940
rect 84120 360126 84148 386922
rect 85132 386306 85160 390374
rect 85362 390130 85390 390388
rect 85362 390102 85436 390130
rect 85120 386300 85172 386306
rect 85120 386242 85172 386248
rect 85408 385898 85436 390102
rect 85396 385892 85448 385898
rect 85396 385834 85448 385840
rect 84108 360120 84160 360126
rect 84108 360062 84160 360068
rect 82910 346488 82966 346497
rect 82910 346423 82966 346432
rect 82924 306374 82952 346423
rect 85500 320142 85528 390895
rect 92018 390824 92074 390833
rect 92074 390782 92368 390810
rect 92018 390759 92074 390768
rect 89718 390688 89774 390697
rect 89608 390646 89718 390674
rect 89774 390658 89944 390674
rect 89774 390652 89956 390658
rect 89774 390646 89904 390652
rect 89718 390623 89774 390632
rect 89732 390563 89760 390623
rect 89904 390594 89956 390600
rect 90456 390652 90508 390658
rect 90456 390594 90508 390600
rect 87984 390510 88136 390538
rect 85592 390374 86112 390402
rect 85592 382265 85620 390374
rect 86834 390130 86862 390388
rect 86972 390374 87584 390402
rect 86834 390102 86908 390130
rect 86880 387122 86908 390102
rect 86868 387116 86920 387122
rect 86868 387058 86920 387064
rect 86866 382936 86922 382945
rect 86866 382871 86922 382880
rect 85578 382256 85634 382265
rect 85578 382191 85634 382200
rect 84844 320136 84896 320142
rect 84844 320078 84896 320084
rect 85488 320136 85540 320142
rect 85488 320078 85540 320084
rect 84106 312488 84162 312497
rect 84106 312423 84162 312432
rect 84014 308408 84070 308417
rect 84014 308343 84070 308352
rect 82924 306346 83412 306374
rect 82648 287026 82768 287054
rect 82360 286272 82412 286278
rect 82360 286214 82412 286220
rect 82176 285728 82228 285734
rect 82176 285670 82228 285676
rect 80992 283478 81144 283506
rect 79046 283455 79102 283464
rect 79060 283395 79088 283455
rect 71870 283248 71926 283257
rect 71608 283206 71760 283234
rect 71870 283183 71926 283192
rect 81990 283112 82046 283121
rect 82372 283098 82400 286214
rect 82046 283070 82400 283098
rect 81990 283047 82046 283056
rect 82648 282985 82676 287026
rect 83094 285832 83150 285841
rect 83094 285767 83150 285776
rect 83108 283506 83136 285767
rect 83384 283778 83412 306346
rect 83462 305824 83518 305833
rect 83462 305759 83518 305768
rect 83476 286278 83504 305759
rect 83464 286272 83516 286278
rect 83464 286214 83516 286220
rect 84028 285841 84056 308343
rect 84014 285832 84070 285841
rect 84014 285767 84070 285776
rect 84120 285705 84148 312423
rect 84856 305658 84884 320078
rect 86774 313984 86830 313993
rect 86774 313919 86830 313928
rect 84844 305652 84896 305658
rect 84844 305594 84896 305600
rect 86224 291644 86276 291650
rect 86224 291586 86276 291592
rect 84568 289876 84620 289882
rect 84568 289818 84620 289824
rect 84292 285728 84344 285734
rect 84106 285696 84162 285705
rect 84292 285670 84344 285676
rect 84106 285631 84162 285640
rect 83384 283750 83504 283778
rect 82800 283478 83136 283506
rect 83476 283506 83504 283750
rect 83476 283478 83904 283506
rect 84304 283234 84332 285670
rect 84580 283506 84608 289818
rect 85856 287972 85908 287978
rect 85856 287914 85908 287920
rect 85868 283506 85896 287914
rect 84580 283478 85008 283506
rect 85560 283478 85896 283506
rect 86236 283506 86264 291586
rect 86788 287978 86816 313919
rect 86776 287972 86828 287978
rect 86776 287914 86828 287920
rect 86788 287094 86816 287914
rect 86776 287088 86828 287094
rect 86776 287030 86828 287036
rect 86880 285705 86908 382871
rect 86972 307737 87000 390374
rect 87984 389201 88012 390510
rect 88352 390374 88872 390402
rect 89732 390374 90344 390402
rect 87970 389192 88026 389201
rect 87970 389127 88026 389136
rect 88248 375352 88300 375358
rect 88248 375294 88300 375300
rect 88260 316810 88288 375294
rect 88352 373289 88380 390374
rect 89626 385928 89682 385937
rect 88432 385892 88484 385898
rect 89626 385863 89682 385872
rect 88432 385834 88484 385840
rect 88338 373280 88394 373289
rect 88338 373215 88394 373224
rect 87604 316804 87656 316810
rect 87604 316746 87656 316752
rect 88248 316804 88300 316810
rect 88248 316746 88300 316752
rect 87616 316062 87644 316746
rect 87604 316056 87656 316062
rect 87604 315998 87656 316004
rect 86958 307728 87014 307737
rect 86958 307663 87014 307672
rect 86960 296064 87012 296070
rect 86960 296006 87012 296012
rect 86866 285696 86922 285705
rect 86866 285631 86922 285640
rect 86972 283506 87000 296006
rect 87326 291136 87382 291145
rect 87326 291071 87382 291080
rect 87340 289921 87368 291071
rect 87616 290465 87644 315998
rect 88246 307048 88302 307057
rect 88246 306983 88302 306992
rect 88260 291145 88288 306983
rect 88444 294681 88472 385834
rect 89442 316704 89498 316713
rect 89442 316639 89498 316648
rect 88430 294672 88486 294681
rect 88430 294607 88486 294616
rect 88246 291136 88302 291145
rect 88246 291071 88302 291080
rect 87602 290456 87658 290465
rect 87602 290391 87658 290400
rect 87326 289912 87382 289921
rect 87326 289847 87382 289856
rect 87340 283506 87368 289847
rect 88614 287872 88670 287881
rect 88614 287807 88670 287816
rect 86236 283478 86664 283506
rect 86972 283478 87216 283506
rect 87340 283478 87768 283506
rect 84304 283206 84456 283234
rect 88430 283112 88486 283121
rect 88320 283070 88430 283098
rect 88628 283098 88656 287807
rect 89456 287054 89484 316639
rect 89180 287026 89484 287054
rect 89180 285977 89208 287026
rect 89166 285968 89222 285977
rect 89166 285903 89222 285912
rect 89180 283506 89208 285903
rect 88872 283478 89208 283506
rect 88486 283070 88656 283098
rect 88430 283047 88486 283056
rect 81990 282976 82046 282985
rect 70914 282934 71084 282962
rect 81696 282934 81990 282962
rect 70858 282911 70914 282920
rect 81990 282911 82046 282920
rect 82634 282976 82690 282985
rect 83462 282976 83518 282985
rect 83352 282934 83462 282962
rect 82634 282911 82690 282920
rect 86314 282976 86370 282985
rect 86112 282934 86314 282962
rect 83462 282911 83518 282920
rect 86314 282911 86370 282920
rect 89074 282976 89130 282985
rect 89640 282962 89668 385863
rect 89732 289649 89760 390374
rect 90468 388929 90496 390594
rect 91066 390130 91094 390388
rect 91204 390374 91632 390402
rect 91066 390102 91140 390130
rect 90454 388920 90510 388929
rect 90454 388855 90510 388864
rect 91112 384305 91140 390102
rect 91098 384296 91154 384305
rect 91098 384231 91154 384240
rect 91204 373994 91232 390374
rect 92032 389174 92060 390759
rect 93104 390374 93440 390402
rect 91940 389146 92060 389174
rect 91940 375358 91968 389146
rect 93412 387569 93440 390374
rect 93964 388346 93992 390918
rect 99470 390895 99526 390904
rect 106002 390960 106058 390969
rect 107382 390960 107438 390969
rect 106058 390918 106136 390946
rect 107088 390918 107382 390946
rect 106002 390895 106058 390904
rect 96802 390824 96858 390833
rect 96600 390782 96802 390810
rect 97078 390824 97134 390833
rect 96858 390782 96936 390810
rect 96802 390759 96858 390768
rect 94148 390374 94392 390402
rect 94792 390374 95128 390402
rect 95252 390374 95864 390402
rect 93952 388340 94004 388346
rect 93952 388282 94004 388288
rect 93398 387560 93454 387569
rect 93398 387495 93454 387504
rect 94148 387138 94176 390374
rect 94228 388340 94280 388346
rect 94228 388282 94280 388288
rect 93872 387110 94176 387138
rect 93124 384328 93176 384334
rect 93124 384270 93176 384276
rect 91928 375352 91980 375358
rect 91928 375294 91980 375300
rect 91112 373966 91232 373994
rect 91006 311128 91062 311137
rect 91006 311063 91062 311072
rect 90362 305688 90418 305697
rect 90362 305623 90418 305632
rect 89718 289640 89774 289649
rect 89718 289575 89774 289584
rect 90270 286104 90326 286113
rect 90270 286039 90326 286048
rect 89810 283520 89866 283529
rect 90284 283506 90312 286039
rect 90376 285734 90404 305623
rect 91020 286113 91048 311063
rect 91112 301617 91140 373966
rect 93136 365702 93164 384270
rect 93124 365696 93176 365702
rect 93124 365638 93176 365644
rect 93872 362234 93900 387110
rect 93952 386912 94004 386918
rect 93952 386854 94004 386860
rect 93964 372502 93992 386854
rect 94240 376718 94268 388282
rect 94792 386918 94820 390374
rect 94780 386912 94832 386918
rect 94780 386854 94832 386860
rect 95146 382392 95202 382401
rect 95146 382327 95202 382336
rect 94228 376712 94280 376718
rect 94228 376654 94280 376660
rect 93952 372496 94004 372502
rect 93952 372438 94004 372444
rect 93860 362228 93912 362234
rect 93860 362170 93912 362176
rect 95160 342310 95188 382327
rect 95148 342304 95200 342310
rect 95148 342246 95200 342252
rect 94504 330540 94556 330546
rect 94504 330482 94556 330488
rect 94516 318102 94544 330482
rect 94504 318096 94556 318102
rect 94504 318038 94556 318044
rect 93766 315344 93822 315353
rect 93766 315279 93822 315288
rect 92480 312588 92532 312594
rect 92480 312530 92532 312536
rect 92388 305652 92440 305658
rect 92388 305594 92440 305600
rect 91098 301608 91154 301617
rect 91098 301543 91154 301552
rect 92296 301572 92348 301578
rect 92296 301514 92348 301520
rect 91928 287020 91980 287026
rect 91928 286962 91980 286968
rect 91006 286104 91062 286113
rect 91006 286039 91062 286048
rect 91376 285932 91428 285938
rect 91376 285874 91428 285880
rect 90364 285728 90416 285734
rect 90364 285670 90416 285676
rect 91388 283506 91416 285874
rect 91940 283506 91968 286962
rect 92308 284209 92336 301514
rect 92400 287026 92428 305594
rect 92492 287774 92520 312530
rect 93124 307080 93176 307086
rect 93124 307022 93176 307028
rect 92572 293956 92624 293962
rect 92572 293898 92624 293904
rect 92480 287768 92532 287774
rect 92480 287710 92532 287716
rect 92388 287020 92440 287026
rect 92388 286962 92440 286968
rect 92294 284200 92350 284209
rect 92294 284135 92350 284144
rect 92386 283656 92442 283665
rect 92386 283591 92442 283600
rect 92400 283506 92428 283591
rect 89866 283478 90312 283506
rect 91080 283478 91416 283506
rect 91632 283478 91968 283506
rect 92184 283478 92428 283506
rect 92584 283506 92612 293898
rect 93136 291650 93164 307022
rect 93780 293962 93808 315279
rect 94502 309768 94558 309777
rect 94502 309703 94558 309712
rect 93768 293956 93820 293962
rect 93768 293898 93820 293904
rect 93124 291644 93176 291650
rect 93124 291586 93176 291592
rect 92940 287768 92992 287774
rect 92940 287710 92992 287716
rect 92952 283506 92980 287710
rect 93950 284336 94006 284345
rect 93950 284271 94006 284280
rect 93964 283506 93992 284271
rect 92584 283478 92736 283506
rect 92952 283478 93288 283506
rect 93840 283478 93992 283506
rect 94042 283520 94098 283529
rect 89810 283455 89866 283464
rect 94516 283506 94544 309703
rect 94596 301504 94648 301510
rect 94596 301446 94648 301452
rect 94608 285938 94636 301446
rect 94596 285932 94648 285938
rect 94596 285874 94648 285880
rect 95160 283506 95188 342246
rect 95252 290057 95280 390374
rect 96712 390176 96764 390182
rect 96712 390118 96764 390124
rect 96724 373994 96752 390118
rect 96908 389065 96936 390782
rect 97134 390782 97764 390810
rect 97078 390759 97134 390768
rect 96894 389056 96950 389065
rect 96894 388991 96950 389000
rect 97630 389056 97686 389065
rect 97630 388991 97686 389000
rect 97262 377496 97318 377505
rect 97644 377466 97672 388991
rect 97736 382974 97764 390782
rect 99484 390538 99512 390895
rect 100392 390584 100444 390590
rect 99360 390510 99604 390538
rect 100096 390532 100392 390538
rect 100096 390526 100444 390532
rect 100096 390510 100432 390526
rect 97874 390182 97902 390388
rect 98624 390374 98960 390402
rect 97862 390176 97914 390182
rect 97862 390118 97914 390124
rect 98932 389201 98960 390374
rect 98918 389192 98974 389201
rect 98918 389127 98974 389136
rect 99470 387968 99526 387977
rect 99470 387903 99526 387912
rect 97724 382968 97776 382974
rect 97724 382910 97776 382916
rect 97262 377431 97318 377440
rect 97632 377460 97684 377466
rect 96632 373966 96752 373994
rect 95330 312488 95386 312497
rect 95330 312423 95386 312432
rect 95344 306374 95372 312423
rect 95344 306346 95648 306374
rect 95238 290048 95294 290057
rect 95238 289983 95294 289992
rect 95332 286748 95384 286754
rect 95332 286690 95384 286696
rect 94098 283478 94544 283506
rect 94700 283478 95188 283506
rect 94042 283455 94098 283464
rect 94700 283393 94728 283478
rect 94686 283384 94742 283393
rect 94686 283319 94742 283328
rect 95344 283234 95372 286690
rect 95620 283506 95648 306346
rect 96632 301578 96660 373966
rect 97276 366994 97304 377431
rect 97632 377402 97684 377408
rect 99286 370560 99342 370569
rect 99286 370495 99342 370504
rect 98368 367804 98420 367810
rect 98368 367746 98420 367752
rect 97264 366988 97316 366994
rect 97264 366930 97316 366936
rect 96712 325712 96764 325718
rect 96712 325654 96764 325660
rect 96620 301572 96672 301578
rect 96620 301514 96672 301520
rect 96724 283506 96752 325654
rect 97264 308440 97316 308446
rect 97264 308382 97316 308388
rect 97172 304292 97224 304298
rect 97172 304234 97224 304240
rect 97184 285818 97212 304234
rect 97276 286754 97304 308382
rect 98276 291236 98328 291242
rect 98276 291178 98328 291184
rect 97264 286748 97316 286754
rect 97264 286690 97316 286696
rect 97184 285790 97304 285818
rect 97276 283506 97304 285790
rect 98288 283778 98316 291178
rect 98242 283750 98316 283778
rect 95620 283478 96048 283506
rect 96724 283478 97152 283506
rect 97276 283478 97704 283506
rect 98242 283492 98270 283750
rect 96894 283384 96950 283393
rect 96600 283342 96894 283370
rect 96894 283319 96950 283328
rect 95344 283206 95496 283234
rect 90730 282976 90786 282985
rect 89130 282934 89668 282962
rect 90528 282934 90730 282962
rect 89074 282911 89130 282920
rect 90730 282911 90786 282920
rect 68848 277366 68968 277394
rect 67822 277264 67878 277273
rect 67822 277199 67878 277208
rect 67836 276078 67864 277199
rect 67824 276072 67876 276078
rect 67824 276014 67876 276020
rect 67730 260128 67786 260137
rect 67730 260063 67786 260072
rect 67744 259486 67772 260063
rect 67732 259480 67784 259486
rect 67732 259422 67784 259428
rect 68190 258768 68246 258777
rect 68190 258703 68246 258712
rect 68204 258058 68232 258703
rect 68192 258052 68244 258058
rect 68192 257994 68244 258000
rect 67730 251152 67786 251161
rect 67730 251087 67786 251096
rect 67640 242956 67692 242962
rect 67640 242898 67692 242904
rect 67548 137352 67600 137358
rect 67548 137294 67600 137300
rect 67652 102202 67680 242898
rect 67744 234054 67772 251087
rect 67822 249520 67878 249529
rect 67822 249455 67878 249464
rect 67836 238746 67864 249455
rect 68468 242956 68520 242962
rect 68468 242898 68520 242904
rect 68480 242298 68508 242898
rect 68480 242270 68816 242298
rect 67824 238740 67876 238746
rect 67824 238682 67876 238688
rect 67732 234048 67784 234054
rect 67732 233990 67784 233996
rect 68940 167074 68968 277366
rect 98380 258777 98408 367746
rect 99196 307148 99248 307154
rect 99196 307090 99248 307096
rect 99208 292574 99236 307090
rect 99024 292546 99236 292574
rect 99024 283506 99052 292546
rect 99300 291242 99328 370495
rect 99484 316713 99512 387903
rect 99576 385694 99604 390510
rect 100666 390416 100722 390425
rect 104254 390416 104310 390425
rect 100722 390388 100832 390402
rect 100722 390374 100846 390388
rect 100666 390351 100722 390360
rect 100818 390182 100846 390374
rect 101048 390374 101384 390402
rect 102120 390374 102272 390402
rect 102856 390374 103468 390402
rect 103592 390374 103928 390402
rect 104144 390374 104254 390402
rect 100806 390176 100858 390182
rect 100772 390124 100806 390130
rect 100772 390118 100858 390124
rect 100772 390102 100846 390118
rect 100772 389298 100800 390102
rect 100760 389292 100812 389298
rect 100760 389234 100812 389240
rect 99564 385688 99616 385694
rect 99564 385630 99616 385636
rect 101048 373994 101076 390374
rect 101956 390176 102008 390182
rect 101956 390118 102008 390124
rect 100772 373966 101076 373994
rect 100772 354006 100800 373966
rect 101968 369850 101996 390118
rect 102048 381540 102100 381546
rect 102048 381482 102100 381488
rect 101956 369844 102008 369850
rect 101956 369786 102008 369792
rect 100760 354000 100812 354006
rect 100760 353942 100812 353948
rect 101404 341556 101456 341562
rect 101404 341498 101456 341504
rect 99470 316704 99526 316713
rect 99470 316639 99526 316648
rect 99288 291236 99340 291242
rect 99288 291178 99340 291184
rect 100114 289912 100170 289921
rect 100114 289847 100170 289856
rect 100024 284436 100076 284442
rect 100024 284378 100076 284384
rect 99104 284368 99156 284374
rect 99104 284310 99156 284316
rect 98624 283478 99052 283506
rect 98736 283008 98788 283014
rect 98736 282950 98788 282956
rect 98918 282976 98974 282985
rect 98748 280158 98776 282950
rect 98918 282911 98974 282920
rect 98736 280152 98788 280158
rect 98736 280094 98788 280100
rect 98932 279970 98960 282911
rect 98748 279942 98960 279970
rect 98748 264246 98776 279942
rect 99116 277394 99144 284310
rect 99380 282940 99432 282946
rect 99380 282882 99432 282888
rect 99392 281518 99420 282882
rect 99380 281512 99432 281518
rect 99380 281454 99432 281460
rect 98840 277366 99144 277394
rect 98840 269822 98868 277366
rect 99470 271280 99526 271289
rect 99470 271215 99526 271224
rect 98828 269816 98880 269822
rect 98828 269758 98880 269764
rect 98736 264240 98788 264246
rect 98736 264182 98788 264188
rect 99378 259040 99434 259049
rect 99378 258975 99434 258984
rect 98366 258768 98422 258777
rect 98366 258703 98422 258712
rect 98380 258194 98408 258703
rect 98368 258188 98420 258194
rect 98368 258130 98420 258136
rect 98736 251184 98788 251190
rect 98736 251126 98788 251132
rect 98090 247072 98146 247081
rect 98090 247007 98146 247016
rect 71134 241768 71190 241777
rect 70840 241726 71134 241754
rect 74906 241768 74962 241777
rect 71134 241703 71190 241712
rect 74828 241726 74906 241754
rect 74828 241618 74856 241726
rect 76654 241768 76710 241777
rect 76360 241726 76654 241754
rect 74906 241703 74962 241712
rect 77666 241768 77722 241777
rect 76654 241703 76710 241712
rect 77312 241726 77666 241754
rect 69184 241590 69520 241618
rect 69294 241496 69350 241505
rect 69294 241431 69350 241440
rect 69020 240032 69072 240038
rect 69020 239974 69072 239980
rect 69032 209098 69060 239974
rect 69308 219434 69336 241431
rect 69492 240310 69520 241590
rect 69584 241590 69736 241618
rect 69952 241590 70288 241618
rect 71332 241590 71392 241618
rect 71792 241590 71944 241618
rect 72496 241590 72832 241618
rect 69584 241505 69612 241590
rect 69570 241496 69626 241505
rect 69570 241431 69626 241440
rect 69480 240304 69532 240310
rect 69480 240246 69532 240252
rect 69952 240038 69980 241590
rect 71332 241505 71360 241590
rect 71318 241496 71374 241505
rect 71318 241431 71374 241440
rect 71332 240038 71360 241431
rect 71792 240145 71820 241590
rect 71778 240136 71834 240145
rect 71778 240071 71834 240080
rect 69940 240032 69992 240038
rect 69940 239974 69992 239980
rect 70492 240032 70544 240038
rect 70492 239974 70544 239980
rect 71320 240032 71372 240038
rect 71320 239974 71372 239980
rect 69124 219406 69336 219434
rect 69020 209092 69072 209098
rect 69020 209034 69072 209040
rect 67732 167068 67784 167074
rect 67732 167010 67784 167016
rect 68928 167068 68980 167074
rect 68928 167010 68980 167016
rect 67744 132841 67772 167010
rect 67824 156664 67876 156670
rect 67824 156606 67876 156612
rect 68652 156664 68704 156670
rect 68652 156606 68704 156612
rect 67730 132832 67786 132841
rect 67730 132767 67786 132776
rect 67730 129024 67786 129033
rect 67730 128959 67786 128968
rect 67640 102196 67692 102202
rect 67640 102138 67692 102144
rect 67546 98016 67602 98025
rect 67546 97951 67602 97960
rect 67454 97200 67510 97209
rect 67454 97135 67510 97144
rect 67364 92880 67416 92886
rect 67364 92822 67416 92828
rect 67468 92342 67496 97135
rect 67456 92336 67508 92342
rect 67456 92278 67508 92284
rect 67272 88324 67324 88330
rect 67272 88266 67324 88272
rect 67560 86737 67588 97951
rect 67546 86728 67602 86737
rect 67546 86663 67602 86672
rect 66076 70372 66128 70378
rect 66076 70314 66128 70320
rect 61384 46232 61436 46238
rect 60738 46200 60794 46209
rect 61384 46174 61436 46180
rect 60738 46135 60794 46144
rect 57244 33108 57296 33114
rect 57244 33050 57296 33056
rect 59360 24132 59412 24138
rect 59360 24074 59412 24080
rect 57980 21412 58032 21418
rect 57980 21354 58032 21360
rect 57992 16574 58020 21354
rect 59372 16574 59400 24074
rect 60752 16574 60780 46135
rect 64880 44872 64932 44878
rect 64880 44814 64932 44820
rect 63500 18624 63552 18630
rect 63500 18566 63552 18572
rect 63512 16574 63540 18566
rect 64892 16574 64920 44814
rect 66260 42084 66312 42090
rect 66260 42026 66312 42032
rect 66272 16574 66300 42026
rect 67640 28280 67692 28286
rect 67640 28222 67692 28228
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 59372 16546 59676 16574
rect 60752 16546 60872 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 52472 6886 52592 6914
rect 51356 2100 51408 2106
rect 51356 2042 51408 2048
rect 51368 480 51396 2042
rect 52564 480 52592 6886
rect 53300 490 53328 16546
rect 53576 598 53788 626
rect 53576 490 53604 598
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 462 53604 490
rect 53760 480 53788 598
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 56796 490 56824 16546
rect 57072 598 57284 626
rect 57072 490 57100 598
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 462 57100 490
rect 57256 480 57284 598
rect 58452 480 58480 16546
rect 59648 480 59676 16546
rect 60844 480 60872 16546
rect 61568 11756 61620 11762
rect 61568 11698 61620 11704
rect 61580 490 61608 11698
rect 63224 3460 63276 3466
rect 63224 3402 63276 3408
rect 61856 598 62068 626
rect 61856 490 61884 598
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 462 61884 490
rect 62040 480 62068 598
rect 63236 480 63264 3402
rect 64340 480 64368 16546
rect 65076 490 65104 16546
rect 65352 598 65564 626
rect 65352 490 65380 598
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 462 65380 490
rect 65536 480 65564 598
rect 66732 480 66760 16546
rect 67652 6914 67680 28222
rect 67744 7614 67772 128959
rect 67836 127673 67864 156606
rect 68664 156058 68692 156606
rect 68652 156052 68704 156058
rect 68652 155994 68704 156000
rect 67914 143848 67970 143857
rect 67914 143783 67970 143792
rect 67822 127664 67878 127673
rect 67822 127599 67878 127608
rect 67928 125225 67956 143783
rect 69124 143449 69152 219406
rect 70398 155952 70454 155961
rect 70398 155887 70454 155896
rect 70412 154873 70440 155887
rect 70398 154864 70454 154873
rect 70398 154799 70454 154808
rect 70308 149728 70360 149734
rect 70308 149670 70360 149676
rect 69110 143440 69166 143449
rect 69110 143375 69166 143384
rect 69018 143032 69074 143041
rect 69018 142967 69074 142976
rect 69032 134994 69060 142967
rect 70214 139632 70270 139641
rect 70214 139567 70270 139576
rect 69204 137284 69256 137290
rect 69204 137226 69256 137232
rect 68986 134966 69060 134994
rect 68986 134708 69014 134966
rect 69216 134722 69244 137226
rect 70228 134722 70256 139567
rect 70320 135153 70348 149670
rect 70306 135144 70362 135153
rect 70306 135079 70362 135088
rect 70308 135040 70360 135046
rect 70306 135008 70308 135017
rect 70360 135008 70362 135017
rect 70306 134943 70362 134952
rect 69216 134694 69552 134722
rect 70104 134694 70256 134722
rect 70412 134722 70440 154799
rect 70504 140894 70532 239974
rect 72804 239873 72832 241590
rect 72896 241590 73048 241618
rect 73540 241590 73600 241618
rect 73816 241590 74152 241618
rect 74704 241590 74856 241618
rect 74920 241590 75256 241618
rect 75472 241590 75808 241618
rect 76576 241590 76912 241618
rect 72790 239864 72846 239873
rect 72790 239799 72846 239808
rect 72896 239465 72924 241590
rect 73540 241398 73568 241590
rect 73528 241392 73580 241398
rect 73528 241334 73580 241340
rect 73540 240009 73568 241334
rect 73526 240000 73582 240009
rect 73526 239935 73582 239944
rect 72882 239456 72938 239465
rect 71044 239420 71096 239426
rect 72882 239391 72938 239400
rect 71044 239362 71096 239368
rect 71056 155961 71084 239362
rect 73816 238754 73844 241590
rect 74540 240168 74592 240174
rect 74446 240136 74502 240145
rect 74540 240110 74592 240116
rect 74446 240071 74502 240080
rect 73172 238726 73844 238754
rect 71780 234048 71832 234054
rect 71778 234016 71780 234025
rect 71832 234016 71834 234025
rect 71778 233951 71834 233960
rect 71792 188358 71820 233951
rect 71780 188352 71832 188358
rect 71780 188294 71832 188300
rect 73172 184278 73200 238726
rect 74460 236706 74488 240071
rect 74448 236700 74500 236706
rect 74448 236642 74500 236648
rect 74552 217190 74580 240110
rect 74736 238754 74764 241590
rect 74920 240174 74948 241590
rect 74908 240168 74960 240174
rect 75472 240145 75500 241590
rect 74908 240110 74960 240116
rect 75458 240136 75514 240145
rect 75458 240071 75514 240080
rect 76576 238921 76604 241590
rect 76562 238912 76618 238921
rect 76562 238847 76618 238856
rect 74644 238726 74764 238754
rect 74540 217184 74592 217190
rect 74540 217126 74592 217132
rect 73160 184272 73212 184278
rect 73160 184214 73212 184220
rect 73344 168428 73396 168434
rect 73344 168370 73396 168376
rect 73068 161492 73120 161498
rect 73068 161434 73120 161440
rect 72422 157448 72478 157457
rect 72422 157383 72478 157392
rect 71042 155952 71098 155961
rect 71042 155887 71098 155896
rect 71780 145580 71832 145586
rect 71780 145522 71832 145528
rect 70492 140888 70544 140894
rect 70492 140830 70544 140836
rect 71412 140072 71464 140078
rect 71412 140014 71464 140020
rect 71318 138272 71374 138281
rect 71318 138207 71374 138216
rect 71332 134722 71360 138207
rect 70412 134694 70656 134722
rect 71024 134694 71360 134722
rect 71424 134722 71452 140014
rect 71792 134722 71820 145522
rect 72332 138712 72384 138718
rect 72332 138654 72384 138660
rect 72344 134722 72372 138654
rect 72436 135046 72464 157383
rect 73080 137986 73108 161434
rect 73356 151814 73384 168370
rect 73356 151786 73752 151814
rect 73618 139360 73674 139369
rect 73618 139295 73674 139304
rect 73080 137970 73200 137986
rect 73068 137964 73200 137970
rect 73120 137958 73200 137964
rect 73068 137906 73120 137912
rect 73080 137875 73108 137906
rect 72424 135040 72476 135046
rect 73172 135028 73200 137958
rect 73632 135028 73660 139295
rect 73172 135000 73246 135028
rect 72424 134982 72476 134988
rect 71424 134694 71576 134722
rect 71792 134694 72128 134722
rect 72344 134694 72680 134722
rect 73218 134708 73246 135000
rect 73586 135000 73660 135028
rect 73586 134708 73614 135000
rect 73724 134722 73752 151786
rect 74644 142154 74672 238726
rect 77312 238649 77340 241726
rect 77666 241703 77722 241712
rect 78402 241768 78458 241777
rect 79874 241768 79930 241777
rect 78458 241726 78568 241754
rect 79672 241726 79874 241754
rect 78402 241703 78458 241712
rect 81990 241768 82046 241777
rect 79930 241726 80008 241754
rect 79874 241703 79930 241712
rect 77588 241590 78016 241618
rect 77298 238640 77354 238649
rect 77298 238575 77354 238584
rect 77300 236700 77352 236706
rect 77300 236642 77352 236648
rect 75920 229764 75972 229770
rect 75920 229706 75972 229712
rect 75932 229158 75960 229706
rect 75920 229152 75972 229158
rect 75920 229094 75972 229100
rect 75932 229066 76052 229094
rect 75644 217184 75696 217190
rect 75644 217126 75696 217132
rect 75656 216714 75684 217126
rect 75644 216708 75696 216714
rect 75644 216650 75696 216656
rect 74722 149696 74778 149705
rect 74722 149631 74778 149640
rect 74552 142126 74672 142154
rect 74552 140026 74580 142126
rect 74460 139998 74580 140026
rect 74460 134881 74488 139998
rect 74736 135028 74764 149631
rect 75552 136740 75604 136746
rect 75552 136682 75604 136688
rect 74690 135000 74764 135028
rect 74446 134872 74502 134881
rect 74446 134807 74502 134816
rect 73724 134694 74152 134722
rect 74690 134708 74718 135000
rect 75564 134722 75592 136682
rect 75656 134745 75684 216650
rect 75918 176216 75974 176225
rect 75918 176151 75974 176160
rect 75828 140072 75880 140078
rect 75828 140014 75880 140020
rect 75840 138014 75868 140014
rect 75932 138106 75960 176151
rect 76024 140146 76052 229066
rect 76288 141432 76340 141438
rect 76288 141374 76340 141380
rect 76012 140140 76064 140146
rect 76012 140082 76064 140088
rect 75920 138100 75972 138106
rect 75920 138042 75972 138048
rect 75748 137986 75868 138014
rect 75748 134858 75776 137986
rect 75748 134830 75822 134858
rect 75256 134694 75592 134722
rect 75642 134736 75698 134745
rect 75794 134722 75822 134830
rect 76300 134722 76328 141374
rect 76380 138100 76432 138106
rect 76380 138042 76432 138048
rect 75794 134708 75960 134722
rect 75808 134694 75960 134708
rect 76176 134694 76328 134722
rect 76392 134722 76420 138042
rect 77312 135028 77340 236642
rect 77588 236609 77616 241590
rect 78416 240145 78444 241703
rect 78692 241590 79120 241618
rect 77666 240136 77722 240145
rect 77666 240071 77722 240080
rect 78402 240136 78458 240145
rect 78402 240071 78458 240080
rect 77574 236600 77630 236609
rect 77574 236535 77630 236544
rect 77680 236230 77708 240071
rect 78692 238754 78720 241590
rect 78600 238726 78720 238754
rect 77668 236224 77720 236230
rect 77668 236166 77720 236172
rect 78600 227050 78628 238726
rect 79980 231198 80008 241726
rect 81452 241726 81990 241754
rect 80164 241590 80224 241618
rect 80348 241590 80776 241618
rect 80992 241590 81328 241618
rect 80060 239828 80112 239834
rect 80060 239770 80112 239776
rect 79968 231192 80020 231198
rect 79968 231134 80020 231140
rect 79324 231124 79376 231130
rect 79324 231066 79376 231072
rect 78588 227044 78640 227050
rect 78588 226986 78640 226992
rect 79336 184958 79364 231066
rect 80072 228410 80100 239770
rect 80164 238513 80192 241590
rect 80150 238504 80206 238513
rect 80150 238439 80206 238448
rect 80164 237969 80192 238439
rect 80150 237960 80206 237969
rect 80150 237895 80206 237904
rect 80348 233238 80376 241590
rect 80992 239834 81020 241590
rect 80980 239828 81032 239834
rect 80980 239770 81032 239776
rect 81452 238754 81480 241726
rect 83738 241768 83794 241777
rect 83536 241740 83738 241754
rect 81990 241703 82046 241712
rect 83522 241726 83738 241740
rect 83522 241618 83550 241726
rect 85946 241768 86002 241777
rect 85744 241726 85946 241754
rect 83738 241703 83794 241712
rect 85946 241703 86002 241712
rect 86590 241768 86646 241777
rect 91558 241768 91614 241777
rect 86646 241740 86848 241754
rect 86646 241726 86862 241740
rect 86590 241703 86646 241712
rect 86834 241618 86862 241726
rect 91614 241726 91816 241754
rect 91558 241703 91614 241712
rect 90270 241632 90326 241641
rect 81360 238726 81480 238754
rect 82096 241590 82432 241618
rect 82924 241590 82984 241618
rect 83476 241604 83550 241618
rect 83476 241590 83536 241604
rect 83752 241590 84088 241618
rect 84304 241590 84640 241618
rect 84856 241590 85192 241618
rect 85868 241590 86296 241618
rect 86834 241604 86908 241618
rect 86848 241590 86908 241604
rect 80336 233232 80388 233238
rect 80336 233174 80388 233180
rect 80060 228404 80112 228410
rect 80060 228346 80112 228352
rect 80704 189780 80756 189786
rect 80704 189722 80756 189728
rect 79324 184952 79376 184958
rect 79324 184894 79376 184900
rect 77942 164384 77998 164393
rect 77942 164319 77998 164328
rect 77956 149734 77984 164319
rect 77944 149728 77996 149734
rect 77944 149670 77996 149676
rect 78680 144424 78732 144430
rect 78680 144366 78732 144372
rect 78036 138780 78088 138786
rect 78036 138722 78088 138728
rect 77266 135000 77340 135028
rect 76392 134694 76728 134722
rect 77266 134708 77294 135000
rect 78048 134722 78076 138722
rect 78496 136672 78548 136678
rect 78496 136614 78548 136620
rect 78508 134722 78536 136614
rect 78692 135028 78720 144366
rect 78772 136740 78824 136746
rect 78772 136682 78824 136688
rect 78784 136649 78812 136682
rect 79336 136678 79364 184894
rect 80060 151156 80112 151162
rect 80060 151098 80112 151104
rect 80072 147674 80100 151098
rect 80716 148374 80744 189722
rect 81360 188358 81388 238726
rect 82096 234598 82124 241590
rect 82820 240168 82872 240174
rect 82820 240110 82872 240116
rect 82084 234592 82136 234598
rect 82084 234534 82136 234540
rect 81348 188352 81400 188358
rect 81348 188294 81400 188300
rect 81992 149796 82044 149802
rect 81992 149738 82044 149744
rect 80704 148368 80756 148374
rect 80704 148310 80756 148316
rect 80072 147646 81020 147674
rect 80520 146328 80572 146334
rect 80520 146270 80572 146276
rect 79966 141400 80022 141409
rect 79966 141335 80022 141344
rect 79598 137320 79654 137329
rect 79598 137255 79600 137264
rect 79652 137255 79654 137264
rect 79600 137226 79652 137232
rect 79324 136672 79376 136678
rect 78770 136640 78826 136649
rect 79324 136614 79376 136620
rect 78770 136575 78826 136584
rect 78692 135000 78766 135028
rect 77832 134694 78076 134722
rect 78200 134694 78536 134722
rect 78738 134708 78766 135000
rect 79612 134722 79640 137226
rect 79980 134722 80008 141335
rect 80428 140752 80480 140758
rect 80428 140694 80480 140700
rect 80440 134994 80468 140694
rect 79304 134694 79640 134722
rect 79856 134694 80008 134722
rect 80394 134966 80468 134994
rect 80394 134708 80422 134966
rect 80532 134722 80560 146270
rect 80992 134722 81020 147646
rect 81900 138712 81952 138718
rect 81900 138654 81952 138660
rect 81912 134994 81940 138654
rect 81866 134966 81940 134994
rect 80532 134694 80776 134722
rect 80992 134694 81328 134722
rect 81866 134708 81894 134966
rect 82004 134722 82032 149738
rect 82096 140865 82124 234534
rect 82832 218754 82860 240110
rect 82924 238377 82952 241590
rect 82910 238368 82966 238377
rect 82910 238303 82966 238312
rect 82820 218748 82872 218754
rect 82820 218690 82872 218696
rect 82174 176760 82230 176769
rect 82174 176695 82230 176704
rect 82188 144430 82216 176695
rect 83476 164898 83504 241590
rect 83752 240174 83780 241590
rect 83740 240168 83792 240174
rect 83740 240110 83792 240116
rect 84200 240168 84252 240174
rect 84200 240110 84252 240116
rect 83556 236224 83608 236230
rect 83556 236166 83608 236172
rect 83568 220153 83596 236166
rect 84212 231130 84240 240110
rect 84304 238649 84332 241590
rect 84856 240174 84884 241590
rect 84844 240168 84896 240174
rect 84844 240110 84896 240116
rect 85868 238754 85896 241590
rect 85592 238726 85896 238754
rect 84290 238640 84346 238649
rect 84290 238575 84346 238584
rect 84200 231124 84252 231130
rect 84200 231066 84252 231072
rect 83554 220144 83610 220153
rect 83554 220079 83610 220088
rect 85592 211857 85620 238726
rect 85578 211848 85634 211857
rect 85578 211783 85634 211792
rect 86880 181558 86908 241590
rect 87064 241590 87400 241618
rect 87616 241590 87952 241618
rect 88352 241590 88504 241618
rect 89056 241590 89392 241618
rect 89608 241590 89668 241618
rect 90160 241590 90270 241618
rect 86960 240168 87012 240174
rect 86960 240110 87012 240116
rect 86972 215966 87000 240110
rect 87064 222154 87092 241590
rect 87616 240174 87644 241590
rect 87604 240168 87656 240174
rect 87604 240110 87656 240116
rect 88352 232558 88380 241590
rect 88430 240136 88486 240145
rect 88430 240071 88486 240080
rect 88340 232552 88392 232558
rect 88340 232494 88392 232500
rect 87604 231192 87656 231198
rect 87604 231134 87656 231140
rect 87052 222148 87104 222154
rect 87052 222090 87104 222096
rect 86960 215960 87012 215966
rect 86960 215902 87012 215908
rect 86868 181552 86920 181558
rect 86868 181494 86920 181500
rect 87616 178702 87644 231134
rect 88248 215960 88300 215966
rect 88248 215902 88300 215908
rect 87604 178696 87656 178702
rect 87604 178638 87656 178644
rect 83554 177304 83610 177313
rect 83554 177239 83610 177248
rect 83464 164892 83516 164898
rect 83464 164834 83516 164840
rect 82912 163600 82964 163606
rect 82912 163542 82964 163548
rect 82820 149524 82872 149530
rect 82820 149466 82872 149472
rect 82176 144424 82228 144430
rect 82176 144366 82228 144372
rect 82082 140856 82138 140865
rect 82082 140791 82138 140800
rect 82832 134994 82860 149466
rect 82924 142866 82952 163542
rect 83002 156088 83058 156097
rect 83002 156023 83058 156032
rect 82912 142860 82964 142866
rect 82912 142802 82964 142808
rect 82786 134966 82860 134994
rect 82004 134694 82432 134722
rect 82786 134708 82814 134966
rect 83016 134722 83044 156023
rect 83568 147674 83596 177239
rect 87144 172576 87196 172582
rect 87144 172518 87196 172524
rect 86314 172408 86370 172417
rect 86314 172343 86370 172352
rect 86328 171193 86356 172343
rect 86314 171184 86370 171193
rect 86314 171119 86370 171128
rect 86224 169788 86276 169794
rect 86224 169730 86276 169736
rect 83476 147646 83596 147674
rect 83476 140758 83504 147646
rect 86130 143576 86186 143585
rect 86130 143511 86186 143520
rect 83556 142860 83608 142866
rect 83556 142802 83608 142808
rect 83464 140752 83516 140758
rect 83464 140694 83516 140700
rect 83568 134722 83596 142802
rect 84842 142080 84898 142089
rect 84842 142015 84898 142024
rect 84750 140040 84806 140049
rect 84750 139975 84806 139984
rect 84764 134722 84792 139975
rect 83016 134694 83352 134722
rect 83568 134694 83904 134722
rect 84456 134694 84792 134722
rect 84856 134722 84884 142015
rect 86144 137970 86172 143511
rect 86132 137964 86184 137970
rect 86132 137906 86184 137912
rect 85488 136672 85540 136678
rect 85488 136614 85540 136620
rect 85500 134722 85528 136614
rect 86144 134722 86172 137906
rect 86236 136678 86264 169730
rect 86328 149530 86356 171119
rect 86958 164520 87014 164529
rect 86958 164455 87014 164464
rect 86868 149728 86920 149734
rect 86868 149670 86920 149676
rect 86316 149524 86368 149530
rect 86316 149466 86368 149472
rect 86880 146266 86908 149670
rect 86868 146260 86920 146266
rect 86868 146202 86920 146208
rect 86880 144974 86908 146202
rect 86868 144968 86920 144974
rect 86868 144910 86920 144916
rect 86866 144800 86922 144809
rect 86866 144735 86922 144744
rect 86880 139466 86908 144735
rect 86868 139460 86920 139466
rect 86868 139402 86920 139408
rect 86880 138014 86908 139402
rect 86788 137986 86908 138014
rect 86224 136672 86276 136678
rect 86224 136614 86276 136620
rect 86788 134722 86816 137986
rect 86972 134994 87000 164455
rect 86972 134966 87046 134994
rect 84856 134694 85008 134722
rect 85376 134694 85528 134722
rect 85928 134694 86172 134722
rect 86480 134694 86816 134722
rect 87018 134708 87046 134966
rect 87156 134722 87184 172518
rect 88260 151065 88288 215902
rect 88444 180130 88472 240071
rect 89364 239494 89392 241590
rect 89640 240009 89668 241590
rect 90822 241632 90878 241641
rect 90270 241567 90326 241576
rect 90376 241590 90712 241618
rect 89626 240000 89682 240009
rect 89626 239935 89682 239944
rect 89352 239488 89404 239494
rect 89352 239430 89404 239436
rect 90376 238754 90404 241590
rect 90822 241567 90878 241576
rect 91204 241590 91264 241618
rect 92032 241590 92368 241618
rect 92584 241590 92920 241618
rect 89732 238726 90404 238754
rect 89628 236496 89680 236502
rect 89628 236438 89680 236444
rect 89640 184210 89668 236438
rect 89732 231198 89760 238726
rect 89720 231192 89772 231198
rect 89720 231134 89772 231140
rect 89628 184204 89680 184210
rect 89628 184146 89680 184152
rect 88432 180124 88484 180130
rect 88432 180066 88484 180072
rect 88340 174548 88392 174554
rect 88340 174490 88392 174496
rect 88246 151056 88302 151065
rect 88246 150991 88302 151000
rect 87696 144968 87748 144974
rect 87696 144910 87748 144916
rect 87708 134722 87736 144910
rect 88352 134722 88380 174490
rect 89718 167104 89774 167113
rect 89718 167039 89774 167048
rect 88984 163532 89036 163538
rect 88984 163474 89036 163480
rect 88996 149705 89024 163474
rect 88982 149696 89038 149705
rect 88982 149631 89038 149640
rect 89166 147792 89222 147801
rect 89166 147727 89222 147736
rect 88432 142316 88484 142322
rect 88432 142258 88484 142264
rect 88444 142089 88472 142258
rect 88430 142080 88486 142089
rect 88430 142015 88486 142024
rect 89074 137320 89130 137329
rect 89074 137255 89130 137264
rect 89088 134858 89116 137255
rect 89042 134830 89116 134858
rect 87156 134694 87584 134722
rect 87708 134694 87952 134722
rect 88352 134694 88504 134722
rect 89042 134708 89070 134830
rect 89180 134722 89208 147727
rect 89732 134722 89760 167039
rect 90364 165640 90416 165646
rect 90364 165582 90416 165588
rect 90376 151162 90404 165582
rect 90364 151156 90416 151162
rect 90364 151098 90416 151104
rect 90836 144809 90864 241567
rect 91098 240136 91154 240145
rect 91098 240071 91154 240080
rect 91112 236502 91140 240071
rect 91100 236496 91152 236502
rect 91100 236438 91152 236444
rect 91100 236360 91152 236366
rect 91100 236302 91152 236308
rect 91112 236065 91140 236302
rect 91098 236056 91154 236065
rect 91204 236026 91232 241590
rect 91928 239488 91980 239494
rect 91926 239456 91928 239465
rect 91980 239456 91982 239465
rect 91926 239391 91982 239400
rect 92032 238754 92060 241590
rect 91388 238726 92060 238754
rect 91098 235991 91154 236000
rect 91192 236020 91244 236026
rect 91192 235962 91244 235968
rect 91388 224330 91416 238726
rect 92584 237386 92612 241590
rect 93458 241466 93486 241604
rect 93872 241590 94024 241618
rect 94148 241590 94576 241618
rect 95128 241590 95188 241618
rect 93124 241460 93176 241466
rect 93124 241402 93176 241408
rect 93446 241460 93498 241466
rect 93446 241402 93498 241408
rect 92572 237380 92624 237386
rect 92572 237322 92624 237328
rect 92386 236464 92442 236473
rect 92386 236399 92442 236408
rect 91376 224324 91428 224330
rect 91376 224266 91428 224272
rect 91744 184272 91796 184278
rect 91744 184214 91796 184220
rect 91192 170400 91244 170406
rect 91192 170342 91244 170348
rect 91204 151814 91232 170342
rect 91204 151786 91692 151814
rect 91008 148368 91060 148374
rect 91008 148310 91060 148316
rect 90822 144800 90878 144809
rect 90822 144735 90878 144744
rect 90822 140856 90878 140865
rect 90822 140791 90878 140800
rect 90836 134722 90864 140791
rect 91020 138014 91048 148310
rect 91020 137986 91140 138014
rect 91006 136912 91062 136921
rect 91006 136847 91062 136856
rect 91020 135930 91048 136847
rect 91112 135969 91140 137986
rect 91098 135960 91154 135969
rect 91008 135924 91060 135930
rect 91098 135895 91154 135904
rect 91282 135960 91338 135969
rect 91282 135895 91338 135904
rect 91008 135866 91060 135872
rect 91192 135584 91244 135590
rect 91192 135526 91244 135532
rect 91204 135318 91232 135526
rect 91192 135312 91244 135318
rect 91192 135254 91244 135260
rect 89180 134694 89608 134722
rect 89732 134694 89976 134722
rect 90528 134694 90864 134722
rect 75642 134671 75698 134680
rect 75932 134638 75960 134694
rect 75920 134632 75972 134638
rect 91204 134586 91232 135254
rect 91296 134722 91324 135895
rect 91664 134858 91692 151786
rect 91756 136202 91784 184214
rect 92400 158778 92428 236399
rect 93136 213926 93164 241402
rect 93124 213920 93176 213926
rect 93124 213862 93176 213868
rect 93872 206378 93900 241590
rect 94148 234161 94176 241590
rect 95160 240038 95188 241590
rect 95252 241604 95680 241618
rect 95252 241590 95694 241604
rect 95148 240032 95200 240038
rect 95148 239974 95200 239980
rect 94778 237280 94834 237289
rect 94778 237215 94834 237224
rect 94792 236366 94820 237215
rect 94780 236360 94832 236366
rect 94780 236302 94832 236308
rect 95252 236026 95280 241590
rect 95666 241466 95694 241590
rect 95896 241590 96232 241618
rect 96632 241590 96784 241618
rect 96908 241590 97336 241618
rect 97552 241590 97888 241618
rect 95654 241460 95706 241466
rect 95654 241402 95706 241408
rect 95896 238754 95924 241590
rect 95344 238726 95924 238754
rect 94688 236020 94740 236026
rect 94688 235962 94740 235968
rect 95240 236020 95292 236026
rect 95240 235962 95292 235968
rect 94134 234152 94190 234161
rect 94134 234087 94190 234096
rect 93860 206372 93912 206378
rect 93860 206314 93912 206320
rect 92664 171148 92716 171154
rect 92664 171090 92716 171096
rect 91836 158772 91888 158778
rect 91836 158714 91888 158720
rect 92388 158772 92440 158778
rect 92388 158714 92440 158720
rect 91744 136196 91796 136202
rect 91744 136138 91796 136144
rect 91848 135590 91876 158714
rect 91928 154624 91980 154630
rect 91928 154566 91980 154572
rect 91940 140078 91968 154566
rect 92478 145616 92534 145625
rect 92478 145551 92534 145560
rect 91928 140072 91980 140078
rect 91928 140014 91980 140020
rect 91836 135584 91888 135590
rect 91836 135526 91888 135532
rect 92492 134994 92520 145551
rect 92492 134966 92566 134994
rect 91664 134830 91784 134858
rect 91756 134722 91784 134830
rect 91296 134694 91632 134722
rect 91756 134694 92184 134722
rect 92538 134708 92566 134966
rect 92676 134722 92704 171090
rect 92756 152584 92808 152590
rect 92756 152526 92808 152532
rect 92768 151814 92796 152526
rect 92768 151786 93256 151814
rect 93228 134722 93256 151786
rect 94320 145648 94372 145654
rect 94320 145590 94372 145596
rect 94332 134722 94360 145590
rect 92676 134694 93104 134722
rect 93228 134694 93656 134722
rect 94332 134694 94576 134722
rect 94412 134632 94464 134638
rect 75920 134574 75972 134580
rect 91080 134558 91232 134586
rect 94208 134580 94412 134586
rect 94208 134574 94464 134580
rect 94208 134558 94452 134574
rect 94700 133226 94728 235962
rect 95240 212560 95292 212566
rect 95240 212502 95292 212508
rect 94870 138136 94926 138145
rect 94870 138071 94926 138080
rect 94884 138014 94912 138071
rect 94884 137986 95004 138014
rect 94700 133198 94912 133226
rect 94780 129736 94832 129742
rect 94780 129678 94832 129684
rect 94792 127786 94820 129678
rect 94608 127758 94820 127786
rect 67914 125216 67970 125225
rect 67914 125151 67970 125160
rect 67822 101008 67878 101017
rect 67822 100943 67878 100952
rect 67836 92041 67864 100943
rect 68558 95840 68614 95849
rect 68558 95775 68614 95784
rect 68572 93854 68600 95775
rect 69018 94480 69074 94489
rect 69018 94415 69074 94424
rect 68008 93832 68060 93838
rect 68008 93774 68060 93780
rect 68388 93826 68600 93854
rect 68020 93401 68048 93774
rect 68006 93392 68062 93401
rect 68006 93327 68062 93336
rect 67822 92032 67878 92041
rect 67822 91967 67878 91976
rect 68020 60625 68048 93327
rect 68388 89593 68416 93826
rect 69032 92954 69060 94415
rect 69020 92948 69072 92954
rect 69020 92890 69072 92896
rect 68468 92880 68520 92886
rect 68520 92828 68968 92834
rect 68468 92822 68968 92828
rect 68480 92806 68968 92822
rect 68940 90302 68968 92806
rect 69032 92806 69184 92834
rect 68928 90296 68980 90302
rect 68928 90238 68980 90244
rect 68374 89584 68430 89593
rect 68374 89519 68430 89528
rect 69032 84182 69060 92806
rect 69722 92698 69750 92820
rect 70274 92750 70302 92820
rect 70262 92744 70314 92750
rect 69722 92670 69888 92698
rect 70262 92686 70314 92692
rect 69860 91089 69888 92670
rect 70274 92562 70302 92686
rect 70826 92562 70854 92820
rect 71194 92698 71222 92820
rect 71148 92670 71222 92698
rect 71746 92698 71774 92820
rect 71746 92670 71820 92698
rect 70274 92534 70348 92562
rect 70826 92534 70900 92562
rect 69846 91080 69902 91089
rect 69846 91015 69902 91024
rect 69860 85377 69888 91015
rect 69846 85368 69902 85377
rect 69846 85303 69902 85312
rect 69020 84176 69072 84182
rect 69020 84118 69072 84124
rect 69018 82104 69074 82113
rect 69018 82039 69074 82048
rect 68006 60616 68062 60625
rect 68006 60551 68062 60560
rect 69032 16574 69060 82039
rect 70320 76566 70348 92534
rect 70872 86601 70900 92534
rect 71148 91050 71176 92670
rect 71792 92449 71820 92670
rect 72298 92562 72326 92820
rect 72850 92562 72878 92820
rect 73402 92698 73430 92820
rect 71884 92534 72326 92562
rect 72804 92534 72878 92562
rect 73356 92670 73430 92698
rect 71778 92440 71834 92449
rect 71778 92375 71834 92384
rect 71136 91044 71188 91050
rect 71136 90986 71188 90992
rect 71044 90296 71096 90302
rect 71044 90238 71096 90244
rect 70858 86592 70914 86601
rect 70858 86527 70914 86536
rect 70308 76560 70360 76566
rect 70308 76502 70360 76508
rect 70398 76528 70454 76537
rect 70398 76463 70454 76472
rect 70412 16574 70440 76463
rect 71056 63510 71084 90238
rect 71792 87961 71820 92375
rect 71778 87952 71834 87961
rect 71778 87887 71834 87896
rect 71884 81326 71912 92534
rect 72804 92410 72832 92534
rect 73356 92449 73384 92670
rect 73770 92562 73798 92820
rect 74322 92721 74350 92820
rect 74874 92721 74902 92820
rect 74308 92712 74364 92721
rect 74308 92647 74364 92656
rect 74860 92712 74916 92721
rect 75426 92698 75454 92820
rect 74860 92647 74916 92656
rect 75380 92670 75592 92698
rect 74322 92562 74350 92647
rect 74632 92608 74684 92614
rect 73770 92534 73844 92562
rect 74322 92534 74396 92562
rect 75380 92585 75408 92670
rect 74632 92550 74684 92556
rect 75366 92576 75422 92585
rect 73342 92440 73398 92449
rect 72792 92404 72844 92410
rect 73342 92375 73398 92384
rect 72792 92346 72844 92352
rect 73816 86902 73844 92534
rect 73804 86896 73856 86902
rect 73804 86838 73856 86844
rect 74368 84194 74396 92534
rect 74368 84166 74488 84194
rect 71872 81320 71924 81326
rect 71872 81262 71924 81268
rect 74460 71777 74488 84166
rect 74540 75200 74592 75206
rect 74540 75142 74592 75148
rect 74446 71768 74502 71777
rect 74446 71703 74502 71712
rect 71044 63504 71096 63510
rect 71044 63446 71096 63452
rect 71780 49020 71832 49026
rect 71780 48962 71832 48968
rect 71792 16574 71820 48962
rect 74552 16574 74580 75142
rect 74644 67590 74672 92550
rect 75366 92511 75422 92520
rect 75564 84194 75592 92670
rect 75794 92614 75822 92820
rect 75782 92608 75834 92614
rect 76346 92562 76374 92820
rect 76898 92721 76926 92820
rect 76884 92712 76940 92721
rect 76884 92647 76940 92656
rect 75782 92550 75834 92556
rect 76300 92534 76374 92562
rect 76898 92562 76926 92647
rect 77450 92562 77478 92820
rect 76898 92534 76972 92562
rect 76300 92313 76328 92534
rect 76286 92304 76342 92313
rect 76286 92239 76342 92248
rect 76944 84194 76972 92534
rect 77312 92534 77478 92562
rect 78002 92562 78030 92820
rect 78370 92562 78398 92820
rect 78922 92562 78950 92820
rect 79474 92562 79502 92820
rect 78002 92534 78076 92562
rect 78370 92534 78444 92562
rect 78922 92534 78996 92562
rect 75564 84166 75868 84194
rect 76944 84166 77248 84194
rect 75840 78674 75868 84166
rect 75828 78668 75880 78674
rect 75828 78610 75880 78616
rect 74632 67584 74684 67590
rect 74632 67526 74684 67532
rect 77220 57934 77248 84166
rect 77312 80073 77340 92534
rect 78048 89457 78076 92534
rect 78416 89729 78444 92534
rect 78968 91089 78996 92534
rect 79428 92534 79502 92562
rect 80026 92562 80054 92820
rect 80152 92608 80204 92614
rect 80026 92534 80100 92562
rect 80578 92562 80606 92820
rect 80946 92614 80974 92820
rect 81498 92698 81526 92820
rect 81452 92670 81526 92698
rect 80152 92550 80204 92556
rect 78954 91080 79010 91089
rect 78954 91015 79010 91024
rect 78402 89720 78458 89729
rect 79428 89690 79456 92534
rect 78402 89655 78458 89664
rect 79416 89684 79468 89690
rect 79416 89626 79468 89632
rect 78034 89448 78090 89457
rect 78034 89383 78090 89392
rect 77298 80064 77354 80073
rect 80072 80034 80100 92534
rect 77298 79999 77354 80008
rect 80060 80028 80112 80034
rect 80060 79970 80112 79976
rect 80164 73166 80192 92550
rect 80256 92534 80606 92562
rect 80934 92608 80986 92614
rect 80934 92550 80986 92556
rect 80256 82754 80284 92534
rect 81452 92449 81480 92670
rect 82050 92562 82078 92820
rect 82602 92698 82630 92820
rect 82602 92670 82676 92698
rect 82050 92534 82124 92562
rect 81438 92440 81494 92449
rect 81438 92375 81494 92384
rect 82096 88097 82124 92534
rect 82648 88262 82676 92670
rect 82970 92562 82998 92820
rect 83522 92562 83550 92820
rect 84074 92562 84102 92820
rect 84626 92562 84654 92820
rect 85178 92562 85206 92820
rect 85546 92562 85574 92820
rect 86098 92562 86126 92820
rect 82970 92534 83044 92562
rect 83522 92534 83596 92562
rect 84074 92534 84148 92562
rect 84626 92534 84700 92562
rect 85178 92534 85252 92562
rect 85546 92534 85620 92562
rect 82636 88256 82688 88262
rect 82636 88198 82688 88204
rect 82082 88088 82138 88097
rect 82082 88023 82138 88032
rect 83016 86873 83044 92534
rect 83568 92449 83596 92534
rect 83554 92440 83610 92449
rect 83554 92375 83610 92384
rect 84120 89622 84148 92534
rect 84672 91050 84700 92534
rect 84660 91044 84712 91050
rect 84660 90986 84712 90992
rect 85224 90370 85252 92534
rect 85212 90364 85264 90370
rect 85212 90306 85264 90312
rect 85592 89690 85620 92534
rect 85684 92534 86126 92562
rect 86650 92562 86678 92820
rect 87202 92698 87230 92820
rect 87202 92670 87276 92698
rect 86650 92534 86724 92562
rect 85580 89684 85632 89690
rect 85580 89626 85632 89632
rect 84108 89616 84160 89622
rect 84108 89558 84160 89564
rect 83464 88256 83516 88262
rect 83464 88198 83516 88204
rect 83002 86864 83058 86873
rect 83002 86799 83058 86808
rect 80244 82748 80296 82754
rect 80244 82690 80296 82696
rect 80152 73160 80204 73166
rect 80152 73102 80204 73108
rect 77208 57928 77260 57934
rect 77208 57870 77260 57876
rect 83476 56574 83504 88198
rect 85684 84017 85712 92534
rect 86696 88262 86724 92534
rect 86684 88256 86736 88262
rect 86684 88198 86736 88204
rect 87248 85542 87276 92670
rect 87570 92562 87598 92820
rect 88122 92562 88150 92820
rect 88674 92682 88702 92820
rect 88662 92676 88714 92682
rect 88662 92618 88714 92624
rect 89226 92562 89254 92820
rect 89626 92712 89682 92721
rect 89626 92647 89628 92656
rect 89680 92647 89682 92656
rect 89628 92618 89680 92624
rect 87340 92534 87598 92562
rect 87800 92534 88150 92562
rect 88352 92534 89254 92562
rect 87236 85536 87288 85542
rect 87236 85478 87288 85484
rect 87340 85354 87368 92534
rect 86972 85326 87368 85354
rect 85670 84008 85726 84017
rect 85670 83943 85726 83952
rect 85580 73840 85632 73846
rect 85580 73782 85632 73788
rect 83464 56568 83516 56574
rect 83464 56510 83516 56516
rect 75184 51808 75236 51814
rect 75184 51750 75236 51756
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 67732 7608 67784 7614
rect 67732 7550 67784 7556
rect 67652 6886 67956 6914
rect 67928 480 67956 6886
rect 69112 4820 69164 4826
rect 69112 4762 69164 4768
rect 69124 480 69152 4762
rect 69860 490 69888 16546
rect 70136 598 70348 626
rect 70136 490 70164 598
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69860 462 70164 490
rect 70320 480 70348 598
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 73344 10396 73396 10402
rect 73344 10338 73396 10344
rect 73356 490 73384 10338
rect 73632 598 73844 626
rect 73632 490 73660 598
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 462 73660 490
rect 73816 480 73844 598
rect 75012 480 75040 16546
rect 75196 3466 75224 51750
rect 75920 39364 75972 39370
rect 75920 39306 75972 39312
rect 75932 16574 75960 39306
rect 81440 29640 81492 29646
rect 81440 29582 81492 29588
rect 78680 22772 78732 22778
rect 78680 22714 78732 22720
rect 78692 16574 78720 22714
rect 81452 16574 81480 29582
rect 82820 26920 82872 26926
rect 82820 26862 82872 26868
rect 82832 16574 82860 26862
rect 85592 16574 85620 73782
rect 86972 63442 87000 85326
rect 87800 84194 87828 92534
rect 87064 84166 87828 84194
rect 87064 66230 87092 84166
rect 88352 82822 88380 92534
rect 88340 82816 88392 82822
rect 88340 82758 88392 82764
rect 88340 72480 88392 72486
rect 88340 72422 88392 72428
rect 87052 66224 87104 66230
rect 87052 66166 87104 66172
rect 86960 63436 87012 63442
rect 86960 63378 87012 63384
rect 87604 53100 87656 53106
rect 87604 53042 87656 53048
rect 75932 16546 76236 16574
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 85592 16546 85712 16574
rect 75184 3460 75236 3466
rect 75184 3402 75236 3408
rect 76208 480 76236 16546
rect 78588 8968 78640 8974
rect 78588 8910 78640 8916
rect 77392 3460 77444 3466
rect 77392 3402 77444 3408
rect 77404 480 77432 3402
rect 78600 480 78628 8910
rect 79244 490 79272 16546
rect 80888 6180 80940 6186
rect 80888 6122 80940 6128
rect 79520 598 79732 626
rect 79520 490 79548 598
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 462 79548 490
rect 79704 480 79732 598
rect 80900 480 80928 6122
rect 81636 490 81664 16546
rect 81912 598 82124 626
rect 81912 490 81940 598
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 462 81940 490
rect 82096 480 82124 598
rect 83292 480 83320 16546
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 84488 480 84516 3470
rect 85684 480 85712 16546
rect 87512 14476 87564 14482
rect 87512 14418 87564 14424
rect 86408 10328 86460 10334
rect 86408 10270 86460 10276
rect 86420 490 86448 10270
rect 86696 598 86908 626
rect 86696 490 86724 598
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 462 86724 490
rect 86880 480 86908 598
rect 87524 490 87552 14418
rect 87616 9042 87644 53042
rect 88352 16574 88380 72422
rect 89640 60722 89668 92618
rect 89778 92562 89806 92820
rect 90146 92682 90174 92820
rect 90134 92676 90186 92682
rect 90134 92618 90186 92624
rect 90698 92562 90726 92820
rect 91250 92562 91278 92820
rect 91802 92750 91830 92820
rect 91790 92744 91842 92750
rect 91790 92686 91842 92692
rect 92354 92562 92382 92820
rect 92722 92698 92750 92820
rect 92722 92670 92796 92698
rect 89778 92534 89852 92562
rect 89824 86970 89852 92534
rect 89916 92534 90726 92562
rect 91112 92534 91278 92562
rect 91480 92534 92382 92562
rect 89812 86964 89864 86970
rect 89812 86906 89864 86912
rect 89916 75857 89944 92534
rect 90362 84824 90418 84833
rect 90362 84759 90418 84768
rect 89902 75848 89958 75857
rect 89902 75783 89958 75792
rect 89628 60716 89680 60722
rect 89628 60658 89680 60664
rect 90376 20670 90404 84759
rect 91112 81433 91140 92534
rect 91480 83881 91508 92534
rect 92768 92313 92796 92670
rect 93274 92562 93302 92820
rect 92952 92534 93302 92562
rect 93826 92562 93854 92820
rect 94378 92698 94406 92820
rect 94608 92698 94636 127758
rect 94884 127514 94912 133198
rect 94976 129674 95004 137986
rect 95148 134632 95200 134638
rect 95148 134574 95200 134580
rect 95160 134026 95188 134574
rect 95148 134020 95200 134026
rect 95148 133962 95200 133968
rect 94964 129668 95016 129674
rect 94964 129610 95016 129616
rect 94378 92670 94636 92698
rect 94700 127486 94912 127514
rect 94700 92562 94728 127486
rect 95252 92750 95280 212502
rect 95344 206038 95372 238726
rect 96528 227792 96580 227798
rect 96528 227734 96580 227740
rect 95700 213920 95752 213926
rect 95700 213862 95752 213868
rect 95712 212566 95740 213862
rect 95700 212560 95752 212566
rect 95700 212502 95752 212508
rect 95884 206304 95936 206310
rect 95884 206246 95936 206252
rect 95896 206038 95924 206246
rect 95332 206032 95384 206038
rect 95332 205974 95384 205980
rect 95884 206032 95936 206038
rect 95884 205974 95936 205980
rect 95896 129742 95924 205974
rect 95974 164520 96030 164529
rect 95974 164455 96030 164464
rect 95988 164257 96016 164455
rect 95974 164248 96030 164257
rect 95974 164183 96030 164192
rect 95976 136196 96028 136202
rect 95976 136138 96028 136144
rect 95884 129736 95936 129742
rect 95884 129678 95936 129684
rect 95330 120320 95386 120329
rect 95330 120255 95386 120264
rect 95240 92744 95292 92750
rect 95240 92686 95292 92692
rect 93826 92534 94728 92562
rect 92754 92304 92810 92313
rect 92754 92239 92810 92248
rect 92952 84194 92980 92534
rect 94502 90400 94558 90409
rect 94502 90335 94504 90344
rect 94556 90335 94558 90344
rect 94504 90306 94556 90312
rect 92492 84166 92980 84194
rect 91466 83872 91522 83881
rect 91466 83807 91522 83816
rect 91098 81424 91154 81433
rect 91098 81359 91154 81368
rect 92492 77246 92520 84166
rect 92480 77240 92532 77246
rect 92480 77182 92532 77188
rect 92480 71052 92532 71058
rect 92480 70994 92532 71000
rect 90364 20664 90416 20670
rect 90364 20606 90416 20612
rect 92492 16574 92520 70994
rect 93860 68332 93912 68338
rect 93860 68274 93912 68280
rect 93872 16574 93900 68274
rect 94516 59362 94544 90306
rect 94700 69018 94728 92534
rect 95344 71738 95372 120255
rect 95424 95260 95476 95266
rect 95424 95202 95476 95208
rect 95436 89593 95464 95202
rect 95988 95198 96016 136138
rect 96540 103601 96568 227734
rect 96632 204950 96660 241590
rect 96908 238066 96936 241590
rect 97552 238754 97580 241590
rect 98104 238754 98132 247007
rect 98644 245676 98696 245682
rect 98644 245618 98696 245624
rect 98426 241534 98454 241604
rect 98414 241528 98466 241534
rect 98414 241470 98466 241476
rect 97000 238726 97580 238754
rect 98012 238726 98132 238754
rect 96896 238060 96948 238066
rect 96896 238002 96948 238008
rect 97000 229226 97028 238726
rect 97908 233912 97960 233918
rect 97908 233854 97960 233860
rect 96988 229220 97040 229226
rect 96988 229162 97040 229168
rect 97000 229094 97028 229162
rect 97000 229066 97304 229094
rect 97276 207058 97304 229066
rect 97264 207052 97316 207058
rect 97264 206994 97316 207000
rect 96620 204944 96672 204950
rect 96620 204886 96672 204892
rect 97816 195288 97868 195294
rect 97816 195230 97868 195236
rect 97264 156460 97316 156466
rect 97264 156402 97316 156408
rect 96712 133884 96764 133890
rect 96712 133826 96764 133832
rect 96724 133113 96752 133826
rect 96710 133104 96766 133113
rect 96710 133039 96766 133048
rect 96712 132388 96764 132394
rect 96712 132330 96764 132336
rect 96724 132297 96752 132330
rect 96710 132288 96766 132297
rect 96710 132223 96766 132232
rect 96802 130928 96858 130937
rect 96802 130863 96858 130872
rect 96816 130422 96844 130863
rect 96804 130416 96856 130422
rect 96804 130358 96856 130364
rect 96712 130212 96764 130218
rect 96712 130154 96764 130160
rect 96724 130121 96752 130154
rect 96710 130112 96766 130121
rect 96710 130047 96766 130056
rect 96618 125488 96674 125497
rect 96618 125423 96674 125432
rect 96632 124914 96660 125423
rect 96620 124908 96672 124914
rect 96620 124850 96672 124856
rect 96526 103592 96582 103601
rect 96526 103527 96528 103536
rect 96580 103527 96582 103536
rect 96528 103498 96580 103504
rect 95976 95192 96028 95198
rect 95976 95134 96028 95140
rect 95422 89584 95478 89593
rect 95422 89519 95478 89528
rect 95988 86834 96016 95134
rect 95976 86828 96028 86834
rect 95976 86770 96028 86776
rect 96632 79966 96660 124850
rect 96710 114064 96766 114073
rect 96710 113999 96766 114008
rect 96724 113830 96752 113999
rect 96712 113824 96764 113830
rect 96712 113766 96764 113772
rect 96620 79960 96672 79966
rect 96620 79902 96672 79908
rect 95332 71732 95384 71738
rect 95332 71674 95384 71680
rect 94688 69012 94740 69018
rect 94688 68954 94740 68960
rect 94504 59356 94556 59362
rect 94504 59298 94556 59304
rect 96620 24200 96672 24206
rect 96620 24142 96672 24148
rect 95240 19984 95292 19990
rect 95240 19926 95292 19932
rect 95252 16574 95280 19926
rect 88352 16546 89208 16574
rect 92492 16546 92796 16574
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 87604 9036 87656 9042
rect 87604 8978 87656 8984
rect 87800 598 88012 626
rect 87800 490 87828 598
rect 86838 -960 86950 480
rect 87524 462 87828 490
rect 87984 480 88012 598
rect 89180 480 89208 16546
rect 91560 15904 91612 15910
rect 91560 15846 91612 15852
rect 89904 13116 89956 13122
rect 89904 13058 89956 13064
rect 89916 490 89944 13058
rect 90192 598 90404 626
rect 90192 490 90220 598
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 462 90220 490
rect 90376 480 90404 598
rect 91572 480 91600 15846
rect 92768 480 92796 16546
rect 93952 2168 94004 2174
rect 93952 2110 94004 2116
rect 93964 480 93992 2110
rect 94700 490 94728 16546
rect 94976 598 95188 626
rect 94976 490 95004 598
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 462 95004 490
rect 95160 480 95188 598
rect 95804 490 95832 16546
rect 96632 6914 96660 24142
rect 96724 14550 96752 113766
rect 96816 84833 96844 130358
rect 97276 128354 97304 156402
rect 97828 147150 97856 195230
rect 97920 156466 97948 233854
rect 98012 220794 98040 238726
rect 98000 220788 98052 220794
rect 98000 220730 98052 220736
rect 98000 202836 98052 202842
rect 98000 202778 98052 202784
rect 98012 202162 98040 202778
rect 98000 202156 98052 202162
rect 98000 202098 98052 202104
rect 97908 156460 97960 156466
rect 97908 156402 97960 156408
rect 97920 155990 97948 156402
rect 97908 155984 97960 155990
rect 97908 155926 97960 155932
rect 97816 147144 97868 147150
rect 97816 147086 97868 147092
rect 97448 146940 97500 146946
rect 97448 146882 97500 146888
rect 97354 144800 97410 144809
rect 97354 144735 97410 144744
rect 97368 131481 97396 144735
rect 97460 135250 97488 146882
rect 97448 135244 97500 135250
rect 97448 135186 97500 135192
rect 97354 131472 97410 131481
rect 97354 131407 97410 131416
rect 97184 128326 97304 128354
rect 97184 123321 97212 128326
rect 97460 127673 97488 135186
rect 97632 128308 97684 128314
rect 97632 128250 97684 128256
rect 97446 127664 97502 127673
rect 97446 127599 97502 127608
rect 97644 127129 97672 128250
rect 97630 127120 97686 127129
rect 97630 127055 97686 127064
rect 97264 126948 97316 126954
rect 97264 126890 97316 126896
rect 97276 126313 97304 126890
rect 97262 126304 97318 126313
rect 97262 126239 97318 126248
rect 97540 125588 97592 125594
rect 97540 125530 97592 125536
rect 97552 124681 97580 125530
rect 97538 124672 97594 124681
rect 97538 124607 97594 124616
rect 97908 124160 97960 124166
rect 97906 124128 97908 124137
rect 97960 124128 97962 124137
rect 97906 124063 97962 124072
rect 97170 123312 97226 123321
rect 97170 123247 97226 123256
rect 97540 122800 97592 122806
rect 97540 122742 97592 122748
rect 97552 122505 97580 122742
rect 97538 122496 97594 122505
rect 97538 122431 97594 122440
rect 97724 121440 97776 121446
rect 97724 121382 97776 121388
rect 97736 120873 97764 121382
rect 97722 120864 97778 120873
rect 97722 120799 97778 120808
rect 97538 120320 97594 120329
rect 97538 120255 97594 120264
rect 97552 120154 97580 120255
rect 97540 120148 97592 120154
rect 97540 120090 97592 120096
rect 97724 120080 97776 120086
rect 97724 120022 97776 120028
rect 97736 119513 97764 120022
rect 97722 119504 97778 119513
rect 97722 119439 97778 119448
rect 97906 118688 97962 118697
rect 97906 118623 97908 118632
rect 97960 118623 97962 118632
rect 97908 118594 97960 118600
rect 97816 117972 97868 117978
rect 97816 117914 97868 117920
rect 97356 117292 97408 117298
rect 97356 117234 97408 117240
rect 97368 117065 97396 117234
rect 97354 117056 97410 117065
rect 97354 116991 97410 117000
rect 97828 114889 97856 117914
rect 97908 117224 97960 117230
rect 97908 117166 97960 117172
rect 97920 116521 97948 117166
rect 97906 116512 97962 116521
rect 97906 116447 97962 116456
rect 97906 115696 97962 115705
rect 97906 115631 97962 115640
rect 97814 114880 97870 114889
rect 97814 114815 97870 114824
rect 97540 114640 97592 114646
rect 97540 114582 97592 114588
rect 97552 113529 97580 114582
rect 97920 114578 97948 115631
rect 97908 114572 97960 114578
rect 97908 114514 97960 114520
rect 97538 113520 97594 113529
rect 97538 113455 97594 113464
rect 97906 112704 97962 112713
rect 97906 112639 97962 112648
rect 96896 111920 96948 111926
rect 96894 111888 96896 111897
rect 96948 111888 96950 111897
rect 97920 111858 97948 112639
rect 96894 111823 96950 111832
rect 97908 111852 97960 111858
rect 97908 111794 97960 111800
rect 97356 111784 97408 111790
rect 97356 111726 97408 111732
rect 97368 111081 97396 111726
rect 97354 111072 97410 111081
rect 97354 111007 97410 111016
rect 97814 109712 97870 109721
rect 97814 109647 97870 109656
rect 96986 107264 97042 107273
rect 96986 107199 97042 107208
rect 97000 106690 97028 107199
rect 97828 106962 97856 109647
rect 97908 108996 97960 109002
rect 97908 108938 97960 108944
rect 97920 108089 97948 108938
rect 97906 108080 97962 108089
rect 97906 108015 97962 108024
rect 97816 106956 97868 106962
rect 97816 106898 97868 106904
rect 96988 106684 97040 106690
rect 96988 106626 97040 106632
rect 97540 106072 97592 106078
rect 97540 106014 97592 106020
rect 96896 105936 96948 105942
rect 97552 105913 97580 106014
rect 96896 105878 96948 105884
rect 97538 105904 97594 105913
rect 96908 105097 96936 105878
rect 97538 105839 97594 105848
rect 96894 105088 96950 105097
rect 96894 105023 96950 105032
rect 97724 104848 97776 104854
rect 97724 104790 97776 104796
rect 97736 104281 97764 104790
rect 97722 104272 97778 104281
rect 97722 104207 97778 104216
rect 97908 103080 97960 103086
rect 97908 103022 97960 103028
rect 97920 102921 97948 103022
rect 97906 102912 97962 102921
rect 97906 102847 97962 102856
rect 97906 102096 97962 102105
rect 97906 102031 97908 102040
rect 97960 102031 97962 102040
rect 97908 102002 97960 102008
rect 97906 101280 97962 101289
rect 98012 101266 98040 202098
rect 98092 111988 98144 111994
rect 98092 111930 98144 111936
rect 98104 110265 98132 111930
rect 98656 111926 98684 245618
rect 98748 240038 98776 251126
rect 99392 246362 99420 258975
rect 99380 246356 99432 246362
rect 99380 246298 99432 246304
rect 99392 245682 99420 246298
rect 99380 245676 99432 245682
rect 99380 245618 99432 245624
rect 98736 240032 98788 240038
rect 98736 239974 98788 239980
rect 99484 233918 99512 271215
rect 100036 267714 100064 284378
rect 100128 273970 100156 289847
rect 100944 283620 100996 283626
rect 100944 283562 100996 283568
rect 100206 283384 100262 283393
rect 100206 283319 100262 283328
rect 100220 277302 100248 283319
rect 100850 282704 100906 282713
rect 100850 282639 100906 282648
rect 100758 281888 100814 281897
rect 100758 281823 100814 281832
rect 100772 281654 100800 281823
rect 100760 281648 100812 281654
rect 100760 281590 100812 281596
rect 100864 281586 100892 282639
rect 100852 281580 100904 281586
rect 100852 281522 100904 281528
rect 100850 281072 100906 281081
rect 100850 281007 100906 281016
rect 100760 280084 100812 280090
rect 100760 280026 100812 280032
rect 100772 279449 100800 280026
rect 100758 279440 100814 279449
rect 100758 279375 100814 279384
rect 100864 278118 100892 281007
rect 100852 278112 100904 278118
rect 100852 278054 100904 278060
rect 100956 277930 100984 283562
rect 100772 277902 100984 277930
rect 100772 277817 100800 277902
rect 100758 277808 100814 277817
rect 100758 277743 100814 277752
rect 100208 277296 100260 277302
rect 100208 277238 100260 277244
rect 100116 273964 100168 273970
rect 100116 273906 100168 273912
rect 100024 267708 100076 267714
rect 100024 267650 100076 267656
rect 100022 262304 100078 262313
rect 100022 262239 100078 262248
rect 99562 249248 99618 249257
rect 99562 249183 99618 249192
rect 99472 233912 99524 233918
rect 99472 233854 99524 233860
rect 98734 223544 98790 223553
rect 98734 223479 98790 223488
rect 98748 222329 98776 223479
rect 98734 222320 98790 222329
rect 98734 222255 98790 222264
rect 98644 111920 98696 111926
rect 98644 111862 98696 111868
rect 98090 110256 98146 110265
rect 98090 110191 98146 110200
rect 98748 105942 98776 222255
rect 98920 220788 98972 220794
rect 98920 220730 98972 220736
rect 98932 220046 98960 220730
rect 98920 220040 98972 220046
rect 98920 219982 98972 219988
rect 98828 211200 98880 211206
rect 98828 211142 98880 211148
rect 98736 105936 98788 105942
rect 98736 105878 98788 105884
rect 98734 104136 98790 104145
rect 98734 104071 98790 104080
rect 97962 101238 98040 101266
rect 97906 101215 97962 101224
rect 97908 100700 97960 100706
rect 97908 100642 97960 100648
rect 97538 100464 97594 100473
rect 97538 100399 97594 100408
rect 97552 99414 97580 100399
rect 97920 99657 97948 100642
rect 97906 99648 97962 99657
rect 97906 99583 97962 99592
rect 98642 99512 98698 99521
rect 98642 99447 98698 99456
rect 97540 99408 97592 99414
rect 97540 99350 97592 99356
rect 96894 99104 96950 99113
rect 96894 99039 96950 99048
rect 96908 98394 96936 99039
rect 96896 98388 96948 98394
rect 96896 98330 96948 98336
rect 97354 98288 97410 98297
rect 97354 98223 97410 98232
rect 97368 98054 97396 98223
rect 97356 98048 97408 98054
rect 97356 97990 97408 97996
rect 97906 97472 97962 97481
rect 97906 97407 97962 97416
rect 96896 96892 96948 96898
rect 96896 96834 96948 96840
rect 96908 96665 96936 96834
rect 97920 96694 97948 97407
rect 97908 96688 97960 96694
rect 96894 96656 96950 96665
rect 97908 96630 97960 96636
rect 96894 96591 96950 96600
rect 97262 95296 97318 95305
rect 97262 95231 97318 95240
rect 96988 94512 97040 94518
rect 96986 94480 96988 94489
rect 97040 94480 97042 94489
rect 96986 94415 97042 94424
rect 96802 84824 96858 84833
rect 96802 84759 96858 84768
rect 97276 64870 97304 95231
rect 97908 93832 97960 93838
rect 97908 93774 97960 93780
rect 97920 93673 97948 93774
rect 97906 93664 97962 93673
rect 97906 93599 97962 93608
rect 98656 82793 98684 99447
rect 98748 89622 98776 104071
rect 98840 96898 98868 211142
rect 98932 202842 98960 219982
rect 98920 202836 98972 202842
rect 98920 202778 98972 202784
rect 99576 103086 99604 249183
rect 100036 117978 100064 262239
rect 100668 247036 100720 247042
rect 100668 246978 100720 246984
rect 100680 245993 100708 246978
rect 100666 245984 100722 245993
rect 100666 245919 100722 245928
rect 100024 117972 100076 117978
rect 100024 117914 100076 117920
rect 100024 106684 100076 106690
rect 100024 106626 100076 106632
rect 99564 103080 99616 103086
rect 99564 103022 99616 103028
rect 99576 102814 99604 103022
rect 99564 102808 99616 102814
rect 99564 102750 99616 102756
rect 98920 98388 98972 98394
rect 98920 98330 98972 98336
rect 98828 96892 98880 96898
rect 98828 96834 98880 96840
rect 98736 89616 98788 89622
rect 98736 89558 98788 89564
rect 98932 82793 98960 98330
rect 100036 93129 100064 106626
rect 100680 102202 100708 245919
rect 100772 230489 100800 277743
rect 100852 277364 100904 277370
rect 100852 277306 100904 277312
rect 100864 276185 100892 277306
rect 101034 276992 101090 277001
rect 101034 276927 101090 276936
rect 100850 276176 100906 276185
rect 100850 276111 100906 276120
rect 100942 275360 100998 275369
rect 100942 275295 100998 275304
rect 100956 274718 100984 275295
rect 101048 275233 101076 276927
rect 101034 275224 101090 275233
rect 101034 275159 101090 275168
rect 100944 274712 100996 274718
rect 100944 274654 100996 274660
rect 100852 274644 100904 274650
rect 100852 274586 100904 274592
rect 100864 274553 100892 274586
rect 100850 274544 100906 274553
rect 100850 274479 100906 274488
rect 101416 273737 101444 341498
rect 102060 305046 102088 381482
rect 102244 355978 102272 390374
rect 103334 382936 103390 382945
rect 103334 382871 103390 382880
rect 102232 355972 102284 355978
rect 102232 355914 102284 355920
rect 101496 305040 101548 305046
rect 101496 304982 101548 304988
rect 102048 305040 102100 305046
rect 102048 304982 102100 304988
rect 101402 273728 101458 273737
rect 101402 273663 101458 273672
rect 100850 272912 100906 272921
rect 100850 272847 100906 272856
rect 100864 272542 100892 272847
rect 100852 272536 100904 272542
rect 100852 272478 100904 272484
rect 101508 271289 101536 304982
rect 102140 287088 102192 287094
rect 102140 287030 102192 287036
rect 101494 271280 101550 271289
rect 101494 271215 101550 271224
rect 100852 270496 100904 270502
rect 100850 270464 100852 270473
rect 100904 270464 100906 270473
rect 100850 270399 100906 270408
rect 100850 268016 100906 268025
rect 100850 267951 100906 267960
rect 100864 267782 100892 267951
rect 100852 267776 100904 267782
rect 100852 267718 100904 267724
rect 101404 267028 101456 267034
rect 101404 266970 101456 266976
rect 101034 266384 101090 266393
rect 101034 266319 101090 266328
rect 100850 265568 100906 265577
rect 100850 265503 100906 265512
rect 100864 264994 100892 265503
rect 100852 264988 100904 264994
rect 100852 264930 100904 264936
rect 100942 264752 100998 264761
rect 100942 264687 100998 264696
rect 100956 263634 100984 264687
rect 100944 263628 100996 263634
rect 100944 263570 100996 263576
rect 100852 263560 100904 263566
rect 100852 263502 100904 263508
rect 100864 263129 100892 263502
rect 100850 263120 100906 263129
rect 100850 263055 100906 263064
rect 100852 261520 100904 261526
rect 100850 261488 100852 261497
rect 101048 261497 101076 266319
rect 101128 265668 101180 265674
rect 101128 265610 101180 265616
rect 101140 262313 101168 265610
rect 101126 262304 101182 262313
rect 101126 262239 101182 262248
rect 100904 261488 100906 261497
rect 100850 261423 100906 261432
rect 101034 261488 101090 261497
rect 101034 261423 101090 261432
rect 100850 260672 100906 260681
rect 100850 260607 100906 260616
rect 100864 259486 100892 260607
rect 100852 259480 100904 259486
rect 100852 259422 100904 259428
rect 101416 257417 101444 266970
rect 101954 259856 102010 259865
rect 101954 259791 102010 259800
rect 101402 257408 101458 257417
rect 101968 257378 101996 259791
rect 101402 257343 101458 257352
rect 101956 257372 102008 257378
rect 100852 256692 100904 256698
rect 100852 256634 100904 256640
rect 100864 255785 100892 256634
rect 100942 256592 100998 256601
rect 100942 256527 100998 256536
rect 100850 255776 100906 255785
rect 100850 255711 100906 255720
rect 100956 255338 100984 256527
rect 100944 255332 100996 255338
rect 100944 255274 100996 255280
rect 100852 255264 100904 255270
rect 100852 255206 100904 255212
rect 100864 254969 100892 255206
rect 100850 254960 100906 254969
rect 100850 254895 100906 254904
rect 100850 253328 100906 253337
rect 100850 253263 100906 253272
rect 100864 252618 100892 253263
rect 100852 252612 100904 252618
rect 100852 252554 100904 252560
rect 100852 251116 100904 251122
rect 100852 251058 100904 251064
rect 100864 250889 100892 251058
rect 100850 250880 100906 250889
rect 100850 250815 100906 250824
rect 100942 250064 100998 250073
rect 100942 249999 100998 250008
rect 100852 249756 100904 249762
rect 100852 249698 100904 249704
rect 100864 248441 100892 249698
rect 100850 248432 100906 248441
rect 100850 248367 100906 248376
rect 100852 245540 100904 245546
rect 100852 245482 100904 245488
rect 100864 245177 100892 245482
rect 100850 245168 100906 245177
rect 100850 245103 100906 245112
rect 100850 243536 100906 243545
rect 100850 243471 100906 243480
rect 100864 243030 100892 243471
rect 100852 243024 100904 243030
rect 100852 242966 100904 242972
rect 100850 242720 100906 242729
rect 100850 242655 100906 242664
rect 100864 242146 100892 242655
rect 100852 242140 100904 242146
rect 100852 242082 100904 242088
rect 100956 238754 100984 249999
rect 101036 245608 101088 245614
rect 101036 245550 101088 245556
rect 101048 244361 101076 245550
rect 101034 244352 101090 244361
rect 101034 244287 101090 244296
rect 100864 238726 100984 238754
rect 100758 230480 100814 230489
rect 100758 230415 100814 230424
rect 100864 227798 100892 238726
rect 100852 227792 100904 227798
rect 100852 227734 100904 227740
rect 101416 167074 101444 257343
rect 101956 257314 102008 257320
rect 101494 216744 101550 216753
rect 101494 216679 101550 216688
rect 101404 167068 101456 167074
rect 101404 167010 101456 167016
rect 100758 151056 100814 151065
rect 100758 150991 100814 151000
rect 100668 102196 100720 102202
rect 100668 102138 100720 102144
rect 100680 100706 100708 102138
rect 100668 100700 100720 100706
rect 100668 100642 100720 100648
rect 100116 98116 100168 98122
rect 100116 98058 100168 98064
rect 100022 93120 100078 93129
rect 100022 93055 100078 93064
rect 100128 86601 100156 98058
rect 100772 88262 100800 150991
rect 101404 147144 101456 147150
rect 101404 147086 101456 147092
rect 100760 88256 100812 88262
rect 100760 88198 100812 88204
rect 100114 86592 100170 86601
rect 100114 86527 100170 86536
rect 98642 82784 98698 82793
rect 98642 82719 98698 82728
rect 98918 82784 98974 82793
rect 98918 82719 98974 82728
rect 98644 79348 98696 79354
rect 98644 79290 98696 79296
rect 97264 64864 97316 64870
rect 97264 64806 97316 64812
rect 97264 51740 97316 51746
rect 97264 51682 97316 51688
rect 96712 14544 96764 14550
rect 96712 14486 96764 14492
rect 96632 6886 97212 6914
rect 97184 1986 97212 6886
rect 97276 2106 97304 51682
rect 98000 37936 98052 37942
rect 98000 37878 98052 37884
rect 98012 16574 98040 37878
rect 98012 16546 98224 16574
rect 97264 2100 97316 2106
rect 97264 2042 97316 2048
rect 97184 1958 97488 1986
rect 96080 598 96292 626
rect 96080 490 96108 598
rect 95118 -960 95230 480
rect 95804 462 96108 490
rect 96264 480 96292 598
rect 97460 480 97488 1958
rect 98196 490 98224 16546
rect 98656 3534 98684 79290
rect 99380 43444 99432 43450
rect 99380 43386 99432 43392
rect 99392 16574 99420 43386
rect 99392 16546 99880 16574
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 98472 598 98684 626
rect 98472 490 98500 598
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 462 98500 490
rect 98656 480 98684 598
rect 99852 480 99880 16546
rect 101416 3534 101444 147086
rect 101508 106078 101536 216679
rect 101588 167068 101640 167074
rect 101588 167010 101640 167016
rect 101600 111994 101628 167010
rect 102152 149802 102180 287030
rect 103348 281489 103376 382871
rect 103440 356726 103468 390374
rect 103900 387802 103928 390374
rect 105266 390416 105322 390425
rect 104310 390374 104572 390402
rect 104880 390374 105216 390402
rect 104254 390351 104310 390360
rect 104268 390291 104296 390351
rect 103888 387796 103940 387802
rect 103888 387738 103940 387744
rect 104544 383654 104572 390374
rect 104808 389836 104860 389842
rect 104808 389778 104860 389784
rect 104544 383626 104756 383654
rect 104728 364342 104756 383626
rect 104716 364336 104768 364342
rect 104716 364278 104768 364284
rect 103520 362228 103572 362234
rect 103520 362170 103572 362176
rect 103428 356720 103480 356726
rect 103428 356662 103480 356668
rect 103428 355972 103480 355978
rect 103428 355914 103480 355920
rect 103334 281480 103390 281489
rect 103334 281415 103390 281424
rect 103348 280265 103376 281415
rect 103334 280256 103390 280265
rect 103334 280191 103390 280200
rect 103440 251190 103468 355914
rect 103428 251184 103480 251190
rect 103428 251126 103480 251132
rect 102784 243024 102836 243030
rect 102784 242966 102836 242972
rect 102796 222902 102824 242966
rect 102876 242956 102928 242962
rect 102876 242898 102928 242904
rect 102888 238746 102916 242898
rect 103428 241528 103480 241534
rect 103428 241470 103480 241476
rect 103440 240038 103468 241470
rect 103428 240032 103480 240038
rect 103428 239974 103480 239980
rect 103532 239465 103560 362170
rect 104820 322250 104848 389778
rect 105188 388657 105216 390374
rect 105322 390374 106044 390402
rect 105266 390351 105322 390360
rect 105174 388648 105230 388657
rect 105174 388583 105230 388592
rect 106016 379409 106044 390374
rect 106002 379400 106058 379409
rect 106002 379335 106058 379344
rect 104808 322244 104860 322250
rect 104808 322186 104860 322192
rect 104164 312656 104216 312662
rect 104164 312598 104216 312604
rect 104176 305658 104204 312598
rect 104164 305652 104216 305658
rect 104164 305594 104216 305600
rect 104716 305652 104768 305658
rect 104716 305594 104768 305600
rect 104624 287768 104676 287774
rect 104624 287710 104676 287716
rect 104164 268388 104216 268394
rect 104164 268330 104216 268336
rect 103612 242140 103664 242146
rect 103612 242082 103664 242088
rect 103518 239456 103574 239465
rect 103518 239391 103574 239400
rect 102876 238740 102928 238746
rect 102876 238682 102928 238688
rect 103532 236745 103560 239391
rect 103518 236736 103574 236745
rect 103518 236671 103574 236680
rect 102784 222896 102836 222902
rect 102784 222838 102836 222844
rect 103624 212498 103652 242082
rect 104176 233209 104204 268330
rect 104636 261526 104664 287710
rect 104728 272513 104756 305594
rect 104714 272504 104770 272513
rect 104714 272439 104770 272448
rect 104820 268258 104848 322186
rect 105636 278044 105688 278050
rect 105636 277986 105688 277992
rect 104808 268252 104860 268258
rect 104808 268194 104860 268200
rect 105544 268252 105596 268258
rect 105544 268194 105596 268200
rect 104820 267782 104848 268194
rect 104808 267776 104860 267782
rect 104808 267718 104860 267724
rect 104808 262132 104860 262138
rect 104808 262074 104860 262080
rect 104624 261520 104676 261526
rect 104624 261462 104676 261468
rect 104820 251802 104848 262074
rect 104256 251796 104308 251802
rect 104256 251738 104308 251744
rect 104808 251796 104860 251802
rect 104808 251738 104860 251744
rect 104268 246809 104296 251738
rect 104820 251258 104848 251738
rect 104808 251252 104860 251258
rect 104808 251194 104860 251200
rect 104254 246800 104310 246809
rect 104254 246735 104310 246744
rect 104162 233200 104218 233209
rect 104162 233135 104218 233144
rect 104162 220144 104218 220153
rect 104162 220079 104218 220088
rect 103612 212492 103664 212498
rect 103612 212434 103664 212440
rect 103624 211206 103652 212434
rect 103612 211200 103664 211206
rect 103612 211142 103664 211148
rect 102232 207052 102284 207058
rect 102232 206994 102284 207000
rect 102140 149796 102192 149802
rect 102140 149738 102192 149744
rect 101588 111988 101640 111994
rect 101588 111930 101640 111936
rect 101496 106072 101548 106078
rect 101496 106014 101548 106020
rect 102244 94518 102272 206994
rect 103520 188352 103572 188358
rect 103520 188294 103572 188300
rect 102782 151056 102838 151065
rect 102782 150991 102838 151000
rect 102324 144220 102376 144226
rect 102324 144162 102376 144168
rect 102232 94512 102284 94518
rect 102232 94454 102284 94460
rect 102336 16574 102364 144162
rect 102796 117881 102824 150991
rect 102966 150512 103022 150521
rect 102966 150447 103022 150456
rect 102980 130218 103008 150447
rect 102968 130212 103020 130218
rect 102968 130154 103020 130160
rect 102782 117872 102838 117881
rect 102782 117807 102838 117816
rect 103532 73166 103560 188294
rect 104176 90409 104204 220079
rect 104992 206372 105044 206378
rect 104992 206314 105044 206320
rect 104254 150648 104310 150657
rect 104254 150583 104310 150592
rect 104268 112470 104296 150583
rect 104256 112464 104308 112470
rect 104256 112406 104308 112412
rect 104256 109744 104308 109750
rect 104256 109686 104308 109692
rect 104162 90400 104218 90409
rect 104162 90335 104218 90344
rect 103520 73160 103572 73166
rect 103520 73102 103572 73108
rect 103518 30968 103574 30977
rect 103518 30903 103574 30912
rect 103532 16574 103560 30903
rect 102336 16546 103376 16574
rect 103532 16546 104112 16574
rect 101404 3528 101456 3534
rect 101034 3496 101090 3505
rect 101404 3470 101456 3476
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 101034 3431 101090 3440
rect 101048 480 101076 3431
rect 102244 480 102272 3470
rect 103348 480 103376 16546
rect 104084 490 104112 16546
rect 104268 3466 104296 109686
rect 104900 108384 104952 108390
rect 104900 108326 104952 108332
rect 104530 90400 104586 90409
rect 104530 90335 104586 90344
rect 104544 89457 104572 90335
rect 104530 89448 104586 89457
rect 104530 89383 104586 89392
rect 104912 16574 104940 108326
rect 105004 83881 105032 206314
rect 105084 178696 105136 178702
rect 105084 178638 105136 178644
rect 105096 91089 105124 178638
rect 105556 157418 105584 268194
rect 105648 241398 105676 277986
rect 106108 267073 106136 390918
rect 107382 390895 107438 390904
rect 111982 390552 112038 390561
rect 111872 390510 111982 390538
rect 111982 390487 112038 390496
rect 106338 390130 106366 390388
rect 107626 390266 107654 390388
rect 107764 390374 108376 390402
rect 107626 390238 107700 390266
rect 106292 390102 106366 390130
rect 106188 387116 106240 387122
rect 106188 387058 106240 387064
rect 106200 383790 106228 387058
rect 106188 383784 106240 383790
rect 106188 383726 106240 383732
rect 106094 267064 106150 267073
rect 106094 266999 106150 267008
rect 106108 266393 106136 266999
rect 106094 266384 106150 266393
rect 106094 266319 106150 266328
rect 105636 241392 105688 241398
rect 105636 241334 105688 241340
rect 106200 238377 106228 383726
rect 106292 241534 106320 390102
rect 107672 389230 107700 390238
rect 107660 389224 107712 389230
rect 107660 389166 107712 389172
rect 107764 380905 107792 390374
rect 109098 390130 109126 390388
rect 109512 390374 109848 390402
rect 109098 390102 109172 390130
rect 108302 389872 108358 389881
rect 108302 389807 108358 389816
rect 107750 380896 107806 380905
rect 107750 380831 107806 380840
rect 107568 373312 107620 373318
rect 107568 373254 107620 373260
rect 107580 349858 107608 373254
rect 107568 349852 107620 349858
rect 107568 349794 107620 349800
rect 106922 317520 106978 317529
rect 106922 317455 106978 317464
rect 106280 241528 106332 241534
rect 106280 241470 106332 241476
rect 106186 238368 106242 238377
rect 106186 238303 106242 238312
rect 106200 237425 106228 238303
rect 106280 238128 106332 238134
rect 106280 238070 106332 238076
rect 106186 237416 106242 237425
rect 106186 237351 106242 237360
rect 105728 206372 105780 206378
rect 105728 206314 105780 206320
rect 105740 205698 105768 206314
rect 105728 205692 105780 205698
rect 105728 205634 105780 205640
rect 105544 157412 105596 157418
rect 105544 157354 105596 157360
rect 105556 120154 105584 157354
rect 105636 140820 105688 140826
rect 105636 140762 105688 140768
rect 105648 132462 105676 140762
rect 105636 132456 105688 132462
rect 105636 132398 105688 132404
rect 105544 120148 105596 120154
rect 105544 120090 105596 120096
rect 105082 91080 105138 91089
rect 105082 91015 105138 91024
rect 105634 89856 105690 89865
rect 105634 89791 105690 89800
rect 105544 89752 105596 89758
rect 105544 89694 105596 89700
rect 104990 83872 105046 83881
rect 104990 83807 105046 83816
rect 105556 82754 105584 89694
rect 105544 82748 105596 82754
rect 105544 82690 105596 82696
rect 105556 56506 105584 82690
rect 105648 80073 105676 89791
rect 105634 80064 105690 80073
rect 105634 79999 105690 80008
rect 105544 56500 105596 56506
rect 105544 56442 105596 56448
rect 106292 16574 106320 238070
rect 106936 228750 106964 317455
rect 107580 251122 107608 349794
rect 108212 311228 108264 311234
rect 108212 311170 108264 311176
rect 108224 308446 108252 311170
rect 108212 308440 108264 308446
rect 108212 308382 108264 308388
rect 108316 269249 108344 389807
rect 109040 387048 109092 387054
rect 109040 386990 109092 386996
rect 108948 376032 109000 376038
rect 108948 375974 109000 375980
rect 108960 352578 108988 375974
rect 109052 371385 109080 386990
rect 109144 383042 109172 390102
rect 109512 387054 109540 390374
rect 110386 390130 110414 390388
rect 110524 390374 111136 390402
rect 111996 390374 112608 390402
rect 110386 390102 110460 390130
rect 110432 387122 110460 390102
rect 110420 387116 110472 387122
rect 110420 387058 110472 387064
rect 109500 387048 109552 387054
rect 110524 387002 110552 390374
rect 109500 386990 109552 386996
rect 110432 386974 110552 387002
rect 109132 383036 109184 383042
rect 109132 382978 109184 382984
rect 109682 371920 109738 371929
rect 109682 371855 109738 371864
rect 109696 371385 109724 371855
rect 109038 371376 109094 371385
rect 109038 371311 109094 371320
rect 109682 371376 109738 371385
rect 109682 371311 109738 371320
rect 108948 352572 109000 352578
rect 108948 352514 109000 352520
rect 108302 269240 108358 269249
rect 108302 269175 108358 269184
rect 108302 266384 108358 266393
rect 108302 266319 108358 266328
rect 107568 251116 107620 251122
rect 107568 251058 107620 251064
rect 107016 247716 107068 247722
rect 107016 247658 107068 247664
rect 107028 238513 107056 247658
rect 107014 238504 107070 238513
rect 107014 238439 107070 238448
rect 107658 234152 107714 234161
rect 107658 234087 107714 234096
rect 107568 229084 107620 229090
rect 107568 229026 107620 229032
rect 107580 228750 107608 229026
rect 106924 228744 106976 228750
rect 106924 228686 106976 228692
rect 107568 228744 107620 228750
rect 107568 228686 107620 228692
rect 106372 228404 106424 228410
rect 106372 228346 106424 228352
rect 106384 89758 106412 228346
rect 106924 178696 106976 178702
rect 106924 178638 106976 178644
rect 106372 89752 106424 89758
rect 106372 89694 106424 89700
rect 106936 68338 106964 178638
rect 107580 145586 107608 228686
rect 107568 145580 107620 145586
rect 107568 145522 107620 145528
rect 107672 92313 107700 234087
rect 108316 225690 108344 266319
rect 108488 258120 108540 258126
rect 108488 258062 108540 258068
rect 108396 253972 108448 253978
rect 108396 253914 108448 253920
rect 108408 245546 108436 253914
rect 108396 245540 108448 245546
rect 108396 245482 108448 245488
rect 108396 238060 108448 238066
rect 108396 238002 108448 238008
rect 108304 225684 108356 225690
rect 108304 225626 108356 225632
rect 108408 211818 108436 238002
rect 108500 234598 108528 258062
rect 108960 255270 108988 352514
rect 108948 255264 109000 255270
rect 108948 255206 109000 255212
rect 109696 253978 109724 371311
rect 110432 369782 110460 386974
rect 110510 385792 110566 385801
rect 110510 385727 110566 385736
rect 110420 369776 110472 369782
rect 110420 369718 110472 369724
rect 110420 356720 110472 356726
rect 110420 356662 110472 356668
rect 110432 356114 110460 356662
rect 110420 356108 110472 356114
rect 110420 356050 110472 356056
rect 109774 263664 109830 263673
rect 109774 263599 109830 263608
rect 109684 253972 109736 253978
rect 109684 253914 109736 253920
rect 109684 252612 109736 252618
rect 109684 252554 109736 252560
rect 109038 237416 109094 237425
rect 109038 237351 109094 237360
rect 108488 234592 108540 234598
rect 108488 234534 108540 234540
rect 108396 211812 108448 211818
rect 108396 211754 108448 211760
rect 108304 193860 108356 193866
rect 108304 193802 108356 193808
rect 107658 92304 107714 92313
rect 107658 92239 107714 92248
rect 106924 68332 106976 68338
rect 106924 68274 106976 68280
rect 108316 51814 108344 193802
rect 108408 93838 108436 211754
rect 108486 144936 108542 144945
rect 108486 144871 108542 144880
rect 108500 126274 108528 144871
rect 108488 126268 108540 126274
rect 108488 126210 108540 126216
rect 108396 93832 108448 93838
rect 108396 93774 108448 93780
rect 109052 88097 109080 237351
rect 109696 225622 109724 252554
rect 109788 242214 109816 263599
rect 109868 253972 109920 253978
rect 109868 253914 109920 253920
rect 109880 249762 109908 253914
rect 109868 249756 109920 249762
rect 109868 249698 109920 249704
rect 109880 249082 109908 249698
rect 109868 249076 109920 249082
rect 109868 249018 109920 249024
rect 109776 242208 109828 242214
rect 109776 242150 109828 242156
rect 110432 241466 110460 356050
rect 110420 241460 110472 241466
rect 110420 241402 110472 241408
rect 110420 238060 110472 238066
rect 110420 238002 110472 238008
rect 109684 225616 109736 225622
rect 109684 225558 109736 225564
rect 109038 88088 109094 88097
rect 109038 88023 109094 88032
rect 109040 68332 109092 68338
rect 109040 68274 109092 68280
rect 108396 64184 108448 64190
rect 108396 64126 108448 64132
rect 108304 51808 108356 51814
rect 108304 51750 108356 51756
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 104256 3460 104308 3466
rect 104256 3402 104308 3408
rect 104360 598 104572 626
rect 104360 490 104388 598
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 462 104388 490
rect 104544 480 104572 598
rect 105740 480 105768 16546
rect 106476 490 106504 16546
rect 108120 10464 108172 10470
rect 108120 10406 108172 10412
rect 106752 598 106964 626
rect 106752 490 106780 598
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 462 106780 490
rect 106936 480 106964 598
rect 108132 480 108160 10406
rect 108408 10402 108436 64126
rect 109052 16574 109080 68274
rect 110432 16574 110460 238002
rect 110524 236609 110552 385727
rect 111996 378146 112024 390374
rect 111984 378140 112036 378146
rect 111984 378082 112036 378088
rect 112444 378140 112496 378146
rect 112444 378082 112496 378088
rect 111064 369776 111116 369782
rect 111064 369718 111116 369724
rect 111076 262138 111104 369718
rect 111800 307828 111852 307834
rect 111800 307770 111852 307776
rect 111812 307154 111840 307770
rect 111800 307148 111852 307154
rect 111800 307090 111852 307096
rect 111800 266348 111852 266354
rect 111800 266290 111852 266296
rect 111812 265674 111840 266290
rect 111800 265668 111852 265674
rect 111800 265610 111852 265616
rect 111064 262132 111116 262138
rect 111064 262074 111116 262080
rect 112456 253978 112484 378082
rect 112534 283248 112590 283257
rect 112534 283183 112590 283192
rect 112444 253972 112496 253978
rect 112444 253914 112496 253920
rect 111800 253292 111852 253298
rect 111800 253234 111852 253240
rect 111064 251116 111116 251122
rect 111064 251058 111116 251064
rect 110510 236600 110566 236609
rect 110510 236535 110566 236544
rect 111076 104922 111104 251058
rect 111156 243568 111208 243574
rect 111156 243510 111208 243516
rect 111168 228410 111196 243510
rect 111156 228404 111208 228410
rect 111156 228346 111208 228352
rect 111156 227044 111208 227050
rect 111156 226986 111208 226992
rect 111064 104916 111116 104922
rect 111064 104858 111116 104864
rect 111168 89729 111196 226986
rect 111246 135960 111302 135969
rect 111246 135895 111302 135904
rect 111260 126954 111288 135895
rect 111248 126948 111300 126954
rect 111248 126890 111300 126896
rect 111154 89720 111210 89729
rect 111154 89655 111210 89664
rect 111812 16574 111840 253234
rect 112548 247790 112576 283183
rect 113100 266354 113128 407050
rect 113192 271930 113220 420815
rect 113284 304201 113312 428159
rect 113362 418976 113418 418985
rect 113362 418911 113418 418920
rect 113376 381546 113404 418911
rect 114480 406473 114508 449958
rect 114572 423065 114600 460158
rect 114928 430500 114980 430506
rect 114928 430442 114980 430448
rect 114940 429321 114968 430442
rect 114926 429312 114982 429321
rect 114926 429247 114982 429256
rect 115112 424992 115164 424998
rect 115110 424960 115112 424969
rect 115164 424960 115166 424969
rect 115110 424895 115166 424904
rect 114558 423056 114614 423065
rect 114558 422991 114614 423000
rect 114650 420064 114706 420073
rect 114650 419999 114706 420008
rect 114558 417888 114614 417897
rect 114558 417823 114614 417832
rect 114466 406464 114522 406473
rect 114466 406399 114522 406408
rect 113454 402384 113510 402393
rect 113454 402319 113510 402328
rect 113468 383722 113496 402319
rect 113456 383716 113508 383722
rect 113456 383658 113508 383664
rect 113364 381540 113416 381546
rect 113364 381482 113416 381488
rect 113468 373994 113496 383658
rect 113376 373966 113496 373994
rect 113376 367810 113404 373966
rect 114468 368484 114520 368490
rect 114468 368426 114520 368432
rect 114480 367810 114508 368426
rect 113364 367804 113416 367810
rect 113364 367746 113416 367752
rect 114468 367804 114520 367810
rect 114468 367746 114520 367752
rect 113270 304192 113326 304201
rect 113270 304127 113326 304136
rect 113824 292596 113876 292602
rect 113824 292538 113876 292544
rect 113180 271924 113232 271930
rect 113180 271866 113232 271872
rect 113088 266348 113140 266354
rect 113088 266290 113140 266296
rect 112720 257372 112772 257378
rect 112720 257314 112772 257320
rect 112626 254008 112682 254017
rect 112626 253943 112682 253952
rect 112536 247784 112588 247790
rect 112536 247726 112588 247732
rect 112640 221474 112668 253943
rect 112732 232529 112760 257314
rect 112718 232520 112774 232529
rect 112718 232455 112774 232464
rect 112628 221468 112680 221474
rect 112628 221410 112680 221416
rect 111892 204944 111944 204950
rect 111892 204886 111944 204892
rect 111904 204338 111932 204886
rect 111892 204332 111944 204338
rect 111892 204274 111944 204280
rect 111904 109585 111932 204274
rect 113836 175302 113864 292538
rect 114572 270502 114600 417823
rect 114664 305658 114692 419999
rect 114926 414896 114982 414905
rect 114926 414831 114982 414840
rect 114940 414730 114968 414831
rect 114928 414724 114980 414730
rect 114928 414666 114980 414672
rect 114836 400988 114888 400994
rect 114836 400930 114888 400936
rect 114848 400489 114876 400930
rect 114834 400480 114890 400489
rect 114834 400415 114890 400424
rect 114940 393314 114968 414666
rect 115216 413817 115244 558826
rect 115308 556850 115336 604415
rect 122840 590028 122892 590034
rect 122840 589970 122892 589976
rect 116584 589960 116636 589966
rect 116584 589902 116636 589908
rect 115296 556844 115348 556850
rect 115296 556786 115348 556792
rect 116214 554024 116270 554033
rect 116214 553959 116270 553968
rect 115294 516760 115350 516769
rect 115294 516695 115350 516704
rect 115308 468489 115336 516695
rect 115294 468480 115350 468489
rect 115294 468415 115350 468424
rect 115308 421977 115336 468415
rect 116032 436144 116084 436150
rect 116032 436086 116084 436092
rect 115756 434716 115808 434722
rect 115756 434658 115808 434664
rect 115768 433401 115796 434658
rect 115754 433392 115810 433401
rect 115754 433327 115810 433336
rect 115848 433288 115900 433294
rect 115848 433230 115900 433236
rect 115860 432313 115888 433230
rect 115846 432304 115902 432313
rect 115846 432239 115902 432248
rect 115848 429140 115900 429146
rect 115848 429082 115900 429088
rect 115860 428233 115888 429082
rect 115846 428224 115902 428233
rect 115846 428159 115902 428168
rect 115846 427136 115902 427145
rect 115846 427071 115902 427080
rect 115860 426494 115888 427071
rect 115848 426488 115900 426494
rect 115848 426430 115900 426436
rect 115756 426420 115808 426426
rect 115756 426362 115808 426368
rect 115768 426057 115796 426362
rect 115754 426048 115810 426057
rect 115754 425983 115810 425992
rect 115848 425060 115900 425066
rect 115848 425002 115900 425008
rect 115860 424153 115888 425002
rect 115846 424144 115902 424153
rect 115846 424079 115902 424088
rect 115848 423632 115900 423638
rect 115848 423574 115900 423580
rect 115860 423065 115888 423574
rect 115846 423056 115902 423065
rect 115846 422991 115902 423000
rect 115294 421968 115350 421977
rect 115294 421903 115350 421912
rect 115848 419484 115900 419490
rect 115848 419426 115900 419432
rect 115860 418985 115888 419426
rect 115846 418976 115902 418985
rect 115846 418911 115902 418920
rect 115848 416832 115900 416838
rect 115846 416800 115848 416809
rect 115900 416800 115902 416809
rect 115846 416735 115902 416744
rect 115846 415712 115902 415721
rect 115846 415647 115848 415656
rect 115900 415647 115902 415656
rect 115848 415618 115900 415624
rect 115202 413808 115258 413817
rect 115202 413743 115258 413752
rect 115846 412720 115902 412729
rect 115846 412655 115848 412664
rect 115900 412655 115902 412664
rect 115848 412626 115900 412632
rect 115756 412616 115808 412622
rect 115756 412558 115808 412564
rect 115768 411641 115796 412558
rect 115754 411632 115810 411641
rect 115754 411567 115810 411576
rect 115848 411256 115900 411262
rect 115848 411198 115900 411204
rect 115860 410553 115888 411198
rect 115846 410544 115902 410553
rect 115846 410479 115902 410488
rect 115940 409896 115992 409902
rect 115940 409838 115992 409844
rect 115848 409760 115900 409766
rect 115846 409728 115848 409737
rect 115900 409728 115902 409737
rect 115846 409663 115902 409672
rect 115846 408640 115902 408649
rect 115846 408575 115902 408584
rect 115860 408542 115888 408575
rect 115848 408536 115900 408542
rect 115848 408478 115900 408484
rect 115202 406464 115258 406473
rect 115202 406399 115258 406408
rect 114848 393286 114968 393314
rect 114848 389842 114876 393286
rect 114836 389836 114888 389842
rect 114836 389778 114888 389784
rect 115216 306474 115244 406399
rect 115846 405648 115902 405657
rect 115952 405634 115980 409838
rect 115902 405606 115980 405634
rect 115846 405583 115902 405592
rect 115846 404560 115902 404569
rect 115846 404495 115902 404504
rect 115860 404394 115888 404495
rect 115848 404388 115900 404394
rect 115848 404330 115900 404336
rect 115846 403472 115902 403481
rect 115846 403407 115902 403416
rect 115860 403034 115888 403407
rect 115848 403028 115900 403034
rect 115848 402970 115900 402976
rect 115940 402280 115992 402286
rect 115940 402222 115992 402228
rect 115386 401296 115442 401305
rect 115386 401231 115442 401240
rect 115400 400246 115428 401231
rect 115388 400240 115440 400246
rect 115388 400182 115440 400188
rect 115846 399392 115902 399401
rect 115952 399378 115980 402222
rect 115902 399350 115980 399378
rect 115846 399327 115902 399336
rect 115848 398336 115900 398342
rect 115846 398304 115848 398313
rect 115900 398304 115902 398313
rect 115846 398239 115902 398248
rect 115846 397216 115902 397225
rect 115846 397151 115902 397160
rect 115756 397112 115808 397118
rect 115756 397054 115808 397060
rect 115768 396409 115796 397054
rect 115754 396400 115810 396409
rect 115754 396335 115810 396344
rect 115860 396098 115888 397151
rect 115848 396092 115900 396098
rect 115848 396034 115900 396040
rect 115846 395312 115902 395321
rect 115846 395247 115902 395256
rect 115860 394806 115888 395247
rect 115848 394800 115900 394806
rect 115848 394742 115900 394748
rect 115848 394664 115900 394670
rect 115848 394606 115900 394612
rect 115860 394233 115888 394606
rect 115846 394224 115902 394233
rect 115846 394159 115902 394168
rect 115846 393136 115902 393145
rect 115902 393094 115980 393122
rect 115846 393071 115902 393080
rect 115952 392766 115980 393094
rect 115940 392760 115992 392766
rect 115940 392702 115992 392708
rect 115846 392048 115902 392057
rect 115846 391983 115848 391992
rect 115900 391983 115902 391992
rect 115848 391954 115900 391960
rect 115952 373318 115980 392702
rect 115940 373312 115992 373318
rect 115940 373254 115992 373260
rect 116044 312662 116072 436086
rect 116124 398336 116176 398342
rect 116124 398278 116176 398284
rect 116136 376038 116164 398278
rect 116228 385801 116256 553959
rect 116596 541686 116624 589902
rect 118700 585200 118752 585206
rect 118700 585142 118752 585148
rect 118712 585041 118740 585142
rect 118698 585032 118754 585041
rect 118698 584967 118754 584976
rect 119342 585032 119398 585041
rect 119342 584967 119398 584976
rect 116584 541680 116636 541686
rect 116584 541622 116636 541628
rect 117320 461644 117372 461650
rect 117320 461586 117372 461592
rect 117332 461009 117360 461586
rect 117318 461000 117374 461009
rect 117318 460935 117374 460944
rect 116584 451308 116636 451314
rect 116584 451250 116636 451256
rect 116596 436150 116624 451250
rect 116584 436144 116636 436150
rect 116584 436086 116636 436092
rect 117332 424998 117360 460935
rect 118698 436248 118754 436257
rect 118698 436183 118754 436192
rect 117504 426420 117556 426426
rect 117504 426362 117556 426368
rect 117320 424992 117372 424998
rect 117320 424934 117372 424940
rect 117412 417240 117464 417246
rect 117412 417182 117464 417188
rect 117424 416838 117452 417182
rect 117412 416832 117464 416838
rect 117412 416774 117464 416780
rect 117228 394052 117280 394058
rect 117228 393994 117280 394000
rect 117240 392766 117268 393994
rect 117228 392760 117280 392766
rect 117228 392702 117280 392708
rect 117424 389881 117452 416774
rect 117410 389872 117466 389881
rect 117410 389807 117466 389816
rect 116214 385792 116270 385801
rect 116214 385727 116270 385736
rect 116124 376032 116176 376038
rect 116124 375974 116176 375980
rect 116676 328500 116728 328506
rect 116676 328442 116728 328448
rect 116584 316056 116636 316062
rect 116584 315998 116636 316004
rect 116032 312656 116084 312662
rect 116032 312598 116084 312604
rect 116596 309194 116624 315998
rect 116584 309188 116636 309194
rect 116584 309130 116636 309136
rect 115204 306468 115256 306474
rect 115204 306410 115256 306416
rect 114652 305652 114704 305658
rect 114652 305594 114704 305600
rect 115216 287774 115244 306410
rect 115938 300248 115994 300257
rect 115938 300183 115994 300192
rect 115204 287768 115256 287774
rect 115204 287710 115256 287716
rect 115296 287768 115348 287774
rect 115296 287710 115348 287716
rect 115204 281648 115256 281654
rect 115204 281590 115256 281596
rect 114560 270496 114612 270502
rect 114560 270438 114612 270444
rect 113916 258188 113968 258194
rect 113916 258130 113968 258136
rect 113824 175296 113876 175302
rect 113824 175238 113876 175244
rect 112444 153332 112496 153338
rect 112444 153274 112496 153280
rect 112456 122126 112484 153274
rect 113836 138786 113864 175238
rect 113928 146402 113956 258130
rect 114652 255196 114704 255202
rect 114652 255138 114704 255144
rect 114560 188352 114612 188358
rect 114560 188294 114612 188300
rect 114006 161528 114062 161537
rect 114006 161463 114062 161472
rect 113916 146396 113968 146402
rect 113916 146338 113968 146344
rect 113824 138780 113876 138786
rect 113824 138722 113876 138728
rect 113824 133204 113876 133210
rect 113824 133146 113876 133152
rect 112444 122120 112496 122126
rect 112444 122062 112496 122068
rect 112444 114640 112496 114646
rect 112444 114582 112496 114588
rect 111890 109576 111946 109585
rect 111890 109511 111946 109520
rect 112456 67522 112484 114582
rect 113836 79354 113864 133146
rect 113928 111790 113956 146338
rect 114020 133890 114048 161463
rect 114008 133884 114060 133890
rect 114008 133826 114060 133832
rect 113916 111784 113968 111790
rect 113916 111726 113968 111732
rect 113916 101448 113968 101454
rect 113916 101390 113968 101396
rect 113928 88330 113956 101390
rect 113916 88324 113968 88330
rect 113916 88266 113968 88272
rect 113824 79348 113876 79354
rect 113824 79290 113876 79296
rect 112444 67516 112496 67522
rect 112444 67458 112496 67464
rect 113180 31068 113232 31074
rect 113180 31010 113232 31016
rect 113192 16574 113220 31010
rect 114572 16574 114600 188294
rect 114664 109002 114692 255138
rect 114744 231124 114796 231130
rect 114744 231066 114796 231072
rect 114652 108996 114704 109002
rect 114652 108938 114704 108944
rect 114756 104145 114784 231066
rect 115216 226953 115244 281590
rect 115308 281489 115336 287710
rect 115294 281480 115350 281489
rect 115294 281415 115350 281424
rect 115294 267880 115350 267889
rect 115294 267815 115350 267824
rect 115308 250510 115336 267815
rect 115296 250504 115348 250510
rect 115296 250446 115348 250452
rect 115202 226944 115258 226953
rect 115202 226879 115258 226888
rect 115848 108996 115900 109002
rect 115848 108938 115900 108944
rect 115860 108322 115888 108938
rect 115848 108316 115900 108322
rect 115848 108258 115900 108264
rect 114742 104136 114798 104145
rect 114742 104071 114798 104080
rect 115952 16574 115980 300183
rect 116596 222154 116624 309130
rect 116688 296070 116716 328442
rect 116676 296064 116728 296070
rect 116676 296006 116728 296012
rect 117228 296064 117280 296070
rect 117228 296006 117280 296012
rect 117240 289202 117268 296006
rect 117228 289196 117280 289202
rect 117228 289138 117280 289144
rect 116674 285832 116730 285841
rect 116674 285767 116730 285776
rect 116688 253230 116716 285767
rect 117516 275233 117544 426362
rect 118608 393984 118660 393990
rect 118608 393926 118660 393932
rect 118620 389230 118648 393926
rect 118608 389224 118660 389230
rect 118608 389166 118660 389172
rect 118712 311234 118740 436183
rect 119356 426426 119384 584967
rect 122102 582720 122158 582729
rect 122102 582655 122158 582664
rect 119436 575544 119488 575550
rect 119436 575486 119488 575492
rect 119448 538218 119476 575486
rect 122116 538898 122144 582655
rect 122104 538892 122156 538898
rect 122104 538834 122156 538840
rect 119436 538212 119488 538218
rect 119436 538154 119488 538160
rect 122104 529304 122156 529310
rect 122104 529246 122156 529252
rect 119344 426420 119396 426426
rect 119344 426362 119396 426368
rect 122116 419422 122144 529246
rect 122748 484424 122800 484430
rect 122748 484366 122800 484372
rect 122196 452736 122248 452742
rect 122196 452678 122248 452684
rect 122208 440910 122236 452678
rect 122760 451897 122788 484366
rect 122746 451888 122802 451897
rect 122746 451823 122802 451832
rect 122760 451353 122788 451823
rect 122746 451344 122802 451353
rect 122746 451279 122802 451288
rect 122196 440904 122248 440910
rect 122196 440846 122248 440852
rect 122196 427100 122248 427106
rect 122196 427042 122248 427048
rect 122104 419416 122156 419422
rect 122104 419358 122156 419364
rect 122208 417246 122236 427042
rect 122196 417240 122248 417246
rect 122196 417182 122248 417188
rect 122104 416084 122156 416090
rect 122104 416026 122156 416032
rect 120080 415676 120132 415682
rect 120080 415618 120132 415624
rect 119344 406428 119396 406434
rect 119344 406370 119396 406376
rect 118792 400920 118844 400926
rect 118792 400862 118844 400868
rect 118804 398342 118832 400862
rect 118792 398336 118844 398342
rect 118792 398278 118844 398284
rect 118792 398132 118844 398138
rect 118792 398074 118844 398080
rect 118804 397118 118832 398074
rect 118792 397112 118844 397118
rect 118792 397054 118844 397060
rect 119356 383489 119384 406370
rect 119988 403096 120040 403102
rect 119988 403038 120040 403044
rect 120000 400994 120028 403038
rect 119988 400988 120040 400994
rect 119988 400930 120040 400936
rect 119342 383480 119398 383489
rect 119342 383415 119398 383424
rect 120092 378026 120120 415618
rect 122116 409766 122144 416026
rect 122104 409760 122156 409766
rect 122104 409702 122156 409708
rect 122104 400240 122156 400246
rect 122104 400182 122156 400188
rect 121644 378820 121696 378826
rect 121644 378762 121696 378768
rect 120000 377998 120120 378026
rect 120000 377369 120028 377998
rect 119986 377360 120042 377369
rect 119986 377295 120042 377304
rect 118792 354000 118844 354006
rect 118792 353942 118844 353948
rect 118804 353326 118832 353942
rect 118792 353320 118844 353326
rect 118792 353262 118844 353268
rect 118700 311228 118752 311234
rect 118700 311170 118752 311176
rect 118700 297424 118752 297430
rect 118700 297366 118752 297372
rect 117502 275224 117558 275233
rect 117502 275159 117558 275168
rect 118056 272536 118108 272542
rect 118056 272478 118108 272484
rect 116676 253224 116728 253230
rect 116676 253166 116728 253172
rect 117964 233164 118016 233170
rect 117964 233106 118016 233112
rect 117976 232558 118004 233106
rect 117964 232552 118016 232558
rect 117964 232494 118016 232500
rect 116032 222148 116084 222154
rect 116032 222090 116084 222096
rect 116584 222148 116636 222154
rect 116584 222090 116636 222096
rect 116044 84114 116072 222090
rect 117320 181552 117372 181558
rect 117320 181494 117372 181500
rect 116124 180124 116176 180130
rect 116124 180066 116176 180072
rect 116136 91050 116164 180066
rect 116858 142760 116914 142769
rect 116858 142695 116914 142704
rect 116872 137329 116900 142695
rect 116858 137320 116914 137329
rect 116858 137255 116914 137264
rect 116124 91044 116176 91050
rect 116124 90986 116176 90992
rect 117332 89690 117360 181494
rect 117320 89684 117372 89690
rect 117320 89626 117372 89632
rect 117780 89684 117832 89690
rect 117780 89626 117832 89632
rect 117792 88330 117820 89626
rect 117780 88324 117832 88330
rect 117780 88266 117832 88272
rect 117976 85542 118004 232494
rect 118068 227050 118096 272478
rect 118056 227044 118108 227050
rect 118056 226986 118108 226992
rect 117964 85536 118016 85542
rect 117964 85478 118016 85484
rect 116032 84108 116084 84114
rect 116032 84050 116084 84056
rect 116044 84017 116072 84050
rect 116030 84008 116086 84017
rect 116030 83943 116086 83952
rect 117320 32496 117372 32502
rect 117320 32438 117372 32444
rect 117332 16574 117360 32438
rect 109052 16546 109356 16574
rect 110432 16546 110552 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 117332 16546 117636 16574
rect 108396 10396 108448 10402
rect 108396 10338 108448 10344
rect 109328 480 109356 16546
rect 110524 480 110552 16546
rect 111616 7676 111668 7682
rect 111616 7618 111668 7624
rect 111628 480 111656 7618
rect 112364 490 112392 16546
rect 112640 598 112852 626
rect 112640 490 112668 598
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 462 112668 490
rect 112824 480 112852 598
rect 114020 480 114048 16546
rect 114756 490 114784 16546
rect 115032 598 115244 626
rect 115032 490 115060 598
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 462 115060 490
rect 115216 480 115244 598
rect 116412 480 116440 16546
rect 117608 480 117636 16546
rect 118712 3534 118740 297366
rect 118804 234161 118832 353262
rect 120000 351898 120028 377295
rect 121656 376718 121684 378762
rect 121644 376712 121696 376718
rect 121644 376654 121696 376660
rect 119988 351892 120040 351898
rect 119988 351834 120040 351840
rect 121460 327140 121512 327146
rect 121460 327082 121512 327088
rect 120722 307864 120778 307873
rect 120722 307799 120778 307808
rect 120736 274650 120764 307799
rect 120724 274644 120776 274650
rect 120724 274586 120776 274592
rect 120172 273964 120224 273970
rect 120172 273906 120224 273912
rect 119344 270496 119396 270502
rect 119344 270438 119396 270444
rect 118790 234152 118846 234161
rect 118790 234087 118846 234096
rect 118792 184272 118844 184278
rect 118792 184214 118844 184220
rect 118700 3528 118752 3534
rect 118700 3470 118752 3476
rect 118804 480 118832 184214
rect 119356 159390 119384 270438
rect 120078 205048 120134 205057
rect 120078 204983 120134 204992
rect 119344 159384 119396 159390
rect 119344 159326 119396 159332
rect 119356 122806 119384 159326
rect 119344 122800 119396 122806
rect 119344 122742 119396 122748
rect 120092 16574 120120 204983
rect 120184 140729 120212 273906
rect 120724 263628 120776 263634
rect 120724 263570 120776 263576
rect 120736 254590 120764 263570
rect 120724 254584 120776 254590
rect 120724 254526 120776 254532
rect 120170 140720 120226 140729
rect 120170 140655 120226 140664
rect 120184 140049 120212 140655
rect 120170 140040 120226 140049
rect 120170 139975 120226 139984
rect 121472 16574 121500 327082
rect 121550 236736 121606 236745
rect 121550 236671 121606 236680
rect 121564 63442 121592 236671
rect 121656 233170 121684 376654
rect 122116 307057 122144 400182
rect 122852 387569 122880 589970
rect 123496 576842 123524 609962
rect 124864 581120 124916 581126
rect 124864 581062 124916 581068
rect 123484 576836 123536 576842
rect 123484 576778 123536 576784
rect 124876 563718 124904 581062
rect 129660 568546 129688 618258
rect 141976 616888 142028 616894
rect 141976 616830 142028 616836
rect 140688 614236 140740 614242
rect 140688 614178 140740 614184
rect 139308 608660 139360 608666
rect 139308 608602 139360 608608
rect 133788 588600 133840 588606
rect 133788 588542 133840 588548
rect 133800 587926 133828 588542
rect 133788 587920 133840 587926
rect 133788 587862 133840 587868
rect 133800 586514 133828 587862
rect 133708 586486 133828 586514
rect 129648 568540 129700 568546
rect 129648 568482 129700 568488
rect 129004 567860 129056 567866
rect 129004 567802 129056 567808
rect 124864 563712 124916 563718
rect 124864 563654 124916 563660
rect 122930 451344 122986 451353
rect 122930 451279 122986 451288
rect 122838 387560 122894 387569
rect 122838 387495 122894 387504
rect 122944 378729 122972 451279
rect 123024 419416 123076 419422
rect 123024 419358 123076 419364
rect 123036 412758 123064 419358
rect 124876 414730 124904 563654
rect 126888 529236 126940 529242
rect 126888 529178 126940 529184
rect 126244 480276 126296 480282
rect 126244 480218 126296 480224
rect 126256 434722 126284 480218
rect 126244 434716 126296 434722
rect 126244 434658 126296 434664
rect 125600 426488 125652 426494
rect 125600 426430 125652 426436
rect 124864 414724 124916 414730
rect 124864 414666 124916 414672
rect 123024 412752 123076 412758
rect 123024 412694 123076 412700
rect 123036 412622 123064 412694
rect 123024 412616 123076 412622
rect 123024 412558 123076 412564
rect 124864 407176 124916 407182
rect 124864 407118 124916 407124
rect 123482 387560 123538 387569
rect 123482 387495 123538 387504
rect 122930 378720 122986 378729
rect 122930 378655 122986 378664
rect 123496 362914 123524 387495
rect 124876 386374 124904 407118
rect 124956 396092 125008 396098
rect 124956 396034 125008 396040
rect 124864 386368 124916 386374
rect 124864 386310 124916 386316
rect 124220 382968 124272 382974
rect 124220 382910 124272 382916
rect 123484 362908 123536 362914
rect 123484 362850 123536 362856
rect 123576 326392 123628 326398
rect 123576 326334 123628 326340
rect 123482 323776 123538 323785
rect 123482 323711 123538 323720
rect 122102 307048 122158 307057
rect 122102 306983 122158 306992
rect 122838 301608 122894 301617
rect 122838 301543 122894 301552
rect 121644 233164 121696 233170
rect 121644 233106 121696 233112
rect 122104 225684 122156 225690
rect 122104 225626 122156 225632
rect 122116 165753 122144 225626
rect 122102 165744 122158 165753
rect 122102 165679 122158 165688
rect 122116 120086 122144 165679
rect 122104 120080 122156 120086
rect 122104 120022 122156 120028
rect 121552 63436 121604 63442
rect 121552 63378 121604 63384
rect 121564 62801 121592 63378
rect 121550 62792 121606 62801
rect 121550 62727 121606 62736
rect 122852 16574 122880 301543
rect 123496 234025 123524 323711
rect 123482 234016 123538 234025
rect 123482 233951 123538 233960
rect 123484 195356 123536 195362
rect 123484 195298 123536 195304
rect 123496 42090 123524 195298
rect 123588 195294 123616 326334
rect 124232 248414 124260 382910
rect 124968 376689 124996 396034
rect 124954 376680 125010 376689
rect 124954 376615 125010 376624
rect 124862 332616 124918 332625
rect 124862 332551 124918 332560
rect 124232 248386 124352 248414
rect 124324 235958 124352 248386
rect 124312 235952 124364 235958
rect 124312 235894 124364 235900
rect 124218 234016 124274 234025
rect 124218 233951 124274 233960
rect 124128 231192 124180 231198
rect 124128 231134 124180 231140
rect 123576 195288 123628 195294
rect 123576 195230 123628 195236
rect 124140 89690 124168 231134
rect 124128 89684 124180 89690
rect 124128 89626 124180 89632
rect 124140 89282 124168 89626
rect 123576 89276 123628 89282
rect 123576 89218 123628 89224
rect 124128 89276 124180 89282
rect 124128 89218 124180 89224
rect 123588 82822 123616 89218
rect 123576 82816 123628 82822
rect 123576 82758 123628 82764
rect 123484 42084 123536 42090
rect 123484 42026 123536 42032
rect 124232 16574 124260 233951
rect 124324 86970 124352 235894
rect 124312 86964 124364 86970
rect 124312 86906 124364 86912
rect 124876 64190 124904 332551
rect 125612 284306 125640 426430
rect 126900 417246 126928 529178
rect 128268 519648 128320 519654
rect 128268 519590 128320 519596
rect 126244 417240 126296 417246
rect 126244 417182 126296 417188
rect 126888 417240 126940 417246
rect 126888 417182 126940 417188
rect 126256 411262 126284 417182
rect 126900 416838 126928 417182
rect 126888 416832 126940 416838
rect 126888 416774 126940 416780
rect 126244 411256 126296 411262
rect 126244 411198 126296 411204
rect 126244 397520 126296 397526
rect 126244 397462 126296 397468
rect 126256 387802 126284 397462
rect 126244 387796 126296 387802
rect 126244 387738 126296 387744
rect 126244 383036 126296 383042
rect 126244 382978 126296 382984
rect 126256 356726 126284 382978
rect 126244 356720 126296 356726
rect 126244 356662 126296 356668
rect 126888 312656 126940 312662
rect 126888 312598 126940 312604
rect 126900 311914 126928 312598
rect 126336 311908 126388 311914
rect 126336 311850 126388 311856
rect 126888 311908 126940 311914
rect 126888 311850 126940 311856
rect 125600 284300 125652 284306
rect 125600 284242 125652 284248
rect 125612 283626 125640 284242
rect 125600 283620 125652 283626
rect 125600 283562 125652 283568
rect 126244 280900 126296 280906
rect 126244 280842 126296 280848
rect 124956 273964 125008 273970
rect 124956 273906 125008 273912
rect 124968 247042 124996 273906
rect 125048 256760 125100 256766
rect 125048 256702 125100 256708
rect 124956 247036 125008 247042
rect 124956 246978 125008 246984
rect 125060 237386 125088 256702
rect 125140 245676 125192 245682
rect 125140 245618 125192 245624
rect 125048 237380 125100 237386
rect 125048 237322 125100 237328
rect 125152 235793 125180 245618
rect 125138 235784 125194 235793
rect 125138 235719 125194 235728
rect 124864 64184 124916 64190
rect 124864 64126 124916 64132
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 119908 480 119936 3470
rect 120644 490 120672 16546
rect 120920 598 121132 626
rect 120920 490 120948 598
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 462 120948 490
rect 121104 480 121132 598
rect 122300 480 122328 16546
rect 123036 490 123064 16546
rect 123312 598 123524 626
rect 123312 490 123340 598
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 462 123340 490
rect 123496 480 123524 598
rect 124692 480 124720 16546
rect 126256 10334 126284 280842
rect 126348 149734 126376 311850
rect 127624 311228 127676 311234
rect 127624 311170 127676 311176
rect 127636 310554 127664 311170
rect 127624 310548 127676 310554
rect 127624 310490 127676 310496
rect 126428 283620 126480 283626
rect 126428 283562 126480 283568
rect 126336 149728 126388 149734
rect 126336 149670 126388 149676
rect 126440 133210 126468 283562
rect 126520 184204 126572 184210
rect 126520 184146 126572 184152
rect 126428 133204 126480 133210
rect 126428 133146 126480 133152
rect 126336 127628 126388 127634
rect 126336 127570 126388 127576
rect 126348 68338 126376 127570
rect 126532 92546 126560 184146
rect 127636 148374 127664 310490
rect 128280 298081 128308 519590
rect 129016 455394 129044 567802
rect 129660 567194 129688 568482
rect 129660 567166 129780 567194
rect 129648 459604 129700 459610
rect 129648 459546 129700 459552
rect 129004 455388 129056 455394
rect 129004 455330 129056 455336
rect 129002 438968 129058 438977
rect 129002 438903 129058 438912
rect 129016 409154 129044 438903
rect 129004 409148 129056 409154
rect 129004 409090 129056 409096
rect 129004 400240 129056 400246
rect 129004 400182 129056 400188
rect 129016 391921 129044 400182
rect 129002 391912 129058 391921
rect 129002 391847 129058 391856
rect 128360 388476 128412 388482
rect 128360 388418 128412 388424
rect 128372 387870 128400 388418
rect 128360 387864 128412 387870
rect 128360 387806 128412 387812
rect 129004 387864 129056 387870
rect 129004 387806 129056 387812
rect 127806 298072 127862 298081
rect 127806 298007 127862 298016
rect 128266 298072 128322 298081
rect 128266 298007 128322 298016
rect 127820 297401 127848 298007
rect 127806 297392 127862 297401
rect 127806 297327 127862 297336
rect 127716 278112 127768 278118
rect 127716 278054 127768 278060
rect 127728 236609 127756 278054
rect 128360 251184 128412 251190
rect 128360 251126 128412 251132
rect 127714 236600 127770 236609
rect 127714 236535 127770 236544
rect 127716 151836 127768 151842
rect 127716 151778 127768 151784
rect 127624 148368 127676 148374
rect 127624 148310 127676 148316
rect 126612 135924 126664 135930
rect 126612 135866 126664 135872
rect 126624 124137 126652 135866
rect 126610 124128 126666 124137
rect 126610 124063 126666 124072
rect 127728 120737 127756 151778
rect 127714 120728 127770 120737
rect 127714 120663 127770 120672
rect 126520 92540 126572 92546
rect 126520 92482 126572 92488
rect 128372 89758 128400 251126
rect 129016 241505 129044 387806
rect 129660 343670 129688 459546
rect 129752 384985 129780 567166
rect 132408 478984 132460 478990
rect 132408 478926 132460 478932
rect 130384 464364 130436 464370
rect 130384 464306 130436 464312
rect 130396 425066 130424 464306
rect 130384 425060 130436 425066
rect 130384 425002 130436 425008
rect 130384 396772 130436 396778
rect 130384 396714 130436 396720
rect 129738 384976 129794 384985
rect 129738 384911 129794 384920
rect 129752 380186 129780 384911
rect 130396 380798 130424 396714
rect 130384 380792 130436 380798
rect 130384 380734 130436 380740
rect 129740 380180 129792 380186
rect 129740 380122 129792 380128
rect 130384 377460 130436 377466
rect 130384 377402 130436 377408
rect 130396 349110 130424 377402
rect 130384 349104 130436 349110
rect 130384 349046 130436 349052
rect 130660 349104 130712 349110
rect 130660 349046 130712 349052
rect 130384 343732 130436 343738
rect 130384 343674 130436 343680
rect 129096 343664 129148 343670
rect 129096 343606 129148 343612
rect 129648 343664 129700 343670
rect 129648 343606 129700 343612
rect 129108 307834 129136 343606
rect 129096 307828 129148 307834
rect 129096 307770 129148 307776
rect 129002 241496 129058 241505
rect 129002 241431 129058 241440
rect 129002 192536 129058 192545
rect 129002 192471 129058 192480
rect 127624 89752 127676 89758
rect 127624 89694 127676 89700
rect 128360 89752 128412 89758
rect 128360 89694 128412 89700
rect 127636 77246 127664 89694
rect 127624 77240 127676 77246
rect 127624 77182 127676 77188
rect 126336 68332 126388 68338
rect 126336 68274 126388 68280
rect 127636 62082 127664 77182
rect 127624 62076 127676 62082
rect 127624 62018 127676 62024
rect 126244 10328 126296 10334
rect 126244 10270 126296 10276
rect 125876 7608 125928 7614
rect 125876 7550 125928 7556
rect 125888 480 125916 7550
rect 129016 490 129044 192471
rect 129108 153338 129136 307770
rect 129188 298852 129240 298858
rect 129188 298794 129240 298800
rect 129200 193866 129228 298794
rect 129280 260160 129332 260166
rect 129280 260102 129332 260108
rect 129292 251190 129320 260102
rect 129280 251184 129332 251190
rect 129280 251126 129332 251132
rect 129188 193860 129240 193866
rect 129188 193802 129240 193808
rect 129096 153332 129148 153338
rect 129096 153274 129148 153280
rect 129108 145654 129136 153274
rect 129096 145648 129148 145654
rect 129096 145590 129148 145596
rect 129094 127664 129150 127673
rect 129094 127599 129150 127608
rect 129108 15910 129136 127599
rect 129096 15904 129148 15910
rect 129096 15846 129148 15852
rect 130396 6186 130424 343674
rect 130474 334792 130530 334801
rect 130474 334727 130530 334736
rect 130488 24206 130516 334727
rect 130568 249076 130620 249082
rect 130568 249018 130620 249024
rect 130580 102066 130608 249018
rect 130672 231198 130700 349046
rect 131854 328672 131910 328681
rect 131854 328607 131910 328616
rect 131120 291168 131172 291174
rect 131120 291110 131172 291116
rect 131132 290494 131160 291110
rect 131120 290488 131172 290494
rect 131120 290430 131172 290436
rect 131120 251252 131172 251258
rect 131120 251194 131172 251200
rect 130660 231192 130712 231198
rect 130660 231134 130712 231140
rect 130568 102060 130620 102066
rect 130568 102002 130620 102008
rect 130580 101522 130608 102002
rect 130568 101516 130620 101522
rect 130568 101458 130620 101464
rect 131132 99498 131160 251194
rect 131764 193860 131816 193866
rect 131764 193802 131816 193808
rect 131040 99470 131160 99498
rect 131040 99414 131068 99470
rect 131028 99408 131080 99414
rect 131028 99350 131080 99356
rect 131040 71738 131068 99350
rect 131028 71732 131080 71738
rect 131028 71674 131080 71680
rect 130476 24200 130528 24206
rect 130476 24142 130528 24148
rect 131776 24138 131804 193802
rect 131868 188358 131896 328607
rect 132420 290494 132448 478926
rect 133708 473249 133736 586486
rect 134524 578264 134576 578270
rect 134524 578206 134576 578212
rect 133788 481704 133840 481710
rect 133788 481646 133840 481652
rect 133142 473240 133198 473249
rect 133142 473175 133198 473184
rect 133694 473240 133750 473249
rect 133694 473175 133750 473184
rect 133156 472025 133184 473175
rect 133142 472016 133198 472025
rect 133142 471951 133198 471960
rect 132498 434752 132554 434761
rect 132498 434687 132554 434696
rect 132408 290488 132460 290494
rect 132408 290430 132460 290436
rect 132040 251864 132092 251870
rect 132040 251806 132092 251812
rect 132052 251258 132080 251806
rect 132040 251252 132092 251258
rect 132040 251194 132092 251200
rect 131856 188352 131908 188358
rect 131856 188294 131908 188300
rect 131764 24132 131816 24138
rect 131764 24074 131816 24080
rect 132512 16574 132540 434687
rect 133156 427106 133184 471951
rect 133144 427100 133196 427106
rect 133144 427042 133196 427048
rect 133142 331256 133198 331265
rect 133142 331191 133198 331200
rect 132512 16546 133000 16574
rect 130384 6180 130436 6186
rect 130384 6122 130436 6128
rect 129200 598 129412 626
rect 129200 490 129228 598
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129016 462 129228 490
rect 129384 480 129412 598
rect 132972 480 133000 16546
rect 133156 11762 133184 331191
rect 133800 293962 133828 481646
rect 133788 293956 133840 293962
rect 133788 293898 133840 293904
rect 133800 293282 133828 293898
rect 133788 293276 133840 293282
rect 133788 293218 133840 293224
rect 133236 264988 133288 264994
rect 133236 264930 133288 264936
rect 133248 232558 133276 264930
rect 133236 232552 133288 232558
rect 133236 232494 133288 232500
rect 133236 152516 133288 152522
rect 133236 152458 133288 152464
rect 133248 118658 133276 152458
rect 133236 118652 133288 118658
rect 133236 118594 133288 118600
rect 133144 11756 133196 11762
rect 133144 11698 133196 11704
rect 134536 5574 134564 578206
rect 137928 577516 137980 577522
rect 137928 577458 137980 577464
rect 137100 573368 137152 573374
rect 137100 573310 137152 573316
rect 137112 572762 137140 573310
rect 136640 572756 136692 572762
rect 136640 572698 136692 572704
rect 137100 572756 137152 572762
rect 137100 572698 137152 572704
rect 136548 504484 136600 504490
rect 136548 504426 136600 504432
rect 135904 470688 135956 470694
rect 135904 470630 135956 470636
rect 135166 458824 135222 458833
rect 135166 458759 135222 458768
rect 134706 297392 134762 297401
rect 134706 297327 134762 297336
rect 134616 261520 134668 261526
rect 134616 261462 134668 261468
rect 134628 139398 134656 261462
rect 134720 200802 134748 297327
rect 135180 267714 135208 458759
rect 135916 407114 135944 470630
rect 135996 409828 136048 409834
rect 135996 409770 136048 409776
rect 136008 409154 136036 409770
rect 135996 409148 136048 409154
rect 135996 409090 136048 409096
rect 135904 407108 135956 407114
rect 135904 407050 135956 407056
rect 135902 327448 135958 327457
rect 135902 327383 135958 327392
rect 135168 267708 135220 267714
rect 135168 267650 135220 267656
rect 135180 267102 135208 267650
rect 135168 267096 135220 267102
rect 135168 267038 135220 267044
rect 134708 200796 134760 200802
rect 134708 200738 134760 200744
rect 134708 168496 134760 168502
rect 134708 168438 134760 168444
rect 134616 139392 134668 139398
rect 134616 139334 134668 139340
rect 134628 133770 134656 139334
rect 134720 133929 134748 168438
rect 134706 133920 134762 133929
rect 134706 133855 134762 133864
rect 134628 133742 134748 133770
rect 134616 133204 134668 133210
rect 134616 133146 134668 133152
rect 134628 32434 134656 133146
rect 134720 132494 134748 133742
rect 134720 132466 134840 132494
rect 134812 113830 134840 132466
rect 134800 113824 134852 113830
rect 134800 113766 134852 113772
rect 135916 54534 135944 327383
rect 136008 325009 136036 409090
rect 135994 325000 136050 325009
rect 135994 324935 136050 324944
rect 135996 313336 136048 313342
rect 135996 313278 136048 313284
rect 136008 301510 136036 313278
rect 135996 301504 136048 301510
rect 135996 301446 136048 301452
rect 135996 284980 136048 284986
rect 135996 284922 136048 284928
rect 136008 127634 136036 284922
rect 136560 275330 136588 504426
rect 136652 394058 136680 572698
rect 137836 518220 137888 518226
rect 137836 518162 137888 518168
rect 136640 394052 136692 394058
rect 136640 393994 136692 394000
rect 137284 394052 137336 394058
rect 137284 393994 137336 394000
rect 137296 369073 137324 393994
rect 137374 373280 137430 373289
rect 137374 373215 137430 373224
rect 137282 369064 137338 369073
rect 137282 368999 137338 369008
rect 137296 354686 137324 368999
rect 137284 354680 137336 354686
rect 137284 354622 137336 354628
rect 137282 316704 137338 316713
rect 137282 316639 137338 316648
rect 137296 283626 137324 316639
rect 137284 283620 137336 283626
rect 137284 283562 137336 283568
rect 137284 280832 137336 280838
rect 137284 280774 137336 280780
rect 136548 275324 136600 275330
rect 136548 275266 136600 275272
rect 136086 149288 136142 149297
rect 136086 149223 136142 149232
rect 135996 127628 136048 127634
rect 135996 127570 136048 127576
rect 136100 117230 136128 149223
rect 136088 117224 136140 117230
rect 136088 117166 136140 117172
rect 135904 54528 135956 54534
rect 135904 54470 135956 54476
rect 134616 32428 134668 32434
rect 134616 32370 134668 32376
rect 134524 5568 134576 5574
rect 134524 5510 134576 5516
rect 136456 5568 136508 5574
rect 136456 5510 136508 5516
rect 136468 480 136496 5510
rect 137296 2174 137324 280774
rect 137388 238649 137416 373215
rect 137848 372774 137876 518162
rect 137940 396778 137968 577458
rect 138664 441720 138716 441726
rect 138664 441662 138716 441668
rect 138676 430574 138704 441662
rect 138664 430568 138716 430574
rect 138664 430510 138716 430516
rect 137928 396772 137980 396778
rect 137928 396714 137980 396720
rect 139320 382265 139348 608602
rect 140596 466540 140648 466546
rect 140596 466482 140648 466488
rect 139306 382256 139362 382265
rect 139306 382191 139362 382200
rect 139320 381721 139348 382191
rect 139306 381712 139362 381721
rect 139306 381647 139362 381656
rect 138756 380180 138808 380186
rect 138756 380122 138808 380128
rect 137836 372768 137888 372774
rect 137836 372710 137888 372716
rect 137466 333296 137522 333305
rect 137466 333231 137522 333240
rect 137480 280906 137508 333231
rect 138664 324420 138716 324426
rect 138664 324362 138716 324368
rect 137558 284336 137614 284345
rect 137558 284271 137614 284280
rect 137468 280900 137520 280906
rect 137468 280842 137520 280848
rect 137468 264308 137520 264314
rect 137468 264250 137520 264256
rect 137374 238640 137430 238649
rect 137374 238575 137430 238584
rect 137388 237969 137416 238575
rect 137374 237960 137430 237969
rect 137374 237895 137430 237904
rect 137376 188352 137428 188358
rect 137376 188294 137428 188300
rect 137388 21418 137416 188294
rect 137480 184278 137508 264250
rect 137572 216034 137600 284271
rect 137560 216028 137612 216034
rect 137560 215970 137612 215976
rect 138020 211064 138072 211070
rect 138018 211032 138020 211041
rect 138072 211032 138074 211041
rect 138018 210967 138074 210976
rect 137468 184272 137520 184278
rect 137468 184214 137520 184220
rect 137468 154692 137520 154698
rect 137468 154634 137520 154640
rect 137480 134473 137508 154634
rect 137466 134464 137522 134473
rect 137466 134399 137522 134408
rect 138676 49026 138704 324362
rect 138768 211070 138796 380122
rect 140042 311944 140098 311953
rect 140042 311879 140098 311888
rect 138846 272504 138902 272513
rect 138846 272439 138902 272448
rect 138860 245546 138888 272439
rect 138848 245540 138900 245546
rect 138848 245482 138900 245488
rect 138756 211064 138808 211070
rect 138756 211006 138808 211012
rect 140056 195362 140084 311879
rect 140136 283620 140188 283626
rect 140136 283562 140188 283568
rect 140044 195356 140096 195362
rect 140044 195298 140096 195304
rect 140148 182850 140176 283562
rect 140608 281518 140636 466482
rect 140700 331129 140728 614178
rect 141884 520940 141936 520946
rect 141884 520882 141936 520888
rect 141424 476128 141476 476134
rect 141424 476070 141476 476076
rect 141436 430506 141464 476070
rect 141424 430500 141476 430506
rect 141424 430442 141476 430448
rect 141896 409834 141924 520882
rect 141884 409828 141936 409834
rect 141884 409770 141936 409776
rect 141424 408536 141476 408542
rect 141424 408478 141476 408484
rect 141436 375193 141464 408478
rect 141608 392012 141660 392018
rect 141608 391954 141660 391960
rect 141422 375184 141478 375193
rect 141422 375119 141478 375128
rect 141516 372768 141568 372774
rect 141516 372710 141568 372716
rect 141240 372496 141292 372502
rect 141240 372438 141292 372444
rect 141252 371890 141280 372438
rect 141240 371884 141292 371890
rect 141240 371826 141292 371832
rect 140686 331120 140742 331129
rect 140686 331055 140742 331064
rect 140596 281512 140648 281518
rect 140596 281454 140648 281460
rect 141424 268456 141476 268462
rect 141424 268398 141476 268404
rect 140136 182844 140188 182850
rect 140136 182786 140188 182792
rect 140044 181552 140096 181558
rect 140044 181494 140096 181500
rect 138754 160168 138810 160177
rect 138754 160103 138810 160112
rect 138768 121689 138796 160103
rect 138754 121680 138810 121689
rect 138754 121615 138810 121624
rect 140056 53106 140084 181494
rect 140044 53100 140096 53106
rect 140044 53042 140096 53048
rect 138664 49020 138716 49026
rect 138664 48962 138716 48968
rect 141436 43450 141464 268398
rect 141528 262886 141556 372710
rect 141620 360194 141648 391954
rect 141988 385762 142016 616830
rect 142068 615528 142120 615534
rect 142068 615470 142120 615476
rect 141976 385756 142028 385762
rect 141976 385698 142028 385704
rect 142080 371890 142108 615470
rect 143446 610056 143502 610065
rect 143446 609991 143502 610000
rect 143356 594108 143408 594114
rect 143356 594050 143408 594056
rect 143368 593434 143396 594050
rect 143356 593428 143408 593434
rect 143356 593370 143408 593376
rect 143264 507136 143316 507142
rect 143264 507078 143316 507084
rect 142894 475280 142950 475289
rect 142894 475215 142950 475224
rect 142804 460216 142856 460222
rect 142804 460158 142856 460164
rect 142816 419490 142844 460158
rect 142908 457502 142936 475215
rect 142896 457496 142948 457502
rect 142896 457438 142948 457444
rect 142896 444508 142948 444514
rect 142896 444450 142948 444456
rect 142804 419484 142856 419490
rect 142804 419426 142856 419432
rect 142804 412752 142856 412758
rect 142804 412694 142856 412700
rect 142068 371884 142120 371890
rect 142068 371826 142120 371832
rect 141608 360188 141660 360194
rect 141608 360130 141660 360136
rect 142816 358766 142844 412694
rect 142804 358760 142856 358766
rect 142804 358702 142856 358708
rect 142804 337408 142856 337414
rect 142804 337350 142856 337356
rect 141608 336796 141660 336802
rect 141608 336738 141660 336744
rect 141620 263566 141648 336738
rect 142066 307048 142122 307057
rect 142066 306983 142122 306992
rect 142080 295361 142108 306983
rect 141698 295352 141754 295361
rect 141698 295287 141754 295296
rect 142066 295352 142122 295361
rect 142066 295287 142122 295296
rect 141712 267034 141740 295287
rect 141700 267028 141752 267034
rect 141700 266970 141752 266976
rect 141608 263560 141660 263566
rect 141608 263502 141660 263508
rect 141516 262880 141568 262886
rect 141516 262822 141568 262828
rect 141516 261520 141568 261526
rect 141516 261462 141568 261468
rect 141528 127673 141556 261462
rect 141514 127664 141570 127673
rect 141514 127599 141570 127608
rect 141424 43444 141476 43450
rect 141424 43386 141476 43392
rect 137376 21412 137428 21418
rect 137376 21354 137428 21360
rect 142816 10470 142844 337350
rect 142908 287026 142936 444450
rect 143276 406434 143304 507078
rect 143368 475289 143396 593370
rect 143354 475280 143410 475289
rect 143354 475215 143410 475224
rect 143368 474881 143396 475215
rect 143354 474872 143410 474881
rect 143354 474807 143410 474816
rect 143356 445052 143408 445058
rect 143356 444994 143408 445000
rect 143368 444514 143396 444994
rect 143356 444508 143408 444514
rect 143356 444450 143408 444456
rect 143264 406428 143316 406434
rect 143264 406370 143316 406376
rect 142988 392624 143040 392630
rect 142988 392566 143040 392572
rect 143000 364274 143028 392566
rect 142988 364268 143040 364274
rect 142988 364210 143040 364216
rect 143460 341630 143488 609991
rect 144734 605976 144790 605985
rect 144734 605911 144790 605920
rect 144748 605878 144776 605911
rect 144736 605872 144788 605878
rect 144736 605814 144788 605820
rect 144644 537532 144696 537538
rect 144644 537474 144696 537480
rect 144656 535430 144684 537474
rect 143540 535424 143592 535430
rect 143540 535366 143592 535372
rect 144644 535424 144696 535430
rect 144644 535366 144696 535372
rect 143552 400926 143580 535366
rect 144642 449168 144698 449177
rect 144642 449103 144698 449112
rect 143540 400920 143592 400926
rect 143540 400862 143592 400868
rect 144184 394800 144236 394806
rect 144184 394742 144236 394748
rect 144196 361593 144224 394742
rect 144274 378040 144330 378049
rect 144274 377975 144330 377984
rect 144288 373289 144316 377975
rect 144274 373280 144330 373289
rect 144274 373215 144330 373224
rect 144182 361584 144238 361593
rect 144182 361519 144238 361528
rect 143448 341624 143500 341630
rect 143448 341566 143500 341572
rect 143080 335368 143132 335374
rect 143080 335310 143132 335316
rect 142896 287020 142948 287026
rect 142896 286962 142948 286968
rect 142908 286346 142936 286962
rect 142986 286376 143042 286385
rect 142896 286340 142948 286346
rect 142986 286311 143042 286320
rect 142896 286282 142948 286288
rect 142896 263016 142948 263022
rect 142896 262958 142948 262964
rect 142908 44878 142936 262958
rect 143000 178702 143028 286311
rect 143092 256698 143120 335310
rect 144090 331120 144146 331129
rect 144090 331055 144146 331064
rect 144104 329905 144132 331055
rect 143538 329896 143594 329905
rect 143538 329831 143594 329840
rect 144090 329896 144146 329905
rect 144090 329831 144146 329840
rect 143080 256692 143132 256698
rect 143080 256634 143132 256640
rect 142988 178696 143040 178702
rect 142988 178638 143040 178644
rect 142986 162888 143042 162897
rect 142986 162823 143042 162832
rect 143000 128314 143028 162823
rect 142988 128308 143040 128314
rect 142988 128250 143040 128256
rect 143552 51746 143580 329831
rect 144656 325694 144684 449103
rect 144748 378049 144776 605814
rect 144734 378040 144790 378049
rect 144734 377975 144790 377984
rect 144656 325666 144776 325694
rect 144748 310457 144776 325666
rect 144734 310448 144790 310457
rect 144734 310383 144790 310392
rect 144748 309777 144776 310383
rect 144734 309768 144790 309777
rect 144734 309703 144790 309712
rect 144736 305108 144788 305114
rect 144736 305050 144788 305056
rect 144182 272504 144238 272513
rect 144182 272439 144238 272448
rect 144196 108390 144224 272439
rect 144184 108384 144236 108390
rect 144184 108326 144236 108332
rect 143540 51740 143592 51746
rect 143540 51682 143592 51688
rect 142896 44872 142948 44878
rect 142896 44814 142948 44820
rect 142804 10464 142856 10470
rect 142804 10406 142856 10412
rect 144748 3534 144776 305050
rect 144840 257961 144868 622406
rect 151728 619676 151780 619682
rect 151728 619618 151780 619624
rect 148968 600364 149020 600370
rect 148968 600306 149020 600312
rect 148692 583024 148744 583030
rect 148692 582966 148744 582972
rect 146944 569968 146996 569974
rect 146944 569910 146996 569916
rect 146956 545766 146984 569910
rect 146944 545760 146996 545766
rect 146944 545702 146996 545708
rect 146116 542428 146168 542434
rect 146116 542370 146168 542376
rect 146128 423570 146156 542370
rect 146944 538892 146996 538898
rect 146944 538834 146996 538840
rect 146956 522986 146984 538834
rect 146944 522980 146996 522986
rect 146944 522922 146996 522928
rect 147404 522980 147456 522986
rect 147404 522922 147456 522928
rect 146208 509924 146260 509930
rect 146208 509866 146260 509872
rect 146116 423564 146168 423570
rect 146116 423506 146168 423512
rect 146116 420980 146168 420986
rect 146116 420922 146168 420928
rect 145562 311128 145618 311137
rect 145562 311063 145618 311072
rect 144826 257952 144882 257961
rect 144826 257887 144882 257896
rect 145576 189786 145604 311063
rect 145654 283520 145710 283529
rect 145654 283455 145710 283464
rect 145564 189780 145616 189786
rect 145564 189722 145616 189728
rect 145564 188148 145616 188154
rect 145564 188090 145616 188096
rect 145576 22778 145604 188090
rect 145668 181558 145696 283455
rect 146128 250578 146156 420922
rect 146220 333305 146248 509866
rect 147416 474706 147444 522922
rect 147494 516760 147550 516769
rect 147494 516695 147550 516704
rect 146944 474700 146996 474706
rect 146944 474642 146996 474648
rect 147404 474700 147456 474706
rect 147404 474642 147456 474648
rect 146956 473482 146984 474642
rect 146944 473476 146996 473482
rect 146944 473418 146996 473424
rect 146956 433294 146984 473418
rect 146944 433288 146996 433294
rect 146944 433230 146996 433236
rect 147036 412684 147088 412690
rect 147036 412626 147088 412632
rect 146944 404388 146996 404394
rect 146944 404330 146996 404336
rect 146956 373289 146984 404330
rect 147048 399498 147076 412626
rect 147036 399492 147088 399498
rect 147036 399434 147088 399440
rect 147508 390561 147536 516695
rect 147588 515432 147640 515438
rect 147588 515374 147640 515380
rect 147494 390552 147550 390561
rect 147494 390487 147550 390496
rect 147508 389337 147536 390487
rect 147494 389328 147550 389337
rect 147494 389263 147550 389272
rect 147036 385756 147088 385762
rect 147036 385698 147088 385704
rect 146942 373280 146998 373289
rect 146942 373215 146998 373224
rect 146206 333296 146262 333305
rect 146206 333231 146262 333240
rect 146942 309360 146998 309369
rect 146942 309295 146998 309304
rect 146116 250572 146168 250578
rect 146116 250514 146168 250520
rect 145656 181552 145708 181558
rect 145656 181494 145708 181500
rect 145654 151872 145710 151881
rect 145654 151807 145710 151816
rect 145668 117298 145696 151807
rect 145656 117292 145708 117298
rect 145656 117234 145708 117240
rect 146956 50386 146984 309295
rect 147048 271182 147076 385698
rect 147126 317520 147182 317529
rect 147126 317455 147182 317464
rect 147036 271176 147088 271182
rect 147036 271118 147088 271124
rect 147036 256012 147088 256018
rect 147036 255954 147088 255960
rect 147048 193866 147076 255954
rect 147140 253298 147168 317455
rect 147600 308446 147628 515374
rect 148704 438870 148732 582966
rect 148874 523696 148930 523705
rect 148874 523631 148930 523640
rect 148784 478236 148836 478242
rect 148784 478178 148836 478184
rect 147680 438864 147732 438870
rect 147680 438806 147732 438812
rect 148692 438864 148744 438870
rect 148692 438806 148744 438812
rect 147692 438190 147720 438806
rect 147680 438184 147732 438190
rect 147680 438126 147732 438132
rect 148324 416832 148376 416838
rect 148324 416774 148376 416780
rect 148336 381585 148364 416774
rect 148322 381576 148378 381585
rect 148322 381511 148378 381520
rect 148508 331288 148560 331294
rect 148508 331230 148560 331236
rect 147588 308440 147640 308446
rect 147588 308382 147640 308388
rect 148324 298784 148376 298790
rect 148324 298726 148376 298732
rect 147128 253292 147180 253298
rect 147128 253234 147180 253240
rect 147036 193860 147088 193866
rect 147036 193802 147088 193808
rect 146944 50380 146996 50386
rect 146944 50322 146996 50328
rect 145564 22772 145616 22778
rect 145564 22714 145616 22720
rect 148336 7682 148364 298726
rect 148414 285016 148470 285025
rect 148520 284986 148548 331230
rect 148796 316034 148824 478178
rect 148888 338162 148916 523631
rect 148980 376718 149008 600306
rect 150440 596828 150492 596834
rect 150440 596770 150492 596776
rect 150452 596222 150480 596770
rect 150440 596216 150492 596222
rect 150440 596158 150492 596164
rect 150348 586560 150400 586566
rect 150348 586502 150400 586508
rect 150256 543788 150308 543794
rect 150256 543730 150308 543736
rect 150162 455560 150218 455569
rect 150162 455495 150218 455504
rect 149060 398132 149112 398138
rect 149060 398074 149112 398080
rect 149072 398041 149100 398074
rect 149058 398032 149114 398041
rect 149058 397967 149114 397976
rect 149704 387184 149756 387190
rect 149704 387126 149756 387132
rect 148968 376712 149020 376718
rect 148968 376654 149020 376660
rect 148980 369782 149008 376654
rect 149716 376417 149744 387126
rect 149702 376408 149758 376417
rect 149702 376343 149758 376352
rect 148968 369776 149020 369782
rect 148968 369718 149020 369724
rect 148876 338156 148928 338162
rect 148876 338098 148928 338104
rect 149702 333432 149758 333441
rect 149702 333367 149758 333376
rect 148876 316056 148928 316062
rect 148796 316024 148876 316034
rect 148928 316024 148930 316033
rect 148796 316006 148874 316024
rect 148874 315959 148930 315968
rect 148690 313304 148746 313313
rect 148690 313239 148746 313248
rect 148598 285968 148654 285977
rect 148598 285903 148654 285912
rect 148414 284951 148470 284960
rect 148508 284980 148560 284986
rect 148428 188358 148456 284951
rect 148508 284922 148560 284928
rect 148508 255332 148560 255338
rect 148508 255274 148560 255280
rect 148520 228313 148548 255274
rect 148612 243545 148640 285903
rect 148704 283626 148732 313239
rect 148692 283620 148744 283626
rect 148692 283562 148744 283568
rect 148598 243536 148654 243545
rect 148598 243471 148654 243480
rect 148506 228304 148562 228313
rect 148506 228239 148562 228248
rect 148508 193860 148560 193866
rect 148508 193802 148560 193808
rect 148416 188352 148468 188358
rect 148416 188294 148468 188300
rect 148520 133210 148548 193802
rect 148598 153776 148654 153785
rect 148598 153711 148654 153720
rect 148508 133204 148560 133210
rect 148508 133146 148560 133152
rect 148612 132394 148640 153711
rect 148692 133204 148744 133210
rect 148692 133146 148744 133152
rect 148600 132388 148652 132394
rect 148600 132330 148652 132336
rect 148416 131164 148468 131170
rect 148416 131106 148468 131112
rect 148428 37942 148456 131106
rect 148704 125594 148732 133146
rect 148692 125588 148744 125594
rect 148692 125530 148744 125536
rect 148508 101516 148560 101522
rect 148508 101458 148560 101464
rect 148520 77246 148548 101458
rect 148508 77240 148560 77246
rect 148508 77182 148560 77188
rect 149716 47598 149744 333367
rect 150176 320142 150204 455495
rect 150268 383722 150296 543730
rect 150360 398041 150388 586502
rect 150346 398032 150402 398041
rect 150346 397967 150402 397976
rect 150452 383790 150480 596158
rect 151084 574116 151136 574122
rect 151084 574058 151136 574064
rect 151096 535401 151124 574058
rect 151082 535392 151138 535401
rect 151082 535327 151138 535336
rect 151084 472048 151136 472054
rect 151084 471990 151136 471996
rect 151096 449274 151124 471990
rect 151634 450120 151690 450129
rect 151634 450055 151690 450064
rect 151084 449268 151136 449274
rect 151084 449210 151136 449216
rect 151084 423564 151136 423570
rect 151084 423506 151136 423512
rect 151096 422346 151124 423506
rect 151084 422340 151136 422346
rect 151084 422282 151136 422288
rect 150440 383784 150492 383790
rect 150440 383726 150492 383732
rect 150256 383716 150308 383722
rect 150256 383658 150308 383664
rect 150452 383654 150480 383726
rect 150360 383626 150480 383654
rect 150360 371142 150388 383626
rect 151096 382226 151124 422282
rect 151176 403028 151228 403034
rect 151176 402970 151228 402976
rect 150808 382220 150860 382226
rect 150808 382162 150860 382168
rect 151084 382220 151136 382226
rect 151084 382162 151136 382168
rect 150820 381546 150848 382162
rect 150808 381540 150860 381546
rect 150808 381482 150860 381488
rect 150348 371136 150400 371142
rect 150348 371078 150400 371084
rect 151188 369782 151216 402970
rect 151176 369776 151228 369782
rect 151176 369718 151228 369724
rect 151266 347848 151322 347857
rect 151266 347783 151322 347792
rect 150440 338156 150492 338162
rect 150440 338098 150492 338104
rect 150164 320136 150216 320142
rect 150164 320078 150216 320084
rect 149796 316056 149848 316062
rect 149796 315998 149848 316004
rect 149808 213926 149836 315998
rect 149888 259480 149940 259486
rect 149888 259422 149940 259428
rect 149900 227730 149928 259422
rect 149888 227724 149940 227730
rect 149888 227666 149940 227672
rect 149796 213920 149848 213926
rect 149796 213862 149848 213868
rect 149796 200796 149848 200802
rect 149796 200738 149848 200744
rect 149808 109750 149836 200738
rect 150452 113801 150480 338098
rect 151176 323060 151228 323066
rect 151176 323002 151228 323008
rect 151084 303680 151136 303686
rect 151084 303622 151136 303628
rect 150532 277296 150584 277302
rect 150532 277238 150584 277244
rect 150544 175234 150572 277238
rect 150532 175228 150584 175234
rect 150532 175170 150584 175176
rect 150544 174554 150572 175170
rect 150532 174548 150584 174554
rect 150532 174490 150584 174496
rect 150438 113792 150494 113801
rect 150438 113727 150494 113736
rect 149796 109744 149848 109750
rect 149796 109686 149848 109692
rect 149704 47592 149756 47598
rect 149704 47534 149756 47540
rect 148416 37936 148468 37942
rect 148416 37878 148468 37884
rect 151096 26926 151124 303622
rect 151188 243574 151216 323002
rect 151280 277302 151308 347783
rect 151648 334626 151676 450055
rect 151740 425066 151768 619618
rect 178776 618384 178828 618390
rect 178776 618326 178828 618332
rect 177488 616956 177540 616962
rect 177488 616898 177540 616904
rect 152556 614168 152608 614174
rect 152556 614110 152608 614116
rect 152462 533352 152518 533361
rect 152462 533287 152518 533296
rect 151728 425060 151780 425066
rect 151728 425002 151780 425008
rect 151636 334620 151688 334626
rect 151636 334562 151688 334568
rect 151268 277296 151320 277302
rect 151268 277238 151320 277244
rect 151176 243568 151228 243574
rect 151176 243510 151228 243516
rect 151174 241632 151230 241641
rect 151174 241567 151230 241576
rect 151188 220153 151216 241567
rect 151174 220144 151230 220153
rect 151174 220079 151230 220088
rect 151174 144936 151230 144945
rect 151174 144871 151230 144880
rect 151188 121446 151216 144871
rect 151176 121440 151228 121446
rect 151176 121382 151228 121388
rect 151174 98288 151230 98297
rect 151174 98223 151230 98232
rect 151188 86737 151216 98223
rect 151174 86728 151230 86737
rect 151174 86663 151230 86672
rect 151084 26920 151136 26926
rect 151084 26862 151136 26868
rect 148324 7676 148376 7682
rect 148324 7618 148376 7624
rect 152476 3670 152504 533287
rect 152568 420986 152596 614110
rect 153844 612876 153896 612882
rect 153844 612818 153896 612824
rect 153016 514072 153068 514078
rect 153016 514014 153068 514020
rect 152924 421592 152976 421598
rect 152924 421534 152976 421540
rect 152556 420980 152608 420986
rect 152556 420922 152608 420928
rect 152738 321600 152794 321609
rect 152738 321535 152794 321544
rect 152554 318200 152610 318209
rect 152554 318135 152610 318144
rect 152568 317529 152596 318135
rect 152554 317520 152610 317529
rect 152554 317455 152610 317464
rect 152646 301200 152702 301209
rect 152646 301135 152702 301144
rect 152556 262948 152608 262954
rect 152556 262890 152608 262896
rect 152568 4826 152596 262890
rect 152660 196654 152688 301135
rect 152752 263022 152780 321535
rect 152936 318209 152964 421534
rect 153028 405686 153056 514014
rect 153856 456113 153884 612818
rect 173806 611416 173862 611425
rect 173806 611351 173862 611360
rect 160742 608696 160798 608705
rect 160742 608631 160798 608640
rect 155866 607336 155922 607345
rect 155866 607271 155922 607280
rect 153934 570616 153990 570625
rect 153934 570551 153990 570560
rect 153948 458153 153976 570551
rect 155776 541680 155828 541686
rect 155776 541622 155828 541628
rect 154488 494760 154540 494766
rect 154488 494702 154540 494708
rect 153934 458144 153990 458153
rect 153934 458079 153990 458088
rect 154028 457496 154080 457502
rect 154028 457438 154080 457444
rect 153842 456104 153898 456113
rect 153842 456039 153898 456048
rect 153108 420980 153160 420986
rect 153108 420922 153160 420928
rect 153120 420889 153148 420922
rect 153106 420880 153162 420889
rect 153106 420815 153162 420824
rect 153108 417444 153160 417450
rect 153108 417386 153160 417392
rect 153016 405680 153068 405686
rect 153016 405622 153068 405628
rect 153016 396024 153068 396030
rect 153016 395966 153068 395972
rect 153028 394738 153056 395966
rect 153016 394732 153068 394738
rect 153016 394674 153068 394680
rect 153028 364274 153056 394674
rect 153016 364268 153068 364274
rect 153016 364210 153068 364216
rect 152922 318200 152978 318209
rect 152922 318135 152978 318144
rect 153120 289785 153148 417386
rect 153856 409154 153884 456039
rect 154040 429146 154068 457438
rect 154396 454708 154448 454714
rect 154396 454650 154448 454656
rect 154408 429146 154436 454650
rect 154028 429140 154080 429146
rect 154028 429082 154080 429088
rect 154396 429140 154448 429146
rect 154396 429082 154448 429088
rect 154028 414044 154080 414050
rect 154028 413986 154080 413992
rect 153844 409148 153896 409154
rect 153844 409090 153896 409096
rect 153936 383716 153988 383722
rect 153936 383658 153988 383664
rect 153198 335472 153254 335481
rect 153198 335407 153254 335416
rect 153212 330546 153240 335407
rect 153200 330540 153252 330546
rect 153200 330482 153252 330488
rect 153290 326360 153346 326369
rect 153290 326295 153346 326304
rect 153304 322386 153332 326295
rect 153292 322380 153344 322386
rect 153292 322322 153344 322328
rect 153844 321632 153896 321638
rect 153844 321574 153896 321580
rect 153106 289776 153162 289785
rect 153106 289711 153162 289720
rect 153120 289105 153148 289711
rect 153106 289096 153162 289105
rect 153106 289031 153162 289040
rect 152832 274712 152884 274718
rect 152832 274654 152884 274660
rect 152740 263016 152792 263022
rect 152740 262958 152792 262964
rect 152844 240786 152872 274654
rect 152832 240780 152884 240786
rect 152832 240722 152884 240728
rect 152648 196648 152700 196654
rect 152648 196590 152700 196596
rect 152648 161560 152700 161566
rect 152648 161502 152700 161508
rect 152660 124166 152688 161502
rect 153856 131170 153884 321574
rect 153948 265674 153976 383658
rect 154040 380866 154068 413986
rect 154396 410576 154448 410582
rect 154396 410518 154448 410524
rect 154408 409902 154436 410518
rect 154396 409896 154448 409902
rect 154396 409838 154448 409844
rect 154304 404320 154356 404326
rect 154304 404262 154356 404268
rect 154316 403102 154344 404262
rect 154304 403096 154356 403102
rect 154304 403038 154356 403044
rect 154316 384441 154344 403038
rect 154302 384432 154358 384441
rect 154302 384367 154358 384376
rect 154028 380860 154080 380866
rect 154028 380802 154080 380808
rect 154408 368393 154436 409838
rect 154394 368384 154450 368393
rect 154394 368319 154450 368328
rect 154500 343641 154528 494702
rect 155684 484492 155736 484498
rect 155684 484434 155736 484440
rect 155592 433288 155644 433294
rect 155592 433230 155644 433236
rect 155604 432614 155632 433230
rect 155592 432608 155644 432614
rect 155592 432550 155644 432556
rect 155604 402974 155632 432550
rect 155696 417450 155724 484434
rect 155788 433294 155816 541622
rect 155776 433288 155828 433294
rect 155776 433230 155828 433236
rect 155776 429888 155828 429894
rect 155776 429830 155828 429836
rect 155684 417444 155736 417450
rect 155684 417386 155736 417392
rect 155604 402946 155724 402974
rect 155222 398984 155278 398993
rect 155222 398919 155278 398928
rect 155236 361554 155264 398919
rect 155696 387705 155724 402946
rect 155682 387696 155738 387705
rect 155682 387631 155738 387640
rect 155696 387025 155724 387631
rect 155682 387016 155738 387025
rect 155682 386951 155738 386960
rect 155224 361548 155276 361554
rect 155224 361490 155276 361496
rect 154486 343632 154542 343641
rect 154486 343567 154542 343576
rect 154500 342961 154528 343567
rect 154486 342952 154542 342961
rect 154486 342887 154542 342896
rect 155408 341624 155460 341630
rect 155408 341566 155460 341572
rect 154026 338736 154082 338745
rect 154026 338671 154082 338680
rect 154040 333266 154068 338671
rect 154028 333260 154080 333266
rect 154028 333202 154080 333208
rect 154486 330576 154542 330585
rect 154486 330511 154542 330520
rect 154500 326398 154528 330511
rect 154488 326392 154540 326398
rect 154488 326334 154540 326340
rect 154488 324352 154540 324358
rect 154488 324294 154540 324300
rect 154500 320890 154528 324294
rect 155316 322992 155368 322998
rect 155316 322934 155368 322940
rect 154488 320884 154540 320890
rect 154488 320826 154540 320832
rect 154118 319424 154174 319433
rect 154118 319359 154174 319368
rect 154028 315376 154080 315382
rect 154028 315318 154080 315324
rect 154040 277370 154068 315318
rect 154132 315314 154160 319359
rect 154120 315308 154172 315314
rect 154120 315250 154172 315256
rect 155222 314800 155278 314809
rect 155222 314735 155278 314744
rect 154028 277364 154080 277370
rect 154028 277306 154080 277312
rect 154028 269884 154080 269890
rect 154028 269826 154080 269832
rect 153936 265668 153988 265674
rect 153936 265610 153988 265616
rect 153936 264240 153988 264246
rect 153936 264182 153988 264188
rect 153948 231198 153976 264182
rect 153936 231192 153988 231198
rect 153936 231134 153988 231140
rect 154040 188154 154068 269826
rect 154028 188148 154080 188154
rect 154028 188090 154080 188096
rect 154028 173936 154080 173942
rect 154028 173878 154080 173884
rect 154040 170406 154068 173878
rect 154028 170400 154080 170406
rect 154028 170342 154080 170348
rect 154396 169856 154448 169862
rect 154396 169798 154448 169804
rect 154408 163606 154436 169798
rect 154488 164960 154540 164966
rect 154488 164902 154540 164908
rect 154396 163600 154448 163606
rect 154396 163542 154448 163548
rect 154500 162761 154528 164902
rect 154486 162752 154542 162761
rect 154486 162687 154542 162696
rect 154486 158808 154542 158817
rect 154486 158743 154542 158752
rect 153934 154728 153990 154737
rect 153934 154663 153990 154672
rect 153948 145625 153976 154663
rect 154500 152590 154528 158743
rect 154488 152584 154540 152590
rect 154488 152526 154540 152532
rect 153934 145616 153990 145625
rect 153934 145551 153990 145560
rect 153936 143608 153988 143614
rect 153936 143550 153988 143556
rect 153844 131164 153896 131170
rect 153844 131106 153896 131112
rect 152648 124160 152700 124166
rect 152648 124102 152700 124108
rect 153948 111790 153976 143550
rect 153936 111784 153988 111790
rect 153936 111726 153988 111732
rect 153844 109744 153896 109750
rect 153844 109686 153896 109692
rect 153856 81394 153884 109686
rect 153844 81388 153896 81394
rect 153844 81330 153896 81336
rect 155236 13122 155264 314735
rect 155328 280090 155356 322934
rect 155420 315518 155448 341566
rect 155408 315512 155460 315518
rect 155408 315454 155460 315460
rect 155316 280084 155368 280090
rect 155316 280026 155368 280032
rect 155316 276684 155368 276690
rect 155316 276626 155368 276632
rect 155328 39370 155356 276626
rect 155500 276072 155552 276078
rect 155500 276014 155552 276020
rect 155406 261488 155462 261497
rect 155406 261423 155462 261432
rect 155420 217326 155448 261423
rect 155512 249082 155540 276014
rect 155788 275398 155816 429830
rect 155880 360126 155908 607271
rect 159364 594856 159416 594862
rect 159364 594798 159416 594804
rect 157156 583840 157208 583846
rect 157156 583782 157208 583788
rect 157064 492040 157116 492046
rect 157064 491982 157116 491988
rect 156604 457428 156656 457434
rect 156604 457370 156656 457376
rect 156616 396030 156644 457370
rect 156604 396024 156656 396030
rect 156604 395966 156656 395972
rect 156696 389836 156748 389842
rect 156696 389778 156748 389784
rect 156602 367024 156658 367033
rect 156602 366959 156658 366968
rect 156052 360664 156104 360670
rect 156052 360606 156104 360612
rect 155868 360120 155920 360126
rect 155868 360062 155920 360068
rect 155868 356720 155920 356726
rect 155868 356662 155920 356668
rect 155880 332602 155908 356662
rect 155880 332574 156000 332602
rect 155776 275392 155828 275398
rect 155776 275334 155828 275340
rect 155500 249076 155552 249082
rect 155500 249018 155552 249024
rect 155972 245614 156000 332574
rect 156064 278050 156092 360606
rect 156616 307057 156644 366959
rect 156708 361486 156736 389778
rect 156696 361480 156748 361486
rect 156696 361422 156748 361428
rect 156708 360670 156736 361422
rect 156696 360664 156748 360670
rect 156696 360606 156748 360612
rect 157076 322318 157104 491982
rect 157168 389162 157196 583782
rect 158720 583772 158772 583778
rect 158720 583714 158772 583720
rect 158536 581664 158588 581670
rect 158536 581606 158588 581612
rect 157248 570648 157300 570654
rect 157248 570590 157300 570596
rect 157156 389156 157208 389162
rect 157156 389098 157208 389104
rect 157260 367033 157288 570590
rect 158444 465724 158496 465730
rect 158444 465666 158496 465672
rect 157984 403028 158036 403034
rect 157984 402970 158036 402976
rect 157340 379500 157392 379506
rect 157340 379442 157392 379448
rect 157352 379030 157380 379442
rect 157996 379030 158024 402970
rect 158076 385076 158128 385082
rect 158076 385018 158128 385024
rect 157340 379024 157392 379030
rect 157340 378966 157392 378972
rect 157984 379024 158036 379030
rect 157984 378966 158036 378972
rect 157246 367024 157302 367033
rect 157246 366959 157302 366968
rect 157064 322312 157116 322318
rect 157064 322254 157116 322260
rect 157076 321638 157104 322254
rect 157064 321632 157116 321638
rect 157064 321574 157116 321580
rect 156602 307048 156658 307057
rect 156602 306983 156658 306992
rect 156604 294704 156656 294710
rect 156604 294646 156656 294652
rect 156616 284306 156644 294646
rect 157248 292528 157300 292534
rect 157248 292470 157300 292476
rect 157260 291242 157288 292470
rect 157248 291236 157300 291242
rect 157248 291178 157300 291184
rect 156604 284300 156656 284306
rect 156604 284242 156656 284248
rect 156052 278044 156104 278050
rect 156052 277986 156104 277992
rect 156604 274032 156656 274038
rect 156604 273974 156656 273980
rect 155960 245608 156012 245614
rect 155960 245550 156012 245556
rect 155972 244934 156000 245550
rect 155960 244928 156012 244934
rect 155960 244870 156012 244876
rect 155408 217320 155460 217326
rect 155408 217262 155460 217268
rect 155866 136504 155922 136513
rect 155866 136439 155922 136448
rect 155880 135289 155908 136439
rect 155866 135280 155922 135289
rect 155866 135215 155922 135224
rect 155880 122806 155908 135215
rect 155868 122800 155920 122806
rect 155868 122742 155920 122748
rect 155316 39364 155368 39370
rect 155316 39306 155368 39312
rect 156616 32502 156644 273974
rect 156694 240816 156750 240825
rect 156694 240751 156750 240760
rect 156708 215286 156736 240751
rect 156696 215280 156748 215286
rect 156696 215222 156748 215228
rect 156708 136513 156736 215222
rect 157260 160206 157288 291178
rect 157352 243370 157380 378966
rect 158088 371210 158116 385018
rect 158076 371204 158128 371210
rect 158076 371146 158128 371152
rect 158076 331900 158128 331906
rect 158076 331842 158128 331848
rect 157984 272604 158036 272610
rect 157984 272546 158036 272552
rect 157340 243364 157392 243370
rect 157340 243306 157392 243312
rect 157352 242962 157380 243306
rect 157340 242956 157392 242962
rect 157340 242898 157392 242904
rect 156788 160200 156840 160206
rect 156788 160142 156840 160148
rect 157248 160200 157300 160206
rect 157248 160142 157300 160148
rect 156694 136504 156750 136513
rect 156694 136439 156750 136448
rect 156800 134026 156828 160142
rect 156788 134020 156840 134026
rect 156788 133962 156840 133968
rect 156604 32496 156656 32502
rect 156604 32438 156656 32444
rect 157996 31074 158024 272546
rect 158088 160721 158116 331842
rect 158456 331809 158484 465666
rect 158548 392630 158576 581606
rect 158732 578950 158760 583714
rect 158720 578944 158772 578950
rect 158720 578886 158772 578892
rect 158626 565040 158682 565049
rect 158626 564975 158682 564984
rect 158536 392624 158588 392630
rect 158536 392566 158588 392572
rect 158442 331800 158498 331809
rect 158442 331735 158498 331744
rect 158640 266393 158668 564975
rect 158720 534064 158772 534070
rect 158720 534006 158772 534012
rect 158732 533594 158760 534006
rect 158720 533588 158772 533594
rect 158720 533530 158772 533536
rect 158732 404326 158760 533530
rect 158812 451920 158864 451926
rect 158810 451888 158812 451897
rect 158864 451888 158866 451897
rect 158810 451823 158866 451832
rect 158720 404320 158772 404326
rect 158720 404262 158772 404268
rect 159376 394058 159404 594798
rect 159916 578944 159968 578950
rect 159916 578886 159968 578892
rect 159456 554804 159508 554810
rect 159456 554746 159508 554752
rect 159468 533594 159496 554746
rect 159456 533588 159508 533594
rect 159456 533530 159508 533536
rect 159928 451897 159956 578886
rect 160756 558890 160784 608631
rect 169024 604512 169076 604518
rect 169024 604454 169076 604460
rect 165526 600536 165582 600545
rect 165526 600471 165582 600480
rect 161388 597576 161440 597582
rect 161388 597518 161440 597524
rect 160744 558884 160796 558890
rect 160744 558826 160796 558832
rect 160100 549908 160152 549914
rect 160100 549850 160152 549856
rect 160112 549302 160140 549850
rect 160100 549296 160152 549302
rect 160100 549238 160152 549244
rect 160744 549296 160796 549302
rect 160744 549238 160796 549244
rect 160008 486464 160060 486470
rect 160008 486406 160060 486412
rect 159914 451888 159970 451897
rect 159914 451823 159970 451832
rect 159914 443048 159970 443057
rect 159914 442983 159970 442992
rect 159364 394052 159416 394058
rect 159364 393994 159416 394000
rect 158720 381540 158772 381546
rect 158720 381482 158772 381488
rect 158732 311166 158760 381482
rect 159928 316713 159956 442983
rect 159914 316704 159970 316713
rect 159914 316639 159970 316648
rect 159362 312080 159418 312089
rect 159362 312015 159418 312024
rect 158720 311160 158772 311166
rect 158720 311102 158772 311108
rect 159376 298858 159404 312015
rect 159364 298852 159416 298858
rect 159364 298794 159416 298800
rect 159364 293276 159416 293282
rect 159364 293218 159416 293224
rect 158626 266384 158682 266393
rect 158626 266319 158682 266328
rect 158720 250572 158772 250578
rect 158720 250514 158772 250520
rect 158168 243364 158220 243370
rect 158168 243306 158220 243312
rect 158180 227662 158208 243306
rect 158732 235929 158760 250514
rect 158718 235920 158774 235929
rect 158718 235855 158774 235864
rect 158732 234705 158760 235855
rect 158718 234696 158774 234705
rect 158718 234631 158774 234640
rect 158168 227656 158220 227662
rect 158168 227598 158220 227604
rect 158180 226370 158208 227598
rect 158168 226364 158220 226370
rect 158168 226306 158220 226312
rect 158628 226364 158680 226370
rect 158628 226306 158680 226312
rect 158074 160712 158130 160721
rect 158074 160647 158130 160656
rect 158088 126954 158116 160647
rect 158076 126948 158128 126954
rect 158076 126890 158128 126896
rect 158640 101454 158668 226306
rect 159376 143449 159404 293218
rect 160020 289134 160048 486406
rect 160756 468518 160784 549238
rect 161204 500268 161256 500274
rect 161204 500210 161256 500216
rect 160744 468512 160796 468518
rect 160744 468454 160796 468460
rect 160744 458312 160796 458318
rect 160744 458254 160796 458260
rect 160756 445738 160784 458254
rect 160100 445732 160152 445738
rect 160100 445674 160152 445680
rect 160744 445732 160796 445738
rect 160744 445674 160796 445680
rect 160112 444446 160140 445674
rect 160100 444440 160152 444446
rect 160100 444382 160152 444388
rect 160112 294642 160140 444382
rect 161216 391950 161244 500210
rect 161294 471200 161350 471209
rect 161294 471135 161350 471144
rect 161204 391944 161256 391950
rect 161204 391886 161256 391892
rect 161216 391241 161244 391886
rect 161202 391232 161258 391241
rect 161202 391167 161258 391176
rect 160374 390416 160430 390425
rect 160374 390351 160430 390360
rect 160388 389201 160416 390351
rect 160374 389192 160430 389201
rect 160374 389127 160430 389136
rect 160192 334620 160244 334626
rect 160192 334562 160244 334568
rect 160204 334014 160232 334562
rect 160192 334008 160244 334014
rect 160192 333950 160244 333956
rect 160744 334008 160796 334014
rect 160744 333950 160796 333956
rect 160190 306912 160246 306921
rect 160190 306847 160246 306856
rect 160204 304298 160232 306847
rect 160192 304292 160244 304298
rect 160192 304234 160244 304240
rect 160100 294636 160152 294642
rect 160100 294578 160152 294584
rect 159456 289128 159508 289134
rect 159456 289070 159508 289076
rect 160008 289128 160060 289134
rect 160008 289070 160060 289076
rect 158718 143440 158774 143449
rect 158718 143375 158774 143384
rect 159362 143440 159418 143449
rect 159362 143375 159418 143384
rect 158732 142769 158760 143375
rect 158718 142760 158774 142769
rect 158718 142695 158774 142704
rect 159468 141438 159496 289070
rect 159638 234696 159694 234705
rect 159638 234631 159694 234640
rect 159548 220176 159600 220182
rect 159548 220118 159600 220124
rect 159560 219434 159588 220118
rect 159548 219428 159600 219434
rect 159548 219370 159600 219376
rect 159560 153241 159588 219370
rect 159652 204241 159680 234631
rect 159638 204232 159694 204241
rect 159638 204167 159694 204176
rect 159546 153232 159602 153241
rect 159546 153167 159602 153176
rect 159456 141432 159508 141438
rect 159456 141374 159508 141380
rect 159362 139496 159418 139505
rect 159362 139431 159418 139440
rect 159376 111897 159404 139431
rect 159560 121446 159588 153167
rect 159652 139505 159680 204167
rect 160756 143313 160784 333950
rect 160928 326392 160980 326398
rect 161308 326369 161336 471135
rect 161400 402354 161428 597518
rect 165540 595474 165568 600471
rect 165528 595468 165580 595474
rect 165528 595410 165580 595416
rect 165540 594930 165568 595410
rect 165528 594924 165580 594930
rect 165528 594866 165580 594872
rect 166264 594924 166316 594930
rect 166264 594866 166316 594872
rect 164884 592136 164936 592142
rect 164884 592078 164936 592084
rect 163504 590708 163556 590714
rect 163504 590650 163556 590656
rect 161480 579760 161532 579766
rect 161480 579702 161532 579708
rect 161492 410582 161520 579702
rect 162768 558204 162820 558210
rect 162768 558146 162820 558152
rect 162216 551336 162268 551342
rect 162216 551278 162268 551284
rect 162228 550662 162256 551278
rect 161572 550656 161624 550662
rect 161572 550598 161624 550604
rect 162216 550656 162268 550662
rect 162216 550598 162268 550604
rect 161480 410576 161532 410582
rect 161480 410518 161532 410524
rect 161480 405680 161532 405686
rect 161480 405622 161532 405628
rect 161388 402348 161440 402354
rect 161388 402290 161440 402296
rect 161386 389192 161442 389201
rect 161386 389127 161442 389136
rect 161400 371210 161428 389127
rect 161492 376553 161520 405622
rect 161584 390425 161612 550598
rect 162676 498840 162728 498846
rect 162676 498782 162728 498788
rect 162688 397322 162716 498782
rect 162780 404326 162808 558146
rect 162860 539640 162912 539646
rect 162860 539582 162912 539588
rect 162872 534478 162900 539582
rect 162860 534472 162912 534478
rect 162860 534414 162912 534420
rect 163516 457434 163544 590650
rect 163596 572824 163648 572830
rect 163596 572766 163648 572772
rect 163504 457428 163556 457434
rect 163504 457370 163556 457376
rect 163608 443057 163636 572766
rect 163872 535424 163924 535430
rect 163872 535366 163924 535372
rect 163884 534478 163912 535366
rect 163872 534472 163924 534478
rect 163872 534414 163924 534420
rect 163594 443048 163650 443057
rect 163594 442983 163650 442992
rect 162768 404320 162820 404326
rect 162768 404262 162820 404268
rect 162780 403034 162808 404262
rect 162768 403028 162820 403034
rect 162768 402970 162820 402976
rect 162124 397316 162176 397322
rect 162124 397258 162176 397264
rect 162676 397316 162728 397322
rect 162676 397258 162728 397264
rect 162136 396098 162164 397258
rect 162124 396092 162176 396098
rect 162124 396034 162176 396040
rect 161570 390416 161626 390425
rect 161570 390351 161626 390360
rect 161572 389156 161624 389162
rect 161572 389098 161624 389104
rect 161478 376544 161534 376553
rect 161478 376479 161534 376488
rect 161584 373930 161612 389098
rect 162136 385082 162164 396034
rect 162216 396024 162268 396030
rect 162216 395966 162268 395972
rect 162124 385076 162176 385082
rect 162124 385018 162176 385024
rect 162122 376544 162178 376553
rect 162122 376479 162178 376488
rect 161572 373924 161624 373930
rect 161572 373866 161624 373872
rect 161388 371204 161440 371210
rect 161388 371146 161440 371152
rect 161480 366988 161532 366994
rect 161480 366930 161532 366936
rect 160928 326334 160980 326340
rect 161294 326360 161350 326369
rect 160836 281648 160888 281654
rect 160836 281590 160888 281596
rect 160848 266354 160876 281590
rect 160836 266348 160888 266354
rect 160836 266290 160888 266296
rect 160836 263628 160888 263634
rect 160836 263570 160888 263576
rect 160742 143304 160798 143313
rect 160742 143239 160798 143248
rect 159638 139496 159694 139505
rect 159638 139431 159694 139440
rect 159548 121440 159600 121446
rect 159548 121382 159600 121388
rect 159362 111888 159418 111897
rect 159362 111823 159418 111832
rect 160744 111852 160796 111858
rect 160744 111794 160796 111800
rect 159364 111104 159416 111110
rect 159364 111046 159416 111052
rect 158628 101448 158680 101454
rect 158628 101390 158680 101396
rect 159376 85474 159404 111046
rect 159364 85468 159416 85474
rect 159364 85410 159416 85416
rect 160756 70310 160784 111794
rect 160848 73846 160876 263570
rect 160940 146985 160968 326334
rect 161294 326295 161350 326304
rect 161492 245682 161520 366930
rect 162136 327321 162164 376479
rect 162228 366994 162256 395966
rect 163884 393990 163912 534414
rect 164056 474768 164108 474774
rect 164056 474710 164108 474716
rect 163964 442264 164016 442270
rect 163964 442206 164016 442212
rect 163976 441658 164004 442206
rect 163964 441652 164016 441658
rect 163964 441594 164016 441600
rect 163872 393984 163924 393990
rect 163872 393926 163924 393932
rect 163870 384976 163926 384985
rect 163870 384911 163926 384920
rect 163884 384305 163912 384911
rect 163870 384296 163926 384305
rect 163870 384231 163926 384240
rect 162768 373924 162820 373930
rect 162768 373866 162820 373872
rect 162216 366988 162268 366994
rect 162216 366930 162268 366936
rect 162122 327312 162178 327321
rect 162122 327247 162178 327256
rect 162136 323785 162164 327247
rect 162122 323776 162178 323785
rect 162122 323711 162178 323720
rect 162122 317520 162178 317529
rect 162122 317455 162178 317464
rect 162136 280838 162164 317455
rect 162216 315512 162268 315518
rect 162216 315454 162268 315460
rect 162228 299470 162256 315454
rect 162216 299464 162268 299470
rect 162216 299406 162268 299412
rect 162124 280832 162176 280838
rect 162124 280774 162176 280780
rect 162122 253872 162178 253881
rect 162122 253807 162178 253816
rect 161480 245676 161532 245682
rect 161480 245618 161532 245624
rect 161480 233232 161532 233238
rect 161480 233174 161532 233180
rect 160926 146976 160982 146985
rect 160926 146911 160982 146920
rect 160940 113830 160968 146911
rect 160928 113824 160980 113830
rect 160928 113766 160980 113772
rect 161492 80034 161520 233174
rect 161480 80028 161532 80034
rect 161480 79970 161532 79976
rect 160836 73840 160888 73846
rect 160836 73782 160888 73788
rect 160744 70304 160796 70310
rect 160744 70246 160796 70252
rect 157984 31068 158036 31074
rect 157984 31010 158036 31016
rect 162136 17270 162164 253807
rect 162228 193866 162256 299406
rect 162676 245676 162728 245682
rect 162676 245618 162728 245624
rect 162688 244361 162716 245618
rect 162674 244352 162730 244361
rect 162674 244287 162730 244296
rect 162780 242010 162808 373866
rect 163884 365634 163912 384231
rect 163872 365628 163924 365634
rect 163872 365570 163924 365576
rect 163596 294636 163648 294642
rect 163596 294578 163648 294584
rect 163504 285728 163556 285734
rect 163504 285670 163556 285676
rect 163516 268394 163544 285670
rect 163608 280090 163636 294578
rect 163688 290488 163740 290494
rect 163976 290465 164004 441594
rect 164068 292534 164096 474710
rect 164146 457464 164202 457473
rect 164146 457399 164202 457408
rect 164056 292528 164108 292534
rect 164056 292470 164108 292476
rect 163688 290430 163740 290436
rect 163962 290456 164018 290465
rect 163700 280838 163728 290430
rect 163962 290391 164018 290400
rect 163688 280832 163740 280838
rect 163688 280774 163740 280780
rect 163596 280084 163648 280090
rect 163596 280026 163648 280032
rect 164056 280084 164108 280090
rect 164056 280026 164108 280032
rect 164068 279478 164096 280026
rect 164056 279472 164108 279478
rect 164056 279414 164108 279420
rect 163504 268388 163556 268394
rect 163504 268330 163556 268336
rect 162858 266384 162914 266393
rect 162858 266319 162914 266328
rect 162308 242004 162360 242010
rect 162308 241946 162360 241952
rect 162768 242004 162820 242010
rect 162768 241946 162820 241952
rect 162320 241534 162348 241946
rect 162308 241528 162360 241534
rect 162308 241470 162360 241476
rect 162320 233238 162348 241470
rect 162308 233232 162360 233238
rect 162308 233174 162360 233180
rect 162216 193860 162268 193866
rect 162216 193802 162268 193808
rect 162872 19990 162900 266319
rect 163504 252612 163556 252618
rect 163504 252554 163556 252560
rect 163516 218657 163544 252554
rect 163502 218648 163558 218657
rect 163502 218583 163558 218592
rect 163516 107642 163544 218583
rect 164068 166326 164096 279414
rect 164160 262206 164188 457399
rect 164896 384985 164924 592078
rect 165068 542496 165120 542502
rect 165068 542438 165120 542444
rect 164976 527944 165028 527950
rect 164976 527886 165028 527892
rect 164988 460934 165016 527886
rect 165080 465730 165108 542438
rect 165620 524408 165672 524414
rect 165620 524350 165672 524356
rect 165528 491972 165580 491978
rect 165528 491914 165580 491920
rect 165068 465724 165120 465730
rect 165068 465666 165120 465672
rect 164988 460906 165108 460934
rect 165080 446486 165108 460906
rect 165068 446480 165120 446486
rect 165068 446422 165120 446428
rect 164976 430568 165028 430574
rect 164976 430510 165028 430516
rect 164882 384976 164938 384985
rect 164882 384911 164938 384920
rect 164884 328568 164936 328574
rect 164884 328510 164936 328516
rect 164148 262200 164200 262206
rect 164148 262142 164200 262148
rect 164056 166320 164108 166326
rect 164056 166262 164108 166268
rect 163504 107636 163556 107642
rect 163504 107578 163556 107584
rect 164896 98122 164924 328510
rect 164988 289202 165016 430510
rect 165080 422294 165108 446422
rect 165436 431248 165488 431254
rect 165436 431190 165488 431196
rect 165448 430574 165476 431190
rect 165436 430568 165488 430574
rect 165436 430510 165488 430516
rect 165080 422266 165476 422294
rect 165448 411942 165476 422266
rect 165436 411936 165488 411942
rect 165436 411878 165488 411884
rect 165448 316742 165476 411878
rect 165540 336161 165568 491914
rect 165632 464234 165660 524350
rect 165620 464228 165672 464234
rect 165620 464170 165672 464176
rect 165632 463758 165660 464170
rect 165620 463752 165672 463758
rect 165620 463694 165672 463700
rect 165620 425128 165672 425134
rect 165620 425070 165672 425076
rect 165526 336152 165582 336161
rect 165526 336087 165582 336096
rect 165540 336054 165568 336087
rect 165528 336048 165580 336054
rect 165528 335990 165580 335996
rect 165436 316736 165488 316742
rect 165436 316678 165488 316684
rect 164976 289196 165028 289202
rect 164976 289138 165028 289144
rect 165632 284889 165660 425070
rect 166276 387938 166304 594866
rect 168288 585200 168340 585206
rect 168288 585142 168340 585148
rect 166356 574116 166408 574122
rect 166356 574058 166408 574064
rect 166368 414633 166396 574058
rect 166448 556232 166500 556238
rect 166448 556174 166500 556180
rect 166460 524414 166488 556174
rect 167644 552084 167696 552090
rect 167644 552026 167696 552032
rect 166540 541000 166592 541006
rect 166540 540942 166592 540948
rect 166552 529242 166580 540942
rect 166540 529236 166592 529242
rect 166540 529178 166592 529184
rect 166448 524408 166500 524414
rect 166448 524350 166500 524356
rect 166540 487892 166592 487898
rect 166540 487834 166592 487840
rect 166448 464228 166500 464234
rect 166448 464170 166500 464176
rect 166460 460193 166488 464170
rect 166446 460184 166502 460193
rect 166446 460119 166502 460128
rect 166446 453248 166502 453257
rect 166446 453183 166502 453192
rect 166460 452674 166488 453183
rect 166448 452668 166500 452674
rect 166448 452610 166500 452616
rect 166354 414624 166410 414633
rect 166354 414559 166410 414568
rect 166356 393372 166408 393378
rect 166356 393314 166408 393320
rect 166264 387932 166316 387938
rect 166264 387874 166316 387880
rect 166368 368422 166396 393314
rect 165712 368416 165764 368422
rect 165712 368358 165764 368364
rect 166356 368416 166408 368422
rect 166356 368358 166408 368364
rect 165618 284880 165674 284889
rect 165618 284815 165674 284824
rect 165632 284345 165660 284815
rect 165618 284336 165674 284345
rect 165618 284271 165674 284280
rect 165068 269816 165120 269822
rect 165068 269758 165120 269764
rect 164976 264988 165028 264994
rect 164976 264930 165028 264936
rect 164148 98116 164200 98122
rect 164148 98058 164200 98064
rect 164884 98116 164936 98122
rect 164884 98058 164936 98064
rect 164160 81258 164188 98058
rect 164148 81252 164200 81258
rect 164148 81194 164200 81200
rect 164988 71058 165016 264930
rect 165080 238649 165108 269758
rect 165724 240106 165752 368358
rect 166262 330576 166318 330585
rect 166262 330511 166318 330520
rect 166276 329866 166304 330511
rect 166264 329860 166316 329866
rect 166264 329802 166316 329808
rect 166262 302832 166318 302841
rect 166262 302767 166318 302776
rect 166276 251938 166304 302767
rect 166460 296002 166488 452610
rect 166552 428505 166580 487834
rect 167656 483721 167684 552026
rect 168194 529136 168250 529145
rect 168194 529071 168250 529080
rect 168104 504416 168156 504422
rect 168104 504358 168156 504364
rect 167642 483712 167698 483721
rect 167642 483647 167698 483656
rect 167644 463752 167696 463758
rect 167644 463694 167696 463700
rect 166538 428496 166594 428505
rect 166538 428431 166594 428440
rect 166998 369880 167054 369889
rect 166998 369815 167054 369824
rect 166448 295996 166500 296002
rect 166448 295938 166500 295944
rect 166356 284368 166408 284374
rect 166356 284310 166408 284316
rect 166446 284336 166502 284345
rect 166264 251932 166316 251938
rect 166264 251874 166316 251880
rect 165712 240100 165764 240106
rect 165712 240042 165764 240048
rect 165066 238640 165122 238649
rect 165066 238575 165122 238584
rect 165080 160138 165108 238575
rect 165068 160132 165120 160138
rect 165068 160074 165120 160080
rect 165080 133890 165108 160074
rect 165068 133884 165120 133890
rect 165068 133826 165120 133832
rect 164976 71052 165028 71058
rect 164976 70994 165028 71000
rect 166276 36582 166304 251874
rect 166368 251870 166396 284310
rect 166446 284271 166502 284280
rect 166460 267034 166488 284271
rect 166448 267028 166500 267034
rect 166448 266970 166500 266976
rect 166908 256080 166960 256086
rect 166908 256022 166960 256028
rect 166356 251864 166408 251870
rect 166356 251806 166408 251812
rect 166356 249076 166408 249082
rect 166356 249018 166408 249024
rect 166368 76566 166396 249018
rect 166920 231849 166948 256022
rect 166906 231840 166962 231849
rect 166906 231775 166962 231784
rect 166920 219434 166948 231775
rect 166460 219406 166948 219434
rect 166460 137057 166488 219406
rect 167012 211138 167040 369815
rect 167656 318073 167684 463694
rect 168116 397594 168144 504358
rect 168104 397588 168156 397594
rect 168104 397530 168156 397536
rect 168208 392018 168236 529071
rect 168196 392012 168248 392018
rect 168196 391954 168248 391960
rect 167736 387932 167788 387938
rect 167736 387874 167788 387880
rect 167748 386345 167776 387874
rect 168208 387190 168236 391954
rect 168196 387184 168248 387190
rect 168196 387126 168248 387132
rect 167734 386336 167790 386345
rect 167734 386271 167790 386280
rect 167748 371249 167776 386271
rect 167734 371240 167790 371249
rect 167734 371175 167790 371184
rect 167748 369889 167776 371175
rect 167734 369880 167790 369889
rect 167734 369815 167790 369824
rect 168194 369744 168250 369753
rect 168194 369679 168250 369688
rect 167642 318064 167698 318073
rect 167642 317999 167698 318008
rect 167090 285696 167146 285705
rect 167090 285631 167146 285640
rect 167104 261526 167132 285631
rect 167656 284306 167684 317999
rect 167644 284300 167696 284306
rect 167644 284242 167696 284248
rect 168208 266354 168236 369679
rect 168300 368422 168328 585142
rect 169036 449206 169064 604454
rect 170404 594924 170456 594930
rect 170404 594866 170456 594872
rect 169114 579728 169170 579737
rect 169114 579663 169170 579672
rect 169760 579692 169812 579698
rect 169128 489161 169156 579663
rect 169760 579634 169812 579640
rect 169208 565140 169260 565146
rect 169208 565082 169260 565088
rect 169220 513369 169248 565082
rect 169576 561740 169628 561746
rect 169576 561682 169628 561688
rect 169206 513360 169262 513369
rect 169206 513295 169208 513304
rect 169260 513295 169262 513304
rect 169208 513266 169260 513272
rect 169220 513235 169248 513266
rect 169484 505776 169536 505782
rect 169484 505718 169536 505724
rect 169114 489152 169170 489161
rect 169114 489087 169170 489096
rect 169024 449200 169076 449206
rect 169024 449142 169076 449148
rect 169036 427106 169064 449142
rect 169024 427100 169076 427106
rect 169024 427042 169076 427048
rect 169392 424516 169444 424522
rect 169392 424458 169444 424464
rect 169024 401600 169076 401606
rect 169024 401542 169076 401548
rect 168380 389836 168432 389842
rect 168380 389778 168432 389784
rect 168392 389298 168420 389778
rect 168380 389292 168432 389298
rect 168380 389234 168432 389240
rect 168288 368416 168340 368422
rect 168288 368358 168340 368364
rect 169036 365673 169064 401542
rect 169022 365664 169078 365673
rect 169022 365599 169078 365608
rect 168288 268388 168340 268394
rect 168288 268330 168340 268336
rect 168196 266348 168248 266354
rect 168196 266290 168248 266296
rect 168208 264994 168236 266290
rect 168196 264988 168248 264994
rect 168196 264930 168248 264936
rect 167092 261520 167144 261526
rect 167092 261462 167144 261468
rect 167642 260536 167698 260545
rect 167642 260471 167698 260480
rect 167000 211132 167052 211138
rect 167000 211074 167052 211080
rect 166446 137048 166502 137057
rect 166446 136983 166502 136992
rect 166460 109002 166488 136983
rect 166448 108996 166500 109002
rect 166448 108938 166500 108944
rect 166356 76560 166408 76566
rect 166356 76502 166408 76508
rect 166368 74458 166396 76502
rect 167656 75206 167684 260471
rect 168300 235929 168328 268330
rect 168380 262200 168432 262206
rect 168380 262142 168432 262148
rect 168392 260914 168420 262142
rect 168380 260908 168432 260914
rect 168380 260850 168432 260856
rect 168286 235920 168342 235929
rect 168286 235855 168342 235864
rect 168300 234705 168328 235855
rect 167734 234696 167790 234705
rect 167734 234631 167790 234640
rect 168286 234696 168342 234705
rect 168286 234631 168342 234640
rect 167748 179450 167776 234631
rect 167736 179444 167788 179450
rect 167736 179386 167788 179392
rect 167748 125594 167776 179386
rect 167736 125588 167788 125594
rect 167736 125530 167788 125536
rect 167644 75200 167696 75206
rect 167644 75142 167696 75148
rect 166356 74452 166408 74458
rect 166356 74394 166408 74400
rect 166264 36576 166316 36582
rect 166264 36518 166316 36524
rect 162860 19984 162912 19990
rect 162860 19926 162912 19932
rect 162124 17264 162176 17270
rect 162124 17206 162176 17212
rect 155224 13116 155276 13122
rect 155224 13058 155276 13064
rect 168392 8974 168420 260850
rect 169036 257378 169064 365599
rect 169404 326398 169432 424458
rect 169496 389298 169524 505718
rect 169588 424386 169616 561682
rect 169772 542366 169800 579634
rect 169760 542360 169812 542366
rect 169760 542302 169812 542308
rect 169772 541686 169800 542302
rect 169760 541680 169812 541686
rect 169760 541622 169812 541628
rect 170416 503033 170444 594866
rect 172334 589928 172390 589937
rect 172334 589863 172390 589872
rect 170956 560312 171008 560318
rect 170956 560254 171008 560260
rect 170496 539640 170548 539646
rect 170496 539582 170548 539588
rect 170402 503024 170458 503033
rect 170402 502959 170458 502968
rect 170508 471209 170536 539582
rect 170772 501628 170824 501634
rect 170772 501570 170824 501576
rect 170494 471200 170550 471209
rect 170494 471135 170550 471144
rect 169666 465760 169722 465769
rect 169666 465695 169722 465704
rect 169576 424380 169628 424386
rect 169576 424322 169628 424328
rect 169484 389292 169536 389298
rect 169484 389234 169536 389240
rect 169392 326392 169444 326398
rect 169392 326334 169444 326340
rect 169114 311400 169170 311409
rect 169114 311335 169170 311344
rect 169128 269890 169156 311335
rect 169208 300144 169260 300150
rect 169208 300086 169260 300092
rect 169116 269884 169168 269890
rect 169116 269826 169168 269832
rect 169116 267096 169168 267102
rect 169116 267038 169168 267044
rect 169024 257372 169076 257378
rect 169024 257314 169076 257320
rect 169024 240100 169076 240106
rect 169024 240042 169076 240048
rect 169036 239426 169064 240042
rect 169024 239420 169076 239426
rect 169024 239362 169076 239368
rect 169036 84182 169064 239362
rect 169128 235793 169156 267038
rect 169220 264314 169248 300086
rect 169680 287774 169708 465695
rect 170784 439521 170812 501570
rect 170862 471200 170918 471209
rect 170862 471135 170918 471144
rect 170770 439512 170826 439521
rect 170770 439447 170826 439456
rect 170404 435396 170456 435402
rect 170404 435338 170456 435344
rect 170416 423638 170444 435338
rect 170404 423632 170456 423638
rect 170404 423574 170456 423580
rect 169760 397588 169812 397594
rect 169760 397530 169812 397536
rect 169772 372570 169800 397530
rect 170876 396030 170904 471135
rect 170968 465769 170996 560254
rect 171784 553444 171836 553450
rect 171784 553386 171836 553392
rect 171048 518288 171100 518294
rect 171048 518230 171100 518236
rect 170954 465760 171010 465769
rect 170954 465695 171010 465704
rect 170864 396024 170916 396030
rect 170864 395966 170916 395972
rect 170954 390824 171010 390833
rect 170954 390759 171010 390768
rect 170494 386200 170550 386209
rect 170494 386135 170550 386144
rect 170508 385694 170536 386135
rect 170496 385688 170548 385694
rect 170496 385630 170548 385636
rect 169760 372564 169812 372570
rect 169760 372506 169812 372512
rect 169772 371278 169800 372506
rect 169760 371272 169812 371278
rect 169760 371214 169812 371220
rect 170404 371272 170456 371278
rect 170404 371214 170456 371220
rect 170416 325694 170444 371214
rect 170508 366897 170536 385630
rect 170494 366888 170550 366897
rect 170494 366823 170550 366832
rect 170416 325666 170628 325694
rect 170600 314770 170628 325666
rect 170588 314764 170640 314770
rect 170588 314706 170640 314712
rect 170404 300824 170456 300830
rect 170404 300766 170456 300772
rect 169668 287768 169720 287774
rect 169668 287710 169720 287716
rect 169208 264308 169260 264314
rect 169208 264250 169260 264256
rect 169298 260536 169354 260545
rect 169298 260471 169354 260480
rect 169312 260234 169340 260471
rect 169300 260228 169352 260234
rect 169300 260170 169352 260176
rect 170416 256018 170444 300766
rect 170496 289944 170548 289950
rect 170496 289886 170548 289892
rect 170508 260166 170536 289886
rect 170600 285734 170628 314706
rect 170968 306374 170996 390759
rect 171060 383625 171088 518230
rect 171796 492046 171824 553386
rect 172244 497480 172296 497486
rect 172244 497422 172296 497428
rect 171784 492040 171836 492046
rect 171784 491982 171836 491988
rect 171782 462904 171838 462913
rect 171782 462839 171838 462848
rect 171046 383616 171102 383625
rect 171046 383551 171102 383560
rect 171796 369753 171824 462839
rect 171968 393984 172020 393990
rect 171968 393926 172020 393932
rect 171874 386200 171930 386209
rect 171874 386135 171930 386144
rect 171782 369744 171838 369753
rect 171782 369679 171838 369688
rect 171888 365702 171916 386135
rect 171980 375290 172008 393926
rect 172256 386209 172284 497422
rect 172348 457609 172376 589863
rect 173162 581088 173218 581097
rect 173162 581023 173218 581032
rect 172428 574796 172480 574802
rect 172428 574738 172480 574744
rect 172334 457600 172390 457609
rect 172334 457535 172390 457544
rect 172336 450016 172388 450022
rect 172336 449958 172388 449964
rect 172348 449750 172376 449958
rect 172336 449744 172388 449750
rect 172336 449686 172388 449692
rect 172440 393961 172468 574738
rect 173176 554033 173204 581023
rect 173162 554024 173218 554033
rect 173162 553959 173218 553968
rect 173624 548548 173676 548554
rect 173624 548490 173676 548496
rect 173532 502988 173584 502994
rect 173532 502930 173584 502936
rect 173544 401606 173572 502930
rect 173636 441590 173664 548490
rect 173716 445800 173768 445806
rect 173716 445742 173768 445748
rect 173624 441584 173676 441590
rect 173624 441526 173676 441532
rect 173636 440881 173664 441526
rect 173622 440872 173678 440881
rect 173622 440807 173678 440816
rect 173532 401600 173584 401606
rect 173532 401542 173584 401548
rect 173162 398032 173218 398041
rect 173162 397967 173218 397976
rect 172426 393952 172482 393961
rect 172426 393887 172482 393896
rect 172242 386200 172298 386209
rect 172242 386135 172298 386144
rect 173176 379273 173204 397967
rect 173624 387864 173676 387870
rect 173624 387806 173676 387812
rect 173636 387705 173664 387806
rect 173622 387696 173678 387705
rect 173622 387631 173678 387640
rect 173622 381712 173678 381721
rect 173622 381647 173678 381656
rect 173636 381546 173664 381647
rect 173624 381540 173676 381546
rect 173624 381482 173676 381488
rect 173162 379264 173218 379273
rect 173162 379199 173218 379208
rect 171968 375284 172020 375290
rect 171968 375226 172020 375232
rect 171232 365696 171284 365702
rect 171232 365638 171284 365644
rect 171876 365696 171928 365702
rect 171876 365638 171928 365644
rect 170968 306346 171088 306374
rect 170588 285728 170640 285734
rect 170588 285670 170640 285676
rect 171060 285666 171088 306346
rect 171140 296744 171192 296750
rect 171140 296686 171192 296692
rect 171152 293350 171180 296686
rect 171140 293344 171192 293350
rect 171140 293286 171192 293292
rect 171048 285660 171100 285666
rect 171048 285602 171100 285608
rect 170496 260160 170548 260166
rect 170496 260102 170548 260108
rect 170404 256012 170456 256018
rect 170404 255954 170456 255960
rect 170402 250472 170458 250481
rect 170402 250407 170458 250416
rect 169760 237380 169812 237386
rect 169760 237322 169812 237328
rect 169772 237289 169800 237322
rect 169758 237280 169814 237289
rect 169758 237215 169814 237224
rect 169114 235784 169170 235793
rect 169114 235719 169170 235728
rect 169666 235784 169722 235793
rect 169666 235719 169722 235728
rect 169680 143614 169708 235719
rect 169760 214600 169812 214606
rect 169760 214542 169812 214548
rect 169772 213926 169800 214542
rect 169760 213920 169812 213926
rect 169760 213862 169812 213868
rect 169772 163538 169800 213862
rect 169760 163532 169812 163538
rect 169760 163474 169812 163480
rect 169668 143608 169720 143614
rect 169668 143550 169720 143556
rect 169680 136649 169708 143550
rect 169666 136640 169722 136649
rect 169666 136575 169722 136584
rect 169116 106956 169168 106962
rect 169116 106898 169168 106904
rect 169024 84176 169076 84182
rect 169024 84118 169076 84124
rect 169128 75886 169156 106898
rect 169116 75880 169168 75886
rect 169116 75822 169168 75828
rect 170416 35222 170444 250407
rect 170496 150544 170548 150550
rect 170496 150486 170548 150492
rect 170508 130422 170536 150486
rect 170496 130416 170548 130422
rect 170496 130358 170548 130364
rect 170496 114572 170548 114578
rect 170496 114514 170548 114520
rect 170508 68950 170536 114514
rect 171060 93158 171088 285602
rect 171140 258188 171192 258194
rect 171140 258130 171192 258136
rect 171152 257961 171180 258130
rect 171138 257952 171194 257961
rect 171138 257887 171194 257896
rect 171048 93152 171100 93158
rect 171048 93094 171100 93100
rect 170496 68944 170548 68950
rect 170496 68886 170548 68892
rect 170404 35216 170456 35222
rect 170404 35158 170456 35164
rect 171152 28286 171180 257887
rect 171244 239873 171272 365638
rect 172336 351212 172388 351218
rect 172336 351154 172388 351160
rect 171782 341456 171838 341465
rect 171782 341391 171838 341400
rect 171796 302258 171824 341391
rect 172242 330440 172298 330449
rect 172242 330375 172298 330384
rect 172256 329934 172284 330375
rect 172244 329928 172296 329934
rect 172244 329870 172296 329876
rect 171784 302252 171836 302258
rect 171784 302194 171836 302200
rect 172244 302252 172296 302258
rect 172244 302194 172296 302200
rect 172256 300830 172284 302194
rect 172244 300824 172296 300830
rect 172244 300766 172296 300772
rect 171784 293276 171836 293282
rect 171784 293218 171836 293224
rect 171796 273970 171824 293218
rect 171784 273964 171836 273970
rect 171784 273906 171836 273912
rect 172348 273222 172376 351154
rect 172428 333260 172480 333266
rect 172428 333202 172480 333208
rect 172336 273216 172388 273222
rect 172336 273158 172388 273164
rect 172348 272610 172376 273158
rect 172336 272604 172388 272610
rect 172336 272546 172388 272552
rect 171784 247784 171836 247790
rect 171784 247726 171836 247732
rect 171230 239864 171286 239873
rect 171230 239799 171286 239808
rect 171796 224913 171824 247726
rect 171782 224904 171838 224913
rect 171782 224839 171838 224848
rect 172336 216708 172388 216714
rect 172336 216650 172388 216656
rect 172348 211041 172376 216650
rect 172334 211032 172390 211041
rect 172334 210967 172390 210976
rect 172348 92857 172376 210967
rect 172440 179450 172468 333202
rect 172520 308440 172572 308446
rect 172520 308382 172572 308388
rect 172532 307834 172560 308382
rect 172520 307828 172572 307834
rect 172520 307770 172572 307776
rect 172532 262954 172560 307770
rect 173636 286346 173664 381482
rect 173728 331906 173756 445742
rect 173716 331900 173768 331906
rect 173716 331842 173768 331848
rect 173714 322960 173770 322969
rect 173714 322895 173770 322904
rect 173624 286340 173676 286346
rect 173624 286282 173676 286288
rect 173254 270464 173310 270473
rect 173254 270399 173310 270408
rect 172520 262948 172572 262954
rect 172520 262890 172572 262896
rect 173162 244352 173218 244361
rect 173162 244287 173218 244296
rect 172518 239864 172574 239873
rect 172518 239799 172574 239808
rect 172532 239465 172560 239799
rect 172518 239456 172574 239465
rect 172518 239391 172574 239400
rect 172428 179444 172480 179450
rect 172428 179386 172480 179392
rect 172440 176633 172468 179386
rect 172426 176624 172482 176633
rect 172426 176559 172482 176568
rect 172334 92848 172390 92857
rect 172334 92783 172390 92792
rect 172532 81326 172560 239391
rect 172520 81320 172572 81326
rect 172520 81262 172572 81268
rect 173176 33794 173204 244287
rect 173268 238134 173296 270399
rect 173728 244633 173756 322895
rect 173820 311273 173848 611351
rect 177396 607232 177448 607238
rect 177396 607174 177448 607180
rect 177304 603152 177356 603158
rect 177304 603094 177356 603100
rect 175188 594176 175240 594182
rect 175188 594118 175240 594124
rect 175096 592680 175148 592686
rect 175096 592622 175148 592628
rect 175108 592074 175136 592622
rect 175096 592068 175148 592074
rect 175096 592010 175148 592016
rect 175108 586514 175136 592010
rect 175016 586486 175136 586514
rect 175016 469266 175044 586486
rect 175094 482216 175150 482225
rect 175094 482151 175150 482160
rect 174544 469260 174596 469266
rect 174544 469202 174596 469208
rect 175004 469260 175056 469266
rect 175004 469202 175056 469208
rect 174556 441522 174584 469202
rect 175002 450256 175058 450265
rect 175002 450191 175058 450200
rect 175016 449954 175044 450191
rect 175004 449948 175056 449954
rect 175004 449890 175056 449896
rect 174544 441516 174596 441522
rect 174544 441458 174596 441464
rect 174636 419552 174688 419558
rect 174636 419494 174688 419500
rect 173806 311264 173862 311273
rect 173806 311199 173862 311208
rect 174544 295996 174596 296002
rect 174544 295938 174596 295944
rect 173898 288416 173954 288425
rect 173898 288351 173954 288360
rect 173912 287745 173940 288351
rect 173898 287736 173954 287745
rect 173898 287671 173954 287680
rect 173808 280832 173860 280838
rect 173808 280774 173860 280780
rect 173714 244624 173770 244633
rect 173714 244559 173770 244568
rect 173728 244361 173756 244559
rect 173714 244352 173770 244361
rect 173714 244287 173770 244296
rect 173256 238128 173308 238134
rect 173256 238070 173308 238076
rect 173820 136610 173848 280774
rect 173912 256086 173940 287671
rect 173900 256080 173952 256086
rect 173900 256022 173952 256028
rect 174556 138689 174584 295938
rect 174648 288425 174676 419494
rect 175016 316034 175044 449890
rect 175108 342378 175136 482151
rect 175200 383042 175228 594118
rect 176568 581052 176620 581058
rect 176568 580994 176620 581000
rect 176476 545148 176528 545154
rect 176476 545090 176528 545096
rect 176384 479528 176436 479534
rect 176384 479470 176436 479476
rect 176108 447092 176160 447098
rect 176108 447034 176160 447040
rect 176120 446418 176148 447034
rect 176108 446412 176160 446418
rect 176108 446354 176160 446360
rect 176396 389162 176424 479470
rect 176488 447098 176516 545090
rect 176476 447092 176528 447098
rect 176476 447034 176528 447040
rect 176476 437504 176528 437510
rect 176476 437446 176528 437452
rect 176384 389156 176436 389162
rect 176384 389098 176436 389104
rect 175188 383036 175240 383042
rect 175188 382978 175240 382984
rect 175556 345160 175608 345166
rect 175556 345102 175608 345108
rect 175568 343641 175596 345102
rect 175554 343632 175610 343641
rect 175554 343567 175610 343576
rect 175096 342372 175148 342378
rect 175096 342314 175148 342320
rect 175108 338774 175136 342314
rect 175096 338768 175148 338774
rect 175096 338710 175148 338716
rect 176488 324358 176516 437446
rect 176580 414730 176608 580994
rect 177316 445806 177344 603094
rect 177408 588606 177436 607174
rect 177396 588600 177448 588606
rect 177396 588542 177448 588548
rect 177396 582412 177448 582418
rect 177396 582354 177448 582360
rect 177408 538286 177436 582354
rect 177500 581670 177528 616898
rect 177488 581664 177540 581670
rect 177488 581606 177540 581612
rect 178788 547097 178816 618326
rect 178868 569220 178920 569226
rect 178868 569162 178920 569168
rect 178774 547088 178830 547097
rect 178774 547023 178830 547032
rect 178684 546576 178736 546582
rect 178684 546518 178736 546524
rect 177396 538280 177448 538286
rect 177396 538222 177448 538228
rect 177396 512644 177448 512650
rect 177396 512586 177448 512592
rect 177304 445800 177356 445806
rect 177304 445742 177356 445748
rect 177408 421598 177436 512586
rect 177488 482316 177540 482322
rect 177488 482258 177540 482264
rect 177396 421592 177448 421598
rect 177396 421534 177448 421540
rect 177304 416832 177356 416838
rect 177304 416774 177356 416780
rect 176568 414724 176620 414730
rect 176568 414666 176620 414672
rect 177316 409834 177344 416774
rect 177304 409828 177356 409834
rect 177304 409770 177356 409776
rect 177396 406428 177448 406434
rect 177396 406370 177448 406376
rect 176660 402348 176712 402354
rect 176660 402290 176712 402296
rect 176672 401674 176700 402290
rect 176660 401668 176712 401674
rect 176660 401610 176712 401616
rect 177302 390960 177358 390969
rect 177302 390895 177358 390904
rect 175924 324352 175976 324358
rect 175924 324294 175976 324300
rect 176476 324352 176528 324358
rect 176476 324294 176528 324300
rect 175186 316160 175242 316169
rect 175186 316095 175242 316104
rect 175200 316034 175228 316095
rect 175016 316006 175228 316034
rect 174728 309800 174780 309806
rect 174728 309742 174780 309748
rect 174634 288416 174690 288425
rect 174634 288351 174690 288360
rect 174740 272542 174768 309742
rect 175200 302938 175228 316006
rect 175188 302932 175240 302938
rect 175188 302874 175240 302880
rect 175200 302569 175228 302874
rect 175186 302560 175242 302569
rect 175186 302495 175242 302504
rect 175648 300892 175700 300898
rect 175648 300834 175700 300840
rect 175660 297430 175688 300834
rect 175648 297424 175700 297430
rect 175648 297366 175700 297372
rect 175936 296070 175964 324294
rect 177316 322969 177344 390895
rect 177408 385694 177436 406370
rect 177500 393378 177528 482258
rect 177580 447908 177632 447914
rect 177580 447850 177632 447856
rect 177592 437510 177620 447850
rect 177580 437504 177632 437510
rect 177580 437446 177632 437452
rect 178040 427100 178092 427106
rect 178040 427042 178092 427048
rect 178052 426494 178080 427042
rect 178040 426488 178092 426494
rect 178040 426430 178092 426436
rect 177948 401668 178000 401674
rect 177948 401610 178000 401616
rect 177856 400648 177908 400654
rect 177856 400590 177908 400596
rect 177868 400246 177896 400590
rect 177856 400240 177908 400246
rect 177856 400182 177908 400188
rect 177488 393372 177540 393378
rect 177488 393314 177540 393320
rect 177500 391338 177528 393314
rect 177488 391332 177540 391338
rect 177488 391274 177540 391280
rect 177396 385688 177448 385694
rect 177396 385630 177448 385636
rect 177670 382392 177726 382401
rect 177670 382327 177726 382336
rect 177396 334620 177448 334626
rect 177396 334562 177448 334568
rect 177302 322960 177358 322969
rect 177302 322895 177358 322904
rect 176016 317484 176068 317490
rect 176016 317426 176068 317432
rect 175924 296064 175976 296070
rect 175924 296006 175976 296012
rect 175924 282940 175976 282946
rect 175924 282882 175976 282888
rect 174728 272536 174780 272542
rect 174728 272478 174780 272484
rect 174636 267028 174688 267034
rect 174636 266970 174688 266976
rect 174648 233238 174676 266970
rect 175186 256048 175242 256057
rect 175186 255983 175188 255992
rect 175240 255983 175242 255992
rect 175188 255954 175240 255960
rect 174728 250504 174780 250510
rect 174728 250446 174780 250452
rect 174740 241466 174768 250446
rect 174728 241460 174780 241466
rect 174728 241402 174780 241408
rect 174636 233232 174688 233238
rect 174636 233174 174688 233180
rect 175188 233232 175240 233238
rect 175188 233174 175240 233180
rect 174542 138680 174598 138689
rect 174542 138615 174598 138624
rect 174556 138145 174584 138615
rect 174542 138136 174598 138145
rect 174542 138071 174598 138080
rect 173808 136604 173860 136610
rect 173808 136546 173860 136552
rect 173256 117972 173308 117978
rect 173256 117914 173308 117920
rect 173268 77178 173296 117914
rect 175200 115938 175228 233174
rect 175936 229158 175964 282882
rect 176028 280838 176056 317426
rect 176658 312080 176714 312089
rect 176658 312015 176714 312024
rect 176672 311409 176700 312015
rect 176658 311400 176714 311409
rect 176658 311335 176714 311344
rect 176658 309768 176714 309777
rect 176658 309703 176714 309712
rect 176106 306776 176162 306785
rect 176106 306711 176162 306720
rect 176120 298081 176148 306711
rect 176106 298072 176162 298081
rect 176106 298007 176162 298016
rect 176200 294024 176252 294030
rect 176200 293966 176252 293972
rect 176108 292460 176160 292466
rect 176108 292402 176160 292408
rect 176016 280832 176068 280838
rect 176016 280774 176068 280780
rect 176016 253224 176068 253230
rect 176016 253166 176068 253172
rect 175924 229152 175976 229158
rect 175924 229094 175976 229100
rect 175936 188358 175964 229094
rect 176028 207874 176056 253166
rect 176120 249082 176148 292402
rect 176212 280158 176240 293966
rect 176200 280152 176252 280158
rect 176200 280094 176252 280100
rect 176212 249121 176240 280094
rect 176672 268394 176700 309703
rect 177408 289882 177436 334562
rect 177684 312089 177712 382327
rect 177868 382226 177896 400182
rect 177856 382220 177908 382226
rect 177856 382162 177908 382168
rect 177762 342952 177818 342961
rect 177762 342887 177818 342896
rect 177670 312080 177726 312089
rect 177670 312015 177726 312024
rect 177486 310584 177542 310593
rect 177486 310519 177542 310528
rect 177396 289876 177448 289882
rect 177396 289818 177448 289824
rect 177408 277394 177436 289818
rect 177316 277366 177436 277394
rect 176660 268388 176712 268394
rect 176660 268330 176712 268336
rect 176658 260128 176714 260137
rect 176658 260063 176714 260072
rect 176672 259486 176700 260063
rect 176660 259480 176712 259486
rect 176660 259422 176712 259428
rect 176198 249112 176254 249121
rect 176108 249076 176160 249082
rect 176198 249047 176254 249056
rect 176108 249018 176160 249024
rect 176568 208344 176620 208350
rect 176568 208286 176620 208292
rect 176580 207874 176608 208286
rect 176016 207868 176068 207874
rect 176016 207810 176068 207816
rect 176568 207868 176620 207874
rect 176568 207810 176620 207816
rect 175924 188352 175976 188358
rect 175924 188294 175976 188300
rect 175922 156224 175978 156233
rect 175922 156159 175978 156168
rect 175936 124914 175964 156159
rect 176580 146305 176608 207810
rect 176014 146296 176070 146305
rect 176014 146231 176070 146240
rect 176566 146296 176622 146305
rect 176566 146231 176622 146240
rect 176028 145081 176056 146231
rect 176014 145072 176070 145081
rect 176014 145007 176070 145016
rect 176028 141409 176056 145007
rect 176014 141400 176070 141409
rect 176014 141335 176070 141344
rect 176014 138136 176070 138145
rect 176014 138071 176070 138080
rect 176028 131102 176056 138071
rect 176016 131096 176068 131102
rect 176016 131038 176068 131044
rect 176028 130422 176056 131038
rect 176016 130416 176068 130422
rect 176016 130358 176068 130364
rect 176568 130416 176620 130422
rect 176568 130358 176620 130364
rect 175924 124908 175976 124914
rect 175924 124850 175976 124856
rect 175188 115932 175240 115938
rect 175188 115874 175240 115880
rect 173808 81320 173860 81326
rect 173808 81262 173860 81268
rect 173820 78606 173848 81262
rect 173808 78600 173860 78606
rect 173808 78542 173860 78548
rect 173256 77172 173308 77178
rect 173256 77114 173308 77120
rect 176580 65521 176608 130358
rect 176672 76537 176700 259422
rect 177316 144974 177344 277366
rect 177500 276690 177528 310519
rect 177488 276684 177540 276690
rect 177488 276626 177540 276632
rect 177396 275392 177448 275398
rect 177396 275334 177448 275340
rect 177408 237318 177436 275334
rect 177776 255270 177804 342887
rect 177960 341630 177988 401610
rect 178038 398848 178094 398857
rect 178038 398783 178094 398792
rect 178052 390969 178080 398783
rect 178696 397526 178724 546518
rect 178880 538218 178908 569162
rect 180076 542366 180104 702442
rect 182088 608728 182140 608734
rect 182088 608670 182140 608676
rect 180708 605872 180760 605878
rect 180708 605814 180760 605820
rect 180156 599072 180208 599078
rect 180156 599014 180208 599020
rect 180168 560998 180196 599014
rect 180156 560992 180208 560998
rect 180156 560934 180208 560940
rect 180156 554804 180208 554810
rect 180156 554746 180208 554752
rect 180168 545086 180196 554746
rect 180156 545080 180208 545086
rect 180156 545022 180208 545028
rect 179420 542360 179472 542366
rect 179420 542302 179472 542308
rect 180064 542360 180116 542366
rect 180064 542302 180116 542308
rect 178868 538212 178920 538218
rect 178868 538154 178920 538160
rect 179432 535514 179460 542302
rect 180614 539744 180670 539753
rect 180614 539679 180670 539688
rect 179510 538384 179566 538393
rect 179510 538319 179566 538328
rect 179340 535486 179460 535514
rect 178776 534744 178828 534750
rect 178776 534686 178828 534692
rect 178788 400654 178816 534686
rect 179340 532642 179368 535486
rect 179328 532636 179380 532642
rect 179328 532578 179380 532584
rect 178868 519580 178920 519586
rect 178868 519522 178920 519528
rect 178880 454714 178908 519522
rect 178960 483676 179012 483682
rect 178960 483618 179012 483624
rect 178868 454708 178920 454714
rect 178868 454650 178920 454656
rect 178972 432002 179000 483618
rect 178960 431996 179012 432002
rect 178960 431938 179012 431944
rect 178972 430574 179000 431938
rect 178960 430568 179012 430574
rect 178960 430510 179012 430516
rect 179328 426488 179380 426494
rect 179328 426430 179380 426436
rect 178868 404388 178920 404394
rect 178868 404330 178920 404336
rect 178776 400648 178828 400654
rect 178776 400590 178828 400596
rect 178684 397520 178736 397526
rect 178684 397462 178736 397468
rect 178696 393990 178724 397462
rect 178684 393984 178736 393990
rect 178684 393926 178736 393932
rect 178038 390960 178094 390969
rect 178038 390895 178094 390904
rect 178776 371884 178828 371890
rect 178776 371826 178828 371832
rect 177948 341624 178000 341630
rect 177948 341566 178000 341572
rect 178684 317552 178736 317558
rect 178684 317494 178736 317500
rect 178696 282946 178724 317494
rect 178684 282940 178736 282946
rect 178684 282882 178736 282888
rect 178682 269784 178738 269793
rect 178682 269719 178738 269728
rect 178696 257281 178724 269719
rect 178682 257272 178738 257281
rect 178682 257207 178738 257216
rect 177764 255264 177816 255270
rect 177764 255206 177816 255212
rect 177776 254017 177804 255206
rect 177762 254008 177818 254017
rect 177762 253943 177818 253952
rect 177396 237312 177448 237318
rect 177396 237254 177448 237260
rect 177396 233912 177448 233918
rect 177396 233854 177448 233860
rect 177408 211070 177436 233854
rect 177396 211064 177448 211070
rect 177396 211006 177448 211012
rect 177304 144968 177356 144974
rect 177304 144910 177356 144916
rect 177316 138718 177344 144910
rect 177304 138712 177356 138718
rect 177304 138654 177356 138660
rect 177304 104916 177356 104922
rect 177304 104858 177356 104864
rect 177316 80034 177344 104858
rect 177408 92177 177436 211006
rect 177394 92168 177450 92177
rect 177394 92103 177450 92112
rect 178040 82748 178092 82754
rect 178040 82690 178092 82696
rect 177304 80028 177356 80034
rect 177304 79970 177356 79976
rect 178052 78674 178080 82690
rect 178040 78668 178092 78674
rect 178040 78610 178092 78616
rect 176658 76528 176714 76537
rect 176658 76463 176714 76472
rect 176566 65512 176622 65521
rect 176566 65447 176622 65456
rect 173164 33788 173216 33794
rect 173164 33730 173216 33736
rect 171140 28280 171192 28286
rect 171140 28222 171192 28228
rect 178696 18630 178724 257207
rect 178788 240009 178816 371826
rect 178880 294030 178908 404330
rect 179144 390584 179196 390590
rect 179144 390526 179196 390532
rect 179156 387569 179184 390526
rect 179236 389836 179288 389842
rect 179236 389778 179288 389784
rect 179142 387560 179198 387569
rect 179142 387495 179198 387504
rect 179248 378078 179276 389778
rect 179236 378072 179288 378078
rect 179236 378014 179288 378020
rect 178868 294024 178920 294030
rect 178868 293966 178920 293972
rect 179248 280838 179276 378014
rect 179340 317558 179368 426430
rect 179420 417444 179472 417450
rect 179420 417386 179472 417392
rect 179432 416770 179460 417386
rect 179420 416764 179472 416770
rect 179420 416706 179472 416712
rect 179420 392624 179472 392630
rect 179420 392566 179472 392572
rect 179432 392057 179460 392566
rect 179418 392048 179474 392057
rect 179418 391983 179474 391992
rect 179524 390590 179552 538319
rect 180628 534070 180656 539679
rect 180616 534064 180668 534070
rect 180616 534006 180668 534012
rect 180628 485897 180656 534006
rect 180614 485888 180670 485897
rect 180614 485823 180670 485832
rect 180616 469872 180668 469878
rect 180616 469814 180668 469820
rect 180064 450628 180116 450634
rect 180064 450570 180116 450576
rect 180076 436762 180104 450570
rect 180064 436756 180116 436762
rect 180064 436698 180116 436704
rect 180522 435976 180578 435985
rect 180522 435911 180578 435920
rect 180536 417489 180564 435911
rect 180522 417480 180578 417489
rect 180522 417415 180578 417424
rect 180248 399492 180300 399498
rect 180248 399434 180300 399440
rect 179512 390584 179564 390590
rect 179512 390526 179564 390532
rect 180064 385688 180116 385694
rect 180064 385630 180116 385636
rect 179512 360120 179564 360126
rect 179512 360062 179564 360068
rect 179524 359718 179552 360062
rect 179512 359712 179564 359718
rect 179512 359654 179564 359660
rect 179328 317552 179380 317558
rect 179328 317494 179380 317500
rect 179236 280832 179288 280838
rect 179236 280774 179288 280780
rect 179248 277394 179276 280774
rect 179248 277366 179368 277394
rect 178868 242208 178920 242214
rect 178868 242150 178920 242156
rect 178774 240000 178830 240009
rect 178774 239935 178830 239944
rect 178880 224262 178908 242150
rect 179234 237960 179290 237969
rect 179234 237895 179290 237904
rect 179248 230450 179276 237895
rect 179236 230444 179288 230450
rect 179236 230386 179288 230392
rect 178868 224256 178920 224262
rect 178868 224198 178920 224204
rect 178776 103556 178828 103562
rect 178776 103498 178828 103504
rect 178788 81394 178816 103498
rect 179248 96665 179276 230386
rect 178866 96656 178922 96665
rect 178866 96591 178922 96600
rect 179234 96656 179290 96665
rect 179234 96591 179290 96600
rect 178880 92449 178908 96591
rect 178866 92440 178922 92449
rect 178866 92375 178922 92384
rect 179340 82754 179368 277366
rect 179420 262880 179472 262886
rect 179420 262822 179472 262828
rect 179432 262274 179460 262822
rect 179420 262268 179472 262274
rect 179420 262210 179472 262216
rect 179328 82748 179380 82754
rect 179328 82690 179380 82696
rect 178776 81388 178828 81394
rect 178776 81330 178828 81336
rect 179432 29646 179460 262210
rect 179524 247722 179552 359654
rect 180076 292466 180104 385630
rect 180154 384296 180210 384305
rect 180154 384231 180210 384240
rect 180168 359718 180196 384231
rect 180260 380769 180288 399434
rect 180628 388482 180656 469814
rect 180720 394097 180748 605814
rect 181904 575612 181956 575618
rect 181904 575554 181956 575560
rect 181916 480350 181944 575554
rect 181996 557592 182048 557598
rect 181996 557534 182048 557540
rect 181904 480344 181956 480350
rect 181904 480286 181956 480292
rect 181916 470594 181944 480286
rect 181548 470566 181944 470594
rect 181442 464536 181498 464545
rect 181442 464471 181498 464480
rect 180892 396772 180944 396778
rect 180892 396714 180944 396720
rect 180706 394088 180762 394097
rect 180706 394023 180762 394032
rect 180798 393408 180854 393417
rect 180798 393343 180854 393352
rect 180706 392048 180762 392057
rect 180706 391983 180762 391992
rect 180616 388476 180668 388482
rect 180616 388418 180668 388424
rect 180246 380760 180302 380769
rect 180246 380695 180302 380704
rect 180156 359712 180208 359718
rect 180156 359654 180208 359660
rect 180720 349926 180748 391983
rect 180812 367062 180840 393343
rect 180904 389842 180932 396714
rect 180892 389836 180944 389842
rect 180892 389778 180944 389784
rect 180800 367056 180852 367062
rect 180800 366998 180852 367004
rect 181456 351218 181484 464471
rect 181548 435402 181576 470566
rect 181536 435396 181588 435402
rect 181536 435338 181588 435344
rect 182008 405686 182036 557534
rect 182100 425066 182128 608670
rect 183468 604580 183520 604586
rect 183468 604522 183520 604528
rect 182824 582412 182876 582418
rect 182824 582354 182876 582360
rect 182836 570722 182864 582354
rect 183376 572008 183428 572014
rect 183376 571950 183428 571956
rect 182824 570716 182876 570722
rect 182824 570658 182876 570664
rect 183388 570654 183416 571950
rect 182916 570648 182968 570654
rect 182916 570590 182968 570596
rect 183376 570648 183428 570654
rect 183376 570590 183428 570596
rect 182824 554872 182876 554878
rect 182824 554814 182876 554820
rect 182180 451376 182232 451382
rect 182180 451318 182232 451324
rect 182192 448497 182220 451318
rect 182178 448488 182234 448497
rect 182178 448423 182234 448432
rect 182836 435985 182864 554814
rect 182928 484498 182956 570590
rect 183006 485072 183062 485081
rect 183006 485007 183062 485016
rect 182916 484492 182968 484498
rect 182916 484434 182968 484440
rect 182914 469296 182970 469305
rect 182914 469231 182970 469240
rect 182928 454889 182956 469231
rect 183020 467809 183048 485007
rect 183376 484492 183428 484498
rect 183376 484434 183428 484440
rect 183388 484362 183416 484434
rect 183376 484356 183428 484362
rect 183376 484298 183428 484304
rect 183006 467800 183062 467809
rect 183006 467735 183062 467744
rect 183284 465724 183336 465730
rect 183284 465666 183336 465672
rect 182914 454880 182970 454889
rect 182914 454815 182970 454824
rect 182822 435976 182878 435985
rect 182822 435911 182878 435920
rect 182088 425060 182140 425066
rect 182088 425002 182140 425008
rect 182100 424522 182128 425002
rect 182088 424516 182140 424522
rect 182088 424458 182140 424464
rect 182824 424380 182876 424386
rect 182824 424322 182876 424328
rect 182836 422294 182864 424322
rect 182836 422266 183232 422294
rect 183204 410582 183232 422266
rect 183192 410576 183244 410582
rect 183192 410518 183244 410524
rect 181628 405680 181680 405686
rect 181628 405622 181680 405628
rect 181996 405680 182048 405686
rect 181996 405622 182048 405628
rect 181640 404394 181668 405622
rect 181628 404388 181680 404394
rect 181628 404330 181680 404336
rect 182822 389328 182878 389337
rect 182822 389263 182878 389272
rect 182088 383036 182140 383042
rect 182088 382978 182140 382984
rect 181536 367056 181588 367062
rect 181536 366998 181588 367004
rect 181444 351212 181496 351218
rect 181444 351154 181496 351160
rect 180708 349920 180760 349926
rect 180708 349862 180760 349868
rect 180156 347064 180208 347070
rect 180156 347006 180208 347012
rect 180064 292460 180116 292466
rect 180064 292402 180116 292408
rect 180168 271862 180196 347006
rect 180246 289096 180302 289105
rect 180246 289031 180302 289040
rect 180156 271856 180208 271862
rect 180156 271798 180208 271804
rect 180168 258074 180196 271798
rect 180076 258046 180196 258074
rect 179512 247716 179564 247722
rect 179512 247658 179564 247664
rect 179524 247110 179552 247658
rect 179512 247104 179564 247110
rect 179512 247046 179564 247052
rect 180076 238746 180104 258046
rect 180260 256222 180288 289031
rect 180800 271176 180852 271182
rect 180800 271118 180852 271124
rect 180248 256216 180300 256222
rect 180248 256158 180300 256164
rect 180154 254008 180210 254017
rect 180154 253943 180210 253952
rect 180064 238740 180116 238746
rect 180064 238682 180116 238688
rect 180064 218748 180116 218754
rect 180064 218690 180116 218696
rect 180076 86873 180104 218690
rect 180168 202230 180196 253943
rect 180248 240780 180300 240786
rect 180248 240722 180300 240728
rect 180260 229809 180288 240722
rect 180812 238066 180840 271118
rect 181442 254144 181498 254153
rect 181442 254079 181498 254088
rect 180800 238060 180852 238066
rect 180800 238002 180852 238008
rect 180246 229800 180302 229809
rect 180246 229735 180302 229744
rect 180156 202224 180208 202230
rect 180156 202166 180208 202172
rect 180156 184204 180208 184210
rect 180156 184146 180208 184152
rect 180168 181490 180196 184146
rect 180156 181484 180208 181490
rect 180156 181426 180208 181432
rect 180168 117978 180196 181426
rect 180156 117972 180208 117978
rect 180156 117914 180208 117920
rect 180156 108316 180208 108322
rect 180156 108258 180208 108264
rect 180062 86864 180118 86873
rect 180062 86799 180118 86808
rect 180168 78674 180196 108258
rect 180156 78668 180208 78674
rect 180156 78610 180208 78616
rect 181456 77897 181484 254079
rect 181548 241097 181576 366998
rect 181994 320920 182050 320929
rect 181994 320855 182050 320864
rect 181720 271176 181772 271182
rect 181720 271118 181772 271124
rect 181732 270570 181760 271118
rect 181720 270564 181772 270570
rect 181720 270506 181772 270512
rect 182008 269074 182036 320855
rect 181996 269068 182048 269074
rect 181996 269010 182048 269016
rect 182008 268462 182036 269010
rect 181996 268456 182048 268462
rect 181996 268398 182048 268404
rect 182100 247489 182128 382978
rect 182836 371890 182864 389263
rect 182824 371884 182876 371890
rect 182824 371826 182876 371832
rect 183204 340202 183232 410518
rect 183296 390697 183324 465666
rect 183376 440292 183428 440298
rect 183376 440234 183428 440240
rect 183282 390688 183338 390697
rect 183282 390623 183338 390632
rect 183388 366382 183416 440234
rect 183480 439006 183508 604522
rect 184202 597816 184258 597825
rect 184202 597751 184258 597760
rect 184216 468625 184244 597751
rect 184308 578950 184336 702986
rect 202800 702982 202828 703520
rect 201500 702976 201552 702982
rect 201500 702918 201552 702924
rect 202788 702976 202840 702982
rect 202788 702918 202840 702924
rect 188896 702908 188948 702914
rect 188896 702850 188948 702856
rect 184848 615596 184900 615602
rect 184848 615538 184900 615544
rect 184388 605940 184440 605946
rect 184388 605882 184440 605888
rect 184400 596834 184428 605882
rect 184388 596828 184440 596834
rect 184388 596770 184440 596776
rect 184296 578944 184348 578950
rect 184296 578886 184348 578892
rect 184308 572694 184336 578886
rect 184296 572688 184348 572694
rect 184296 572630 184348 572636
rect 184664 554804 184716 554810
rect 184664 554746 184716 554752
rect 184676 486470 184704 554746
rect 184756 489184 184808 489190
rect 184756 489126 184808 489132
rect 184664 486464 184716 486470
rect 184664 486406 184716 486412
rect 184202 468616 184258 468625
rect 184202 468551 184258 468560
rect 184664 461032 184716 461038
rect 184664 460974 184716 460980
rect 184676 458833 184704 460974
rect 184662 458824 184718 458833
rect 184662 458759 184718 458768
rect 184204 456816 184256 456822
rect 184204 456758 184256 456764
rect 184216 445058 184244 456758
rect 184296 450560 184348 450566
rect 184296 450502 184348 450508
rect 184204 445052 184256 445058
rect 184204 444994 184256 445000
rect 184308 443766 184336 450502
rect 184296 443760 184348 443766
rect 184296 443702 184348 443708
rect 183468 439000 183520 439006
rect 183468 438942 183520 438948
rect 183468 437504 183520 437510
rect 183468 437446 183520 437452
rect 183376 366376 183428 366382
rect 183376 366318 183428 366324
rect 183374 351112 183430 351121
rect 183374 351047 183430 351056
rect 183192 340196 183244 340202
rect 183192 340138 183244 340144
rect 182822 306640 182878 306649
rect 182822 306575 182878 306584
rect 182836 281518 182864 306575
rect 182914 291952 182970 291961
rect 182914 291887 182970 291896
rect 182928 283529 182956 291887
rect 182914 283520 182970 283529
rect 182914 283455 182970 283464
rect 182824 281512 182876 281518
rect 182824 281454 182876 281460
rect 182824 256216 182876 256222
rect 182824 256158 182876 256164
rect 182086 247480 182142 247489
rect 182086 247415 182142 247424
rect 182088 242956 182140 242962
rect 182088 242898 182140 242904
rect 181534 241088 181590 241097
rect 181534 241023 181590 241032
rect 181534 231160 181590 231169
rect 181534 231095 181590 231104
rect 181548 204921 181576 231095
rect 181534 204912 181590 204921
rect 181534 204847 181590 204856
rect 181548 97986 181576 204847
rect 181996 101448 182048 101454
rect 181996 101390 182048 101396
rect 182008 100774 182036 101390
rect 181996 100768 182048 100774
rect 181996 100710 182048 100716
rect 181536 97980 181588 97986
rect 181536 97922 181588 97928
rect 181442 77888 181498 77897
rect 181442 77823 181498 77832
rect 182008 60042 182036 100710
rect 182100 95198 182128 242898
rect 182546 236056 182602 236065
rect 182546 235991 182602 236000
rect 182560 231130 182588 235991
rect 182548 231124 182600 231130
rect 182548 231066 182600 231072
rect 182836 213926 182864 256158
rect 182916 247104 182968 247110
rect 182916 247046 182968 247052
rect 182928 237969 182956 247046
rect 183388 240106 183416 351047
rect 183480 300830 183508 437446
rect 184308 431954 184336 443702
rect 184572 443692 184624 443698
rect 184572 443634 184624 443640
rect 184584 437510 184612 443634
rect 184572 437504 184624 437510
rect 184572 437446 184624 437452
rect 184216 431926 184336 431954
rect 184216 313410 184244 431926
rect 184296 409148 184348 409154
rect 184296 409090 184348 409096
rect 184308 373969 184336 409090
rect 184768 402286 184796 489126
rect 184860 449177 184888 615538
rect 187516 610088 187568 610094
rect 187516 610030 187568 610036
rect 185582 602032 185638 602041
rect 185582 601967 185638 601976
rect 185596 574802 185624 601967
rect 186962 600672 187018 600681
rect 186962 600607 187018 600616
rect 186976 587178 187004 600607
rect 186964 587172 187016 587178
rect 186964 587114 187016 587120
rect 187056 586560 187108 586566
rect 187056 586502 187108 586508
rect 186226 578368 186282 578377
rect 186226 578303 186282 578312
rect 185584 574796 185636 574802
rect 185584 574738 185636 574744
rect 185676 560448 185728 560454
rect 185676 560390 185728 560396
rect 185584 494828 185636 494834
rect 185584 494770 185636 494776
rect 184846 449168 184902 449177
rect 184846 449103 184848 449112
rect 184900 449103 184902 449112
rect 184848 449074 184900 449080
rect 184860 449043 184888 449074
rect 185596 407182 185624 494770
rect 185688 480865 185716 560390
rect 186240 511290 186268 578303
rect 186964 578264 187016 578270
rect 186964 578206 187016 578212
rect 186976 567866 187004 578206
rect 187068 577522 187096 586502
rect 187056 577516 187108 577522
rect 187056 577458 187108 577464
rect 186964 567860 187016 567866
rect 186964 567802 187016 567808
rect 187330 555248 187386 555257
rect 187330 555183 187386 555192
rect 187344 523802 187372 555183
rect 187424 547936 187476 547942
rect 187424 547878 187476 547884
rect 187332 523796 187384 523802
rect 187332 523738 187384 523744
rect 186228 511284 186280 511290
rect 186228 511226 186280 511232
rect 186964 498908 187016 498914
rect 186964 498850 187016 498856
rect 185674 480856 185730 480865
rect 185674 480791 185730 480800
rect 186226 475416 186282 475425
rect 186226 475351 186282 475360
rect 186044 472048 186096 472054
rect 186044 471990 186096 471996
rect 186056 438938 186084 471990
rect 186134 449440 186190 449449
rect 186134 449375 186190 449384
rect 186044 438932 186096 438938
rect 186044 438874 186096 438880
rect 186148 407794 186176 449375
rect 186136 407788 186188 407794
rect 186136 407730 186188 407736
rect 185584 407176 185636 407182
rect 185584 407118 185636 407124
rect 184756 402280 184808 402286
rect 184756 402222 184808 402228
rect 184768 401742 184796 402222
rect 184756 401736 184808 401742
rect 184756 401678 184808 401684
rect 184938 390688 184994 390697
rect 184938 390623 184994 390632
rect 184952 389881 184980 390623
rect 184938 389872 184994 389881
rect 184938 389807 184994 389816
rect 184848 388476 184900 388482
rect 184848 388418 184900 388424
rect 184860 387734 184888 388418
rect 184388 387728 184440 387734
rect 184388 387670 184440 387676
rect 184848 387728 184900 387734
rect 184848 387670 184900 387676
rect 184294 373960 184350 373969
rect 184294 373895 184350 373904
rect 184400 354674 184428 387670
rect 185596 385014 185624 407118
rect 186136 406020 186188 406026
rect 186136 405962 186188 405968
rect 185584 385008 185636 385014
rect 185584 384950 185636 384956
rect 184308 354646 184428 354674
rect 184308 353258 184336 354646
rect 184296 353252 184348 353258
rect 184296 353194 184348 353200
rect 184204 313404 184256 313410
rect 184204 313346 184256 313352
rect 183468 300824 183520 300830
rect 183468 300766 183520 300772
rect 184216 287706 184244 313346
rect 184204 287700 184256 287706
rect 184204 287642 184256 287648
rect 184308 280294 184336 353194
rect 184846 345672 184902 345681
rect 184846 345607 184902 345616
rect 184860 294710 184888 345607
rect 185584 320204 185636 320210
rect 185584 320146 185636 320152
rect 184848 294704 184900 294710
rect 184848 294646 184900 294652
rect 184860 294030 184888 294646
rect 184848 294024 184900 294030
rect 184848 293966 184900 293972
rect 184756 287768 184808 287774
rect 184756 287710 184808 287716
rect 184296 280288 184348 280294
rect 184296 280230 184348 280236
rect 183468 278044 183520 278050
rect 183468 277986 183520 277992
rect 183480 277438 183508 277986
rect 183468 277432 183520 277438
rect 183468 277374 183520 277380
rect 183480 243574 183508 277374
rect 184204 275324 184256 275330
rect 184204 275266 184256 275272
rect 184216 269414 184244 275266
rect 184204 269408 184256 269414
rect 184204 269350 184256 269356
rect 183468 243568 183520 243574
rect 183468 243510 183520 243516
rect 183376 240100 183428 240106
rect 183376 240042 183428 240048
rect 182914 237960 182970 237969
rect 182914 237895 182970 237904
rect 182916 224324 182968 224330
rect 182916 224266 182968 224272
rect 182928 218006 182956 224266
rect 182916 218000 182968 218006
rect 182916 217942 182968 217948
rect 182824 213920 182876 213926
rect 182824 213862 182876 213868
rect 183468 213920 183520 213926
rect 183468 213862 183520 213868
rect 182824 178696 182876 178702
rect 182824 178638 182876 178644
rect 182836 158030 182864 178638
rect 182824 158024 182876 158030
rect 182824 157966 182876 157972
rect 182836 126886 182864 157966
rect 182914 143712 182970 143721
rect 182914 143647 182970 143656
rect 182928 135250 182956 143647
rect 182916 135244 182968 135250
rect 182916 135186 182968 135192
rect 182824 126880 182876 126886
rect 182824 126822 182876 126828
rect 183376 113824 183428 113830
rect 183376 113766 183428 113772
rect 183388 113218 183416 113766
rect 183376 113212 183428 113218
rect 183376 113154 183428 113160
rect 182088 95192 182140 95198
rect 182088 95134 182140 95140
rect 182100 94518 182128 95134
rect 182088 94512 182140 94518
rect 182088 94454 182140 94460
rect 181996 60036 182048 60042
rect 181996 59978 182048 59984
rect 183388 29646 183416 113154
rect 183480 108934 183508 213862
rect 184216 144226 184244 269350
rect 184308 242962 184336 280230
rect 184388 254584 184440 254590
rect 184388 254526 184440 254532
rect 184296 242956 184348 242962
rect 184296 242898 184348 242904
rect 184400 225690 184428 254526
rect 184768 229770 184796 287710
rect 185596 287026 185624 320146
rect 185674 309496 185730 309505
rect 185674 309431 185730 309440
rect 185688 299470 185716 309431
rect 185676 299464 185728 299470
rect 185676 299406 185728 299412
rect 186042 290456 186098 290465
rect 186042 290391 186098 290400
rect 186056 290018 186084 290391
rect 186044 290012 186096 290018
rect 186044 289954 186096 289960
rect 185584 287020 185636 287026
rect 185584 286962 185636 286968
rect 184940 265668 184992 265674
rect 184940 265610 184992 265616
rect 184846 240816 184902 240825
rect 184846 240751 184902 240760
rect 184756 229764 184808 229770
rect 184756 229706 184808 229712
rect 184388 225684 184440 225690
rect 184388 225626 184440 225632
rect 184296 147688 184348 147694
rect 184296 147630 184348 147636
rect 184204 144220 184256 144226
rect 184204 144162 184256 144168
rect 184204 135312 184256 135318
rect 184204 135254 184256 135260
rect 183468 108928 183520 108934
rect 183468 108870 183520 108876
rect 183560 93152 183612 93158
rect 183560 93094 183612 93100
rect 183572 60625 183600 93094
rect 183558 60616 183614 60625
rect 183558 60551 183614 60560
rect 179420 29640 179472 29646
rect 179420 29582 179472 29588
rect 183376 29640 183428 29646
rect 183376 29582 183428 29588
rect 178684 18624 178736 18630
rect 178684 18566 178736 18572
rect 168380 8968 168432 8974
rect 168380 8910 168432 8916
rect 152556 4820 152608 4826
rect 152556 4762 152608 4768
rect 150624 3664 150676 3670
rect 150624 3606 150676 3612
rect 152464 3664 152516 3670
rect 152464 3606 152516 3612
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144736 3528 144788 3534
rect 144736 3470 144788 3476
rect 147126 3496 147182 3505
rect 140044 3460 140096 3466
rect 140044 3402 140096 3408
rect 137284 2168 137336 2174
rect 137284 2110 137336 2116
rect 140056 480 140084 3402
rect 143552 480 143580 3470
rect 147126 3431 147182 3440
rect 147140 480 147168 3431
rect 150636 480 150664 3606
rect 184216 3466 184244 135254
rect 184308 120086 184336 147630
rect 184386 143576 184442 143585
rect 184386 143511 184442 143520
rect 184400 133210 184428 143511
rect 184388 133204 184440 133210
rect 184388 133146 184440 133152
rect 184754 120728 184810 120737
rect 184754 120663 184756 120672
rect 184808 120663 184810 120672
rect 184756 120634 184808 120640
rect 184296 120080 184348 120086
rect 184296 120022 184348 120028
rect 184296 102196 184348 102202
rect 184296 102138 184348 102144
rect 184308 92478 184336 102138
rect 184388 98116 184440 98122
rect 184388 98058 184440 98064
rect 184296 92472 184348 92478
rect 184296 92414 184348 92420
rect 184400 92342 184428 98058
rect 184860 92721 184888 240751
rect 184846 92712 184902 92721
rect 184846 92647 184902 92656
rect 184388 92336 184440 92342
rect 184388 92278 184440 92284
rect 184952 72486 184980 265610
rect 185492 257372 185544 257378
rect 185492 257314 185544 257320
rect 185504 248414 185532 257314
rect 185582 257272 185638 257281
rect 185582 257207 185584 257216
rect 185636 257207 185638 257216
rect 185584 257178 185636 257184
rect 186056 252550 186084 289954
rect 186148 267034 186176 405962
rect 186240 302569 186268 475351
rect 186976 440298 187004 498850
rect 187436 496194 187464 547878
rect 187528 510950 187556 610030
rect 188344 607300 188396 607306
rect 188344 607242 188396 607248
rect 187606 599584 187662 599593
rect 187606 599519 187662 599528
rect 187620 599010 187648 599519
rect 187608 599004 187660 599010
rect 187608 598946 187660 598952
rect 187516 510944 187568 510950
rect 187516 510886 187568 510892
rect 187424 496188 187476 496194
rect 187424 496130 187476 496136
rect 187516 487824 187568 487830
rect 187516 487766 187568 487772
rect 187146 468616 187202 468625
rect 187146 468551 187202 468560
rect 187056 454096 187108 454102
rect 187056 454038 187108 454044
rect 186964 440292 187016 440298
rect 186964 440234 187016 440240
rect 186964 439000 187016 439006
rect 186964 438942 187016 438948
rect 186976 420238 187004 438942
rect 186964 420232 187016 420238
rect 186964 420174 187016 420180
rect 187068 406026 187096 454038
rect 187160 443698 187188 468551
rect 187528 456142 187556 487766
rect 187620 458561 187648 598946
rect 188356 585041 188384 607242
rect 188342 585032 188398 585041
rect 188342 584967 188398 584976
rect 188344 579760 188396 579766
rect 188344 579702 188396 579708
rect 188356 571334 188384 579702
rect 188344 571328 188396 571334
rect 188344 571270 188396 571276
rect 188804 567248 188856 567254
rect 188804 567190 188856 567196
rect 187700 565820 187752 565826
rect 187700 565762 187752 565768
rect 187712 565146 187740 565762
rect 187700 565140 187752 565146
rect 187700 565082 187752 565088
rect 187700 564460 187752 564466
rect 187700 564402 187752 564408
rect 187712 558210 187740 564402
rect 187700 558204 187752 558210
rect 187700 558146 187752 558152
rect 188344 557660 188396 557666
rect 188344 557602 188396 557608
rect 188356 554878 188384 557602
rect 188344 554872 188396 554878
rect 188344 554814 188396 554820
rect 188344 549364 188396 549370
rect 188344 549306 188396 549312
rect 187700 549296 187752 549302
rect 187700 549238 187752 549244
rect 187712 548554 187740 549238
rect 187700 548548 187752 548554
rect 187700 548490 187752 548496
rect 188356 540258 188384 549306
rect 188436 545760 188488 545766
rect 188436 545702 188488 545708
rect 188344 540252 188396 540258
rect 188344 540194 188396 540200
rect 188448 537985 188476 545702
rect 188434 537976 188490 537985
rect 188434 537911 188490 537920
rect 188342 536072 188398 536081
rect 188342 536007 188398 536016
rect 187700 533384 187752 533390
rect 187700 533326 187752 533332
rect 187712 532710 187740 533326
rect 187700 532704 187752 532710
rect 187700 532646 187752 532652
rect 188356 511329 188384 536007
rect 188342 511320 188398 511329
rect 188342 511255 188398 511264
rect 188344 466472 188396 466478
rect 188344 466414 188396 466420
rect 188160 460964 188212 460970
rect 188160 460906 188212 460912
rect 187792 459536 187844 459542
rect 187792 459478 187844 459484
rect 187606 458552 187662 458561
rect 187606 458487 187662 458496
rect 187620 457502 187648 458487
rect 187804 458289 187832 459478
rect 187790 458280 187846 458289
rect 187700 458244 187752 458250
rect 187790 458215 187846 458224
rect 187700 458186 187752 458192
rect 187608 457496 187660 457502
rect 187608 457438 187660 457444
rect 187516 456136 187568 456142
rect 187516 456078 187568 456084
rect 187712 456074 187740 458186
rect 188172 457502 188200 460906
rect 188356 460329 188384 466414
rect 188342 460320 188398 460329
rect 188342 460255 188398 460264
rect 188160 457496 188212 457502
rect 188160 457438 188212 457444
rect 188344 456136 188396 456142
rect 188344 456078 188396 456084
rect 187700 456068 187752 456074
rect 187700 456010 187752 456016
rect 187606 446448 187662 446457
rect 187606 446383 187662 446392
rect 187148 443692 187200 443698
rect 187148 443634 187200 443640
rect 187056 406020 187108 406026
rect 187056 405962 187108 405968
rect 187620 402974 187648 446383
rect 187700 438932 187752 438938
rect 187700 438874 187752 438880
rect 187436 402946 187648 402974
rect 186964 401736 187016 401742
rect 186964 401678 187016 401684
rect 186320 392012 186372 392018
rect 186320 391954 186372 391960
rect 186332 390969 186360 391954
rect 186318 390960 186374 390969
rect 186318 390895 186374 390904
rect 186976 383081 187004 401678
rect 187436 387802 187464 402946
rect 187712 393314 187740 438874
rect 188356 436150 188384 456078
rect 188436 454164 188488 454170
rect 188436 454106 188488 454112
rect 188448 447914 188476 454106
rect 188816 450634 188844 567190
rect 188908 565826 188936 702850
rect 189722 612776 189778 612785
rect 189722 612711 189778 612720
rect 188988 611448 189040 611454
rect 188988 611390 189040 611396
rect 188896 565820 188948 565826
rect 188896 565762 188948 565768
rect 188804 450628 188856 450634
rect 188804 450570 188856 450576
rect 188816 449954 188844 450570
rect 188804 449948 188856 449954
rect 188804 449890 188856 449896
rect 188436 447908 188488 447914
rect 188436 447850 188488 447856
rect 188344 436144 188396 436150
rect 188344 436086 188396 436092
rect 188356 429894 188384 436086
rect 188344 429888 188396 429894
rect 188344 429830 188396 429836
rect 188344 398880 188396 398886
rect 188344 398822 188396 398828
rect 187976 393984 188028 393990
rect 187976 393926 188028 393932
rect 187528 393286 187740 393314
rect 187424 387796 187476 387802
rect 187424 387738 187476 387744
rect 187148 387116 187200 387122
rect 187148 387058 187200 387064
rect 187054 387016 187110 387025
rect 187054 386951 187110 386960
rect 186962 383072 187018 383081
rect 186962 383007 187018 383016
rect 187068 371890 187096 386951
rect 187160 373998 187188 387058
rect 187148 373992 187200 373998
rect 187148 373934 187200 373940
rect 187160 373454 187188 373934
rect 187148 373448 187200 373454
rect 187148 373390 187200 373396
rect 187056 371884 187108 371890
rect 187056 371826 187108 371832
rect 187528 334626 187556 393286
rect 187606 390552 187662 390561
rect 187662 390510 187740 390538
rect 187606 390487 187662 390496
rect 187712 386209 187740 390510
rect 187988 389230 188016 393926
rect 187976 389224 188028 389230
rect 187976 389166 188028 389172
rect 187698 386200 187754 386209
rect 187698 386135 187754 386144
rect 187700 380248 187752 380254
rect 187700 380190 187752 380196
rect 187712 378826 187740 380190
rect 187700 378820 187752 378826
rect 187700 378762 187752 378768
rect 188356 375329 188384 398822
rect 188526 394088 188582 394097
rect 188526 394023 188582 394032
rect 188540 387802 188568 394023
rect 189000 393314 189028 611390
rect 189736 597650 189764 612711
rect 201512 609278 201540 702918
rect 218992 702846 219020 703520
rect 218980 702840 219032 702846
rect 218980 702782 219032 702788
rect 224224 702772 224276 702778
rect 224224 702714 224276 702720
rect 206284 702704 206336 702710
rect 206284 702646 206336 702652
rect 206296 619614 206324 702646
rect 215300 702636 215352 702642
rect 215300 702578 215352 702584
rect 222844 702636 222896 702642
rect 222844 702578 222896 702584
rect 205640 619608 205692 619614
rect 205640 619550 205692 619556
rect 206284 619608 206336 619614
rect 206284 619550 206336 619556
rect 205652 618322 205680 619550
rect 205640 618316 205692 618322
rect 205640 618258 205692 618264
rect 205652 615494 205680 618258
rect 213920 615528 213972 615534
rect 205652 615466 206416 615494
rect 213972 615476 214696 615494
rect 213920 615470 214696 615476
rect 213932 615466 214696 615470
rect 204350 611416 204406 611425
rect 204350 611351 204406 611360
rect 202878 610056 202934 610065
rect 202878 609991 202934 610000
rect 201500 609272 201552 609278
rect 201500 609214 201552 609220
rect 198738 608696 198794 608705
rect 198738 608631 198794 608640
rect 200672 608660 200724 608666
rect 191654 607880 191710 607889
rect 191654 607815 191710 607824
rect 191194 603664 191250 603673
rect 191194 603599 191250 603608
rect 191102 599040 191158 599049
rect 191102 598975 191158 598984
rect 189724 597644 189776 597650
rect 189724 597586 189776 597592
rect 189080 542428 189132 542434
rect 189080 542370 189132 542376
rect 189092 538354 189120 542370
rect 189080 538348 189132 538354
rect 189080 538290 189132 538296
rect 189736 469305 189764 597586
rect 190642 596320 190698 596329
rect 190642 596255 190698 596264
rect 190656 596174 190684 596255
rect 190564 596146 190684 596174
rect 190564 589966 190592 596146
rect 190642 595232 190698 595241
rect 190642 595167 190698 595176
rect 190656 594930 190684 595167
rect 190644 594924 190696 594930
rect 190644 594866 190696 594872
rect 191010 591288 191066 591297
rect 191010 591223 191066 591232
rect 191024 590714 191052 591223
rect 191012 590708 191064 590714
rect 191012 590650 191064 590656
rect 190552 589960 190604 589966
rect 190552 589902 190604 589908
rect 190460 586560 190512 586566
rect 190458 586528 190460 586537
rect 190512 586528 190514 586537
rect 190458 586463 190514 586472
rect 191116 578377 191144 598975
rect 191208 586634 191236 603599
rect 191668 596873 191696 607815
rect 196716 607300 196768 607306
rect 196716 607242 196768 607248
rect 196728 604761 196756 607242
rect 196714 604752 196770 604761
rect 196714 604687 196770 604696
rect 191748 601792 191800 601798
rect 191748 601734 191800 601740
rect 191760 598913 191788 601734
rect 192576 600432 192628 600438
rect 192576 600374 192628 600380
rect 194690 600400 194746 600409
rect 192484 599208 192536 599214
rect 192484 599150 192536 599156
rect 191746 598904 191802 598913
rect 191746 598839 191802 598848
rect 191654 596864 191710 596873
rect 191654 596799 191710 596808
rect 191748 594856 191800 594862
rect 191748 594798 191800 594804
rect 191760 594697 191788 594798
rect 191746 594688 191802 594697
rect 191746 594623 191802 594632
rect 191654 593464 191710 593473
rect 191654 593399 191710 593408
rect 191286 589384 191342 589393
rect 191286 589319 191342 589328
rect 191196 586628 191248 586634
rect 191196 586570 191248 586576
rect 191208 586265 191236 586570
rect 191194 586256 191250 586265
rect 191194 586191 191250 586200
rect 191300 583030 191328 589319
rect 191288 583024 191340 583030
rect 191288 582966 191340 582972
rect 191102 578368 191158 578377
rect 191102 578303 191158 578312
rect 191562 578368 191618 578377
rect 191562 578303 191618 578312
rect 191576 578270 191604 578303
rect 191564 578264 191616 578270
rect 191564 578206 191616 578212
rect 191010 576192 191066 576201
rect 191010 576127 191066 576136
rect 191024 575618 191052 576127
rect 191194 575648 191250 575657
rect 191012 575612 191064 575618
rect 191194 575583 191250 575592
rect 191012 575554 191064 575560
rect 191208 575550 191236 575583
rect 191196 575544 191248 575550
rect 191196 575486 191248 575492
rect 191286 574560 191342 574569
rect 191286 574495 191342 574504
rect 191300 574122 191328 574495
rect 191288 574116 191340 574122
rect 191288 574058 191340 574064
rect 191010 573336 191066 573345
rect 191010 573271 191066 573280
rect 191024 572830 191052 573271
rect 191012 572824 191064 572830
rect 191012 572766 191064 572772
rect 191562 572792 191618 572801
rect 191562 572727 191564 572736
rect 191616 572727 191618 572736
rect 191564 572698 191616 572704
rect 191288 572688 191340 572694
rect 191288 572630 191340 572636
rect 191300 572257 191328 572630
rect 191286 572248 191342 572257
rect 191286 572183 191342 572192
rect 190920 571328 190972 571334
rect 190920 571270 190972 571276
rect 190932 570625 190960 571270
rect 191562 570888 191618 570897
rect 191562 570823 191618 570832
rect 191576 570654 191604 570823
rect 191564 570648 191616 570654
rect 190918 570616 190974 570625
rect 191564 570590 191616 570596
rect 190918 570551 190974 570560
rect 190366 568712 190422 568721
rect 190366 568647 190422 568656
rect 189816 536104 189868 536110
rect 189816 536046 189868 536052
rect 189828 518226 189856 536046
rect 190380 530602 190408 568647
rect 190458 567624 190514 567633
rect 190458 567559 190514 567568
rect 190472 565049 190500 567559
rect 190828 565820 190880 565826
rect 190828 565762 190880 565768
rect 190458 565040 190514 565049
rect 190458 564975 190514 564984
rect 190840 564777 190868 565762
rect 191102 564904 191158 564913
rect 191102 564839 191158 564848
rect 190826 564768 190882 564777
rect 190826 564703 190882 564712
rect 191116 564466 191144 564839
rect 191104 564460 191156 564466
rect 191104 564402 191156 564408
rect 191012 563712 191064 563718
rect 191010 563680 191012 563689
rect 191064 563680 191066 563689
rect 191010 563615 191066 563624
rect 191194 560960 191250 560969
rect 191194 560895 191250 560904
rect 191102 560688 191158 560697
rect 191102 560623 191158 560632
rect 191116 560454 191144 560623
rect 191104 560448 191156 560454
rect 191104 560390 191156 560396
rect 191208 560318 191236 560895
rect 191196 560312 191248 560318
rect 191196 560254 191248 560260
rect 190918 558240 190974 558249
rect 190918 558175 190974 558184
rect 190932 557666 190960 558175
rect 190920 557660 190972 557666
rect 190920 557602 190972 557608
rect 191668 557534 191696 593399
rect 191746 592376 191802 592385
rect 191746 592311 191802 592320
rect 191760 592142 191788 592311
rect 191748 592136 191800 592142
rect 191748 592078 191800 592084
rect 192496 591326 192524 599150
rect 192588 592686 192616 600374
rect 194690 600335 194746 600344
rect 192758 599312 192814 599321
rect 192758 599247 192814 599256
rect 192668 599004 192720 599010
rect 192668 598946 192720 598952
rect 192680 594114 192708 598946
rect 192772 594182 192800 599247
rect 194704 599148 194732 600335
rect 196728 599148 196756 604687
rect 198554 600536 198610 600545
rect 198554 600471 198610 600480
rect 197358 600400 197414 600409
rect 197358 600335 197414 600344
rect 193404 599140 193456 599146
rect 193404 599082 193456 599088
rect 192944 598936 192996 598942
rect 192944 598878 192996 598884
rect 192956 597582 192984 598878
rect 193312 598868 193364 598874
rect 193312 598810 193364 598816
rect 193324 597825 193352 598810
rect 193310 597816 193366 597825
rect 193310 597751 193366 597760
rect 192944 597576 192996 597582
rect 192944 597518 192996 597524
rect 192760 594176 192812 594182
rect 192760 594118 192812 594124
rect 192668 594108 192720 594114
rect 192668 594050 192720 594056
rect 193416 592793 193444 599082
rect 197174 599040 197230 599049
rect 193508 598998 194166 599026
rect 195072 598998 195454 599026
rect 195624 599010 196006 599026
rect 195612 599004 196006 599010
rect 193508 598505 193536 598998
rect 195072 598942 195100 598998
rect 195664 598998 196006 599004
rect 197230 598998 197294 599026
rect 197174 598975 197230 598984
rect 195612 598946 195664 598952
rect 197372 598942 197400 600335
rect 197636 599208 197688 599214
rect 197688 599156 198030 599162
rect 197636 599150 198030 599156
rect 197648 599134 198030 599150
rect 198568 599148 198596 600471
rect 198752 599162 198780 608631
rect 200672 608602 200724 608608
rect 199842 604616 199898 604625
rect 199842 604551 199898 604560
rect 198752 599134 199134 599162
rect 199856 599148 199884 604551
rect 200396 600364 200448 600370
rect 200396 600306 200448 600312
rect 200408 599148 200436 600306
rect 200684 599162 200712 608602
rect 201682 600400 201738 600409
rect 201682 600335 201738 600344
rect 200684 599134 201158 599162
rect 201696 599148 201724 600335
rect 202892 599162 202920 609991
rect 203708 603152 203760 603158
rect 203708 603094 203760 603100
rect 202892 599134 202998 599162
rect 203720 599148 203748 603094
rect 204260 600432 204312 600438
rect 204260 600374 204312 600380
rect 204272 599148 204300 600374
rect 204364 599162 204392 611351
rect 206100 604580 206152 604586
rect 206100 604522 206152 604528
rect 204364 599134 204838 599162
rect 206112 599148 206140 604522
rect 206388 599162 206416 615466
rect 207664 614236 207716 614242
rect 207664 614178 207716 614184
rect 207676 599162 207704 614178
rect 209412 607232 209464 607238
rect 209412 607174 209464 607180
rect 208674 603256 208730 603265
rect 208674 603191 208730 603200
rect 206388 599134 206862 599162
rect 207676 599134 208150 599162
rect 208688 599148 208716 603191
rect 209424 599148 209452 607174
rect 214380 605872 214432 605878
rect 214380 605814 214432 605820
rect 211618 602032 211674 602041
rect 211618 601967 211674 601976
rect 211632 601769 211660 601967
rect 211618 601760 211674 601769
rect 211252 601724 211304 601730
rect 211618 601695 211674 601704
rect 211252 601666 211304 601672
rect 209962 600536 210018 600545
rect 209962 600471 210018 600480
rect 209976 599148 210004 600471
rect 211264 599148 211292 601666
rect 211632 599162 211660 601695
rect 212538 599312 212594 599321
rect 212538 599247 212594 599256
rect 211632 599134 211830 599162
rect 212552 599148 212580 599247
rect 213366 599176 213422 599185
rect 213118 599134 213366 599162
rect 214392 599148 214420 605814
rect 214668 599162 214696 615466
rect 215312 600409 215340 702578
rect 219440 616888 219492 616894
rect 219440 616830 219492 616836
rect 219452 615494 219480 616830
rect 219452 615466 219664 615494
rect 217232 610088 217284 610094
rect 217232 610030 217284 610036
rect 215668 606484 215720 606490
rect 215668 606426 215720 606432
rect 215680 605946 215708 606426
rect 215668 605940 215720 605946
rect 215668 605882 215720 605888
rect 215298 600400 215354 600409
rect 215298 600335 215354 600344
rect 214668 599134 215142 599162
rect 215680 599148 215708 605882
rect 216956 604512 217008 604518
rect 216956 604454 217008 604460
rect 216402 600400 216458 600409
rect 216402 600335 216458 600344
rect 216680 600364 216732 600370
rect 216416 599148 216444 600335
rect 216680 600306 216732 600312
rect 213366 599111 213422 599120
rect 216692 599049 216720 600306
rect 216968 599148 216996 604454
rect 217244 599162 217272 610030
rect 218242 609240 218298 609249
rect 218242 609175 218298 609184
rect 218256 599593 218284 609175
rect 219530 600808 219586 600817
rect 219530 600743 219586 600752
rect 218242 599584 218298 599593
rect 218242 599519 218298 599528
rect 217244 599134 217718 599162
rect 218256 599148 218284 599519
rect 219544 599148 219572 600743
rect 219636 599162 219664 615466
rect 221648 612876 221700 612882
rect 221648 612818 221700 612824
rect 221370 600808 221426 600817
rect 221370 600743 221426 600752
rect 219636 599134 220110 599162
rect 221384 599148 221412 600743
rect 221660 599162 221688 612818
rect 222856 612785 222884 702578
rect 222198 612776 222254 612785
rect 222198 612711 222254 612720
rect 222842 612776 222898 612785
rect 222842 612711 222898 612720
rect 222212 602206 222240 612711
rect 222292 609272 222344 609278
rect 222292 609214 222344 609220
rect 222200 602200 222252 602206
rect 222200 602142 222252 602148
rect 222304 600681 222332 609214
rect 223028 602200 223080 602206
rect 223028 602142 223080 602148
rect 222290 600672 222346 600681
rect 222290 600607 222346 600616
rect 222658 600672 222714 600681
rect 222658 600607 222714 600616
rect 221660 599134 222134 599162
rect 202602 599040 202658 599049
rect 202446 598998 202602 599026
rect 207110 599040 207166 599049
rect 205192 599010 205574 599026
rect 202602 598975 202658 598984
rect 205180 599004 205574 599010
rect 205232 598998 205574 599004
rect 210422 599040 210478 599049
rect 207166 598998 207414 599026
rect 207110 598975 207166 598984
rect 214010 599040 214066 599049
rect 210478 598998 210726 599026
rect 213854 598998 214010 599026
rect 210422 598975 210478 598984
rect 214010 598975 214066 598984
rect 216678 599040 216734 599049
rect 216678 598975 216734 598984
rect 218702 599040 218758 599049
rect 220910 599040 220966 599049
rect 218758 598998 218822 599026
rect 220846 598998 220910 599026
rect 218702 598975 218758 598984
rect 222672 599026 222700 600607
rect 223040 599162 223068 602142
rect 224236 601662 224264 702714
rect 233240 702568 233292 702574
rect 233240 702510 233292 702516
rect 233252 616010 233280 702510
rect 235184 702506 235212 703520
rect 242808 703180 242860 703186
rect 242808 703122 242860 703128
rect 235172 702500 235224 702506
rect 235172 702442 235224 702448
rect 241520 622464 241572 622470
rect 241520 622406 241572 622412
rect 236000 618384 236052 618390
rect 236000 618326 236052 618332
rect 233240 616004 233292 616010
rect 233240 615946 233292 615952
rect 233884 616004 233936 616010
rect 233884 615946 233936 615952
rect 233252 615602 233280 615946
rect 233240 615596 233292 615602
rect 233240 615538 233292 615544
rect 232320 614168 232372 614174
rect 232320 614110 232372 614116
rect 230480 611448 230532 611454
rect 230480 611390 230532 611396
rect 226340 608728 226392 608734
rect 226340 608670 226392 608676
rect 224224 601656 224276 601662
rect 224224 601598 224276 601604
rect 225236 601656 225288 601662
rect 225236 601598 225288 601604
rect 224222 599176 224278 599185
rect 223040 599134 223422 599162
rect 224278 599134 224526 599162
rect 225248 599148 225276 601598
rect 226352 599162 226380 608670
rect 229650 601896 229706 601905
rect 229650 601831 229706 601840
rect 227812 600364 227864 600370
rect 227812 600306 227864 600312
rect 226352 599134 226550 599162
rect 227824 599148 227852 600306
rect 228638 599176 228694 599185
rect 228390 599134 228638 599162
rect 224222 599111 224278 599120
rect 229664 599148 229692 601831
rect 230492 599162 230520 611390
rect 231490 600400 231546 600409
rect 231490 600335 231546 600344
rect 230492 599134 230966 599162
rect 231504 599148 231532 600335
rect 232332 599162 232360 614110
rect 233896 601594 233924 615946
rect 234066 607336 234122 607345
rect 234066 607271 234122 607280
rect 233884 601588 233936 601594
rect 233884 601530 233936 601536
rect 232332 599134 232806 599162
rect 234080 599148 234108 607271
rect 235356 601588 235408 601594
rect 235356 601530 235408 601536
rect 235368 599148 235396 601530
rect 236012 599162 236040 618326
rect 241532 615494 241560 622406
rect 241532 615466 241928 615494
rect 239218 606112 239274 606121
rect 239218 606047 239274 606056
rect 238482 604480 238538 604489
rect 238482 604415 238538 604424
rect 237562 600536 237618 600545
rect 237562 600471 237618 600480
rect 236642 600400 236698 600409
rect 236642 600335 236698 600344
rect 236012 599134 236118 599162
rect 236656 599148 236684 600335
rect 237576 599162 237604 600471
rect 237576 599134 237958 599162
rect 238496 599148 238524 604415
rect 239232 599148 239260 606047
rect 241796 604512 241848 604518
rect 241796 604454 241848 604460
rect 241060 603152 241112 603158
rect 241060 603094 241112 603100
rect 239772 600432 239824 600438
rect 239772 600374 239824 600380
rect 239784 599148 239812 600374
rect 241072 599148 241100 603094
rect 241808 599148 241836 604454
rect 241900 599162 241928 615466
rect 242820 604518 242848 703122
rect 248420 702772 248472 702778
rect 248420 702714 248472 702720
rect 242900 616956 242952 616962
rect 242900 616898 242952 616904
rect 242808 604512 242860 604518
rect 242808 604454 242860 604460
rect 242912 599162 242940 616898
rect 245474 605976 245530 605985
rect 245474 605911 245530 605920
rect 243634 600672 243690 600681
rect 243634 600607 243690 600616
rect 241900 599134 242374 599162
rect 242912 599134 243110 599162
rect 243648 599148 243676 600607
rect 244186 600536 244242 600545
rect 244186 600471 244242 600480
rect 244200 599148 244228 600471
rect 245488 599148 245516 605911
rect 246212 603220 246264 603226
rect 246212 603162 246264 603168
rect 246224 599148 246252 603162
rect 248432 599457 248460 702714
rect 255964 702500 256016 702506
rect 255964 702442 256016 702448
rect 251824 700324 251876 700330
rect 251824 700266 251876 700272
rect 251836 619682 251864 700266
rect 251180 619676 251232 619682
rect 251180 619618 251232 619624
rect 251824 619676 251876 619682
rect 251824 619618 251876 619624
rect 251192 615494 251220 619618
rect 251192 615466 251496 615494
rect 248786 600536 248842 600545
rect 248786 600471 248842 600480
rect 248418 599448 248474 599457
rect 248418 599383 248474 599392
rect 248800 599148 248828 600471
rect 250074 600400 250130 600409
rect 250074 600335 250130 600344
rect 251180 600364 251232 600370
rect 249338 599312 249394 599321
rect 249338 599247 249394 599256
rect 249352 599148 249380 599247
rect 250088 599148 250116 600335
rect 251180 600306 251232 600312
rect 251192 599148 251220 600306
rect 251468 599162 251496 615466
rect 254032 611380 254084 611386
rect 254032 611322 254084 611328
rect 252468 601724 252520 601730
rect 252468 601666 252520 601672
rect 251468 599134 251942 599162
rect 252480 599148 252508 601666
rect 253386 600536 253442 600545
rect 253386 600471 253442 600480
rect 228638 599111 228694 599120
rect 229008 599072 229060 599078
rect 224038 599040 224094 599049
rect 222672 599012 222976 599026
rect 222686 599010 222976 599012
rect 222686 599004 222988 599010
rect 222686 598998 222936 599004
rect 220910 598975 220966 598984
rect 205180 598946 205232 598952
rect 223974 598998 224038 599026
rect 226062 599040 226118 599049
rect 225814 598998 226062 599026
rect 224038 598975 224094 598984
rect 226062 598975 226118 598984
rect 226798 599040 226854 599049
rect 226854 598998 227102 599026
rect 247684 599072 247736 599078
rect 230018 599040 230074 599049
rect 229060 599020 229126 599026
rect 229008 599014 229126 599020
rect 229020 598998 229126 599014
rect 226798 598975 226854 598984
rect 232410 599040 232466 599049
rect 230074 598998 230414 599026
rect 232254 598998 232410 599026
rect 230018 598975 230074 598984
rect 232410 598975 232466 598984
rect 233238 599040 233294 599049
rect 234710 599040 234766 599049
rect 233294 598998 233542 599026
rect 233238 598975 233294 598984
rect 236826 599040 236882 599049
rect 234766 598998 234830 599026
rect 234710 598975 234766 598984
rect 240690 599040 240746 599049
rect 236882 598998 237222 599026
rect 240534 598998 240690 599026
rect 236826 598975 236882 598984
rect 244950 598998 245240 599026
rect 247526 599020 247684 599026
rect 247526 599014 247736 599020
rect 247774 599040 247830 599049
rect 247526 598998 247724 599014
rect 240690 598975 240746 598984
rect 222936 598946 222988 598952
rect 245212 598942 245240 598998
rect 250902 599040 250958 599049
rect 247830 598998 248078 599026
rect 250654 598998 250902 599026
rect 247774 598975 247830 598984
rect 250902 598975 250958 598984
rect 252834 599040 252890 599049
rect 252890 598998 253230 599026
rect 252834 598975 252890 598984
rect 195060 598936 195112 598942
rect 195060 598878 195112 598884
rect 197360 598936 197412 598942
rect 197360 598878 197412 598884
rect 245200 598936 245252 598942
rect 245200 598878 245252 598884
rect 193494 598496 193550 598505
rect 246776 598466 246804 598468
rect 193494 598431 193550 598440
rect 246764 598460 246816 598466
rect 246764 598402 246816 598408
rect 253400 596834 253428 600471
rect 253478 600400 253534 600409
rect 253478 600335 253534 600344
rect 253388 596828 253440 596834
rect 253388 596770 253440 596776
rect 193402 592784 193458 592793
rect 193402 592719 193458 592728
rect 192576 592680 192628 592686
rect 192576 592622 192628 592628
rect 253386 592104 253442 592113
rect 253386 592039 253442 592048
rect 192484 591320 192536 591326
rect 192484 591262 192536 591268
rect 253400 586514 253428 592039
rect 253492 591326 253520 600335
rect 253570 599312 253626 599321
rect 253570 599247 253626 599256
rect 253584 599049 253612 599247
rect 253570 599040 253626 599049
rect 253570 598975 253626 598984
rect 253480 591320 253532 591326
rect 253480 591262 253532 591268
rect 253938 587412 253994 587421
rect 253938 587347 253994 587356
rect 253308 586486 253428 586514
rect 191748 585200 191800 585206
rect 191746 585168 191748 585177
rect 191800 585168 191802 585177
rect 191746 585103 191802 585112
rect 191746 583944 191802 583953
rect 191746 583879 191802 583888
rect 191760 583846 191788 583879
rect 191748 583840 191800 583846
rect 191748 583782 191800 583788
rect 191746 582720 191802 582729
rect 191746 582655 191802 582664
rect 191760 582418 191788 582655
rect 191748 582412 191800 582418
rect 191748 582354 191800 582360
rect 191746 581632 191802 581641
rect 191746 581567 191802 581576
rect 191760 581058 191788 581567
rect 191748 581052 191800 581058
rect 191748 580994 191800 581000
rect 191746 578912 191802 578921
rect 191746 578847 191802 578856
rect 191760 578354 191788 578847
rect 191760 578326 191880 578354
rect 191748 578196 191800 578202
rect 191748 578138 191800 578144
rect 191760 578105 191788 578138
rect 191746 578096 191802 578105
rect 191746 578031 191802 578040
rect 191852 577946 191880 578326
rect 191760 577918 191880 577946
rect 191760 567338 191788 577918
rect 191760 567310 191880 567338
rect 191748 567248 191800 567254
rect 191746 567216 191748 567225
rect 191800 567216 191802 567225
rect 191746 567151 191802 567160
rect 191746 562048 191802 562057
rect 191746 561983 191802 561992
rect 191760 561746 191788 561983
rect 191748 561740 191800 561746
rect 191748 561682 191800 561688
rect 191746 557832 191802 557841
rect 191746 557767 191802 557776
rect 191760 557598 191788 557767
rect 191748 557592 191800 557598
rect 191748 557534 191800 557540
rect 191484 557506 191696 557534
rect 190826 554840 190882 554849
rect 190826 554775 190828 554784
rect 190880 554775 190882 554784
rect 190828 554746 190880 554752
rect 190918 553888 190974 553897
rect 190918 553823 190974 553832
rect 190932 553450 190960 553823
rect 190920 553444 190972 553450
rect 190920 553386 190972 553392
rect 191378 550760 191434 550769
rect 191378 550695 191434 550704
rect 191392 550662 191420 550695
rect 191380 550656 191432 550662
rect 191380 550598 191432 550604
rect 191484 548978 191512 557506
rect 191746 556472 191802 556481
rect 191746 556407 191802 556416
rect 191760 556238 191788 556407
rect 191748 556232 191800 556238
rect 191748 556174 191800 556180
rect 191746 552120 191802 552129
rect 191746 552055 191748 552064
rect 191800 552055 191802 552064
rect 191748 552026 191800 552032
rect 191562 549808 191618 549817
rect 191562 549743 191618 549752
rect 191576 549114 191604 549743
rect 191746 549400 191802 549409
rect 191746 549335 191802 549344
rect 191760 549302 191788 549335
rect 191748 549296 191800 549302
rect 191748 549238 191800 549244
rect 191576 549086 191788 549114
rect 191484 548950 191696 548978
rect 191562 548040 191618 548049
rect 191562 547975 191618 547984
rect 191576 547942 191604 547975
rect 191564 547936 191616 547942
rect 191564 547878 191616 547884
rect 191286 547088 191342 547097
rect 191286 547023 191342 547032
rect 191300 546514 191328 547023
rect 191564 546576 191616 546582
rect 191562 546544 191564 546553
rect 191616 546544 191618 546553
rect 191288 546508 191340 546514
rect 191562 546479 191618 546488
rect 191288 546450 191340 546456
rect 191194 545456 191250 545465
rect 191194 545391 191250 545400
rect 191208 545154 191236 545391
rect 191196 545148 191248 545154
rect 191196 545090 191248 545096
rect 190644 545080 190696 545086
rect 190644 545022 190696 545028
rect 190656 544105 190684 545022
rect 191102 544232 191158 544241
rect 191102 544167 191158 544176
rect 190642 544096 190698 544105
rect 190642 544031 190698 544040
rect 191116 543794 191144 544167
rect 191104 543788 191156 543794
rect 191104 543730 191156 543736
rect 191562 542600 191618 542609
rect 191562 542535 191618 542544
rect 191576 542502 191604 542535
rect 191564 542496 191616 542502
rect 191564 542438 191616 542444
rect 190826 541512 190882 541521
rect 190826 541447 190882 541456
rect 190840 541006 190868 541447
rect 190828 541000 190880 541006
rect 190828 540942 190880 540948
rect 191470 540288 191526 540297
rect 191470 540223 191526 540232
rect 191564 540252 191616 540258
rect 191484 539646 191512 540223
rect 191564 540194 191616 540200
rect 191576 540161 191604 540194
rect 191562 540152 191618 540161
rect 191562 540087 191618 540096
rect 191472 539640 191524 539646
rect 191472 539582 191524 539588
rect 190368 530596 190420 530602
rect 190368 530538 190420 530544
rect 191668 529922 191696 548950
rect 191656 529916 191708 529922
rect 191656 529858 191708 529864
rect 189816 518220 189868 518226
rect 189816 518162 189868 518168
rect 189722 469296 189778 469305
rect 189722 469231 189778 469240
rect 189736 416090 189764 469231
rect 190276 463004 190328 463010
rect 190276 462946 190328 462952
rect 190288 442270 190316 462946
rect 191654 458824 191710 458833
rect 191654 458759 191710 458768
rect 190366 456920 190422 456929
rect 190366 456855 190422 456864
rect 190276 442264 190328 442270
rect 190276 442206 190328 442212
rect 190276 440904 190328 440910
rect 190276 440846 190328 440852
rect 189724 416084 189776 416090
rect 189724 416026 189776 416032
rect 189724 414724 189776 414730
rect 189724 414666 189776 414672
rect 189000 393286 189120 393314
rect 188436 387796 188488 387802
rect 188436 387738 188488 387744
rect 188528 387796 188580 387802
rect 188528 387738 188580 387744
rect 188448 378894 188476 387738
rect 188986 385656 189042 385665
rect 188986 385591 189042 385600
rect 189000 385422 189028 385591
rect 188988 385416 189040 385422
rect 188988 385358 189040 385364
rect 188436 378888 188488 378894
rect 188436 378830 188488 378836
rect 189000 378185 189028 385358
rect 188986 378176 189042 378185
rect 188986 378111 189042 378120
rect 189092 378026 189120 393286
rect 189736 391270 189764 414666
rect 189724 391264 189776 391270
rect 189724 391206 189776 391212
rect 190182 387424 190238 387433
rect 190182 387359 190238 387368
rect 188908 377998 189120 378026
rect 188342 375320 188398 375329
rect 188342 375255 188398 375264
rect 187608 373448 187660 373454
rect 187608 373390 187660 373396
rect 187516 334620 187568 334626
rect 187516 334562 187568 334568
rect 187054 308000 187110 308009
rect 187054 307935 187110 307944
rect 186410 305144 186466 305153
rect 186410 305079 186466 305088
rect 186320 305040 186372 305046
rect 186320 304982 186372 304988
rect 186226 302560 186282 302569
rect 186226 302495 186282 302504
rect 186332 302190 186360 304982
rect 186320 302184 186372 302190
rect 186320 302126 186372 302132
rect 186424 297401 186452 305079
rect 186964 300824 187016 300830
rect 186964 300766 187016 300772
rect 186410 297392 186466 297401
rect 186410 297327 186466 297336
rect 186228 294704 186280 294710
rect 186228 294646 186280 294652
rect 186240 294030 186268 294646
rect 186228 294024 186280 294030
rect 186228 293966 186280 293972
rect 186136 267028 186188 267034
rect 186136 266970 186188 266976
rect 186044 252544 186096 252550
rect 186044 252486 186096 252492
rect 185504 248386 185624 248414
rect 185596 234598 185624 248386
rect 186240 242457 186268 293966
rect 186320 286340 186372 286346
rect 186320 286282 186372 286288
rect 186332 259146 186360 286282
rect 186320 259140 186372 259146
rect 186320 259082 186372 259088
rect 186320 250572 186372 250578
rect 186320 250514 186372 250520
rect 186332 250481 186360 250514
rect 186318 250472 186374 250481
rect 186318 250407 186374 250416
rect 186976 247110 187004 300766
rect 187068 286385 187096 307935
rect 187516 305040 187568 305046
rect 187514 305008 187516 305017
rect 187568 305008 187570 305017
rect 187514 304943 187570 304952
rect 187620 298178 187648 373390
rect 188356 372570 188384 375255
rect 188434 373280 188490 373289
rect 188434 373215 188490 373224
rect 188344 372564 188396 372570
rect 188344 372506 188396 372512
rect 188448 362953 188476 373215
rect 188434 362944 188490 362953
rect 188434 362879 188490 362888
rect 188908 337414 188936 377998
rect 190196 376553 190224 387359
rect 190288 384441 190316 440846
rect 190274 384432 190330 384441
rect 190274 384367 190330 384376
rect 189722 376544 189778 376553
rect 189722 376479 189778 376488
rect 190182 376544 190238 376553
rect 190182 376479 190238 376488
rect 188988 348424 189040 348430
rect 188988 348366 189040 348372
rect 188896 337408 188948 337414
rect 188896 337350 188948 337356
rect 188436 318844 188488 318850
rect 188436 318786 188488 318792
rect 188344 316056 188396 316062
rect 188344 315998 188396 316004
rect 187792 314696 187844 314702
rect 187792 314638 187844 314644
rect 187700 311976 187752 311982
rect 187700 311918 187752 311924
rect 187712 309806 187740 311918
rect 187700 309800 187752 309806
rect 187700 309742 187752 309748
rect 187698 309224 187754 309233
rect 187698 309159 187754 309168
rect 187712 309126 187740 309159
rect 187700 309120 187752 309126
rect 187700 309062 187752 309068
rect 187804 307086 187832 314638
rect 188356 312594 188384 315998
rect 188448 315382 188476 318786
rect 188436 315376 188488 315382
rect 188436 315318 188488 315324
rect 188344 312588 188396 312594
rect 188344 312530 188396 312536
rect 188896 308440 188948 308446
rect 188896 308382 188948 308388
rect 187792 307080 187844 307086
rect 187792 307022 187844 307028
rect 188068 306400 188120 306406
rect 188068 306342 188120 306348
rect 188080 305697 188108 306342
rect 188066 305688 188122 305697
rect 188066 305623 188122 305632
rect 187790 305280 187846 305289
rect 187790 305215 187846 305224
rect 187700 302320 187752 302326
rect 187700 302262 187752 302268
rect 187712 300150 187740 302262
rect 187700 300144 187752 300150
rect 187700 300086 187752 300092
rect 187804 298790 187832 305215
rect 188344 299668 188396 299674
rect 188344 299610 188396 299616
rect 187792 298784 187844 298790
rect 187792 298726 187844 298732
rect 187608 298172 187660 298178
rect 187608 298114 187660 298120
rect 187620 293282 187648 298114
rect 187608 293276 187660 293282
rect 187608 293218 187660 293224
rect 187608 289196 187660 289202
rect 187608 289138 187660 289144
rect 187054 286376 187110 286385
rect 187054 286311 187110 286320
rect 187620 285938 187648 289138
rect 187608 285932 187660 285938
rect 187608 285874 187660 285880
rect 187148 259140 187200 259146
rect 187148 259082 187200 259088
rect 187160 258126 187188 259082
rect 187148 258120 187200 258126
rect 187148 258062 187200 258068
rect 187056 256760 187108 256766
rect 187056 256702 187108 256708
rect 186964 247104 187016 247110
rect 186964 247046 187016 247052
rect 186226 242448 186282 242457
rect 186226 242383 186282 242392
rect 186318 242176 186374 242185
rect 186318 242111 186374 242120
rect 186332 241602 186360 242111
rect 186320 241596 186372 241602
rect 186320 241538 186372 241544
rect 185584 234592 185636 234598
rect 185584 234534 185636 234540
rect 185596 221513 185624 234534
rect 185582 221504 185638 221513
rect 185582 221439 185638 221448
rect 185596 100706 185624 221439
rect 185676 188352 185728 188358
rect 185676 188294 185728 188300
rect 185688 117298 185716 188294
rect 186332 186998 186360 241538
rect 186976 198014 187004 247046
rect 187068 241505 187096 256702
rect 187160 249966 187188 258062
rect 187148 249960 187200 249966
rect 187148 249902 187200 249908
rect 187148 248464 187200 248470
rect 187148 248406 187200 248412
rect 187054 241496 187110 241505
rect 187054 241431 187110 241440
rect 187160 234569 187188 248406
rect 187620 247518 187648 285874
rect 187608 247512 187660 247518
rect 187608 247454 187660 247460
rect 187698 245848 187754 245857
rect 187698 245783 187754 245792
rect 187712 245546 187740 245783
rect 187700 245540 187752 245546
rect 187700 245482 187752 245488
rect 187146 234560 187202 234569
rect 187146 234495 187202 234504
rect 188356 200802 188384 299610
rect 188436 275052 188488 275058
rect 188436 274994 188488 275000
rect 188448 234025 188476 274994
rect 188908 274038 188936 308382
rect 188896 274032 188948 274038
rect 188896 273974 188948 273980
rect 188896 253020 188948 253026
rect 188896 252962 188948 252968
rect 188908 252618 188936 252962
rect 188896 252612 188948 252618
rect 188896 252554 188948 252560
rect 188908 234433 188936 252554
rect 189000 245857 189028 348366
rect 189078 270464 189134 270473
rect 189078 270399 189134 270408
rect 189092 269249 189120 270399
rect 189078 269240 189134 269249
rect 189078 269175 189134 269184
rect 189078 253872 189134 253881
rect 189078 253807 189134 253816
rect 189092 252657 189120 253807
rect 189736 253026 189764 376479
rect 189814 351248 189870 351257
rect 189814 351183 189870 351192
rect 189828 303754 189856 351183
rect 190380 333266 190408 456855
rect 191470 456104 191526 456113
rect 191470 456039 191526 456048
rect 191484 449018 191512 456039
rect 191562 449168 191618 449177
rect 191562 449103 191564 449112
rect 191616 449103 191618 449112
rect 191564 449074 191616 449080
rect 191484 448990 191604 449018
rect 191576 447846 191604 448990
rect 191564 447840 191616 447846
rect 191562 447808 191564 447817
rect 191616 447808 191618 447817
rect 191562 447743 191618 447752
rect 191012 447092 191064 447098
rect 191012 447034 191064 447040
rect 191024 446457 191052 447034
rect 191010 446448 191066 446457
rect 191010 446383 191066 446392
rect 191012 445732 191064 445738
rect 191012 445674 191064 445680
rect 191024 445097 191052 445674
rect 191010 445088 191066 445097
rect 191010 445023 191066 445032
rect 191564 442264 191616 442270
rect 191564 442206 191616 442212
rect 191576 442105 191604 442206
rect 191562 442096 191618 442105
rect 191562 442031 191618 442040
rect 191564 441584 191616 441590
rect 191564 441526 191616 441532
rect 191576 440745 191604 441526
rect 191562 440736 191618 440745
rect 191562 440671 191618 440680
rect 191668 438954 191696 458759
rect 191576 438926 191696 438954
rect 191576 434602 191604 438926
rect 191656 438864 191708 438870
rect 191656 438806 191708 438812
rect 191668 438025 191696 438806
rect 191654 438016 191710 438025
rect 191654 437951 191710 437960
rect 191654 436656 191710 436665
rect 191654 436591 191710 436600
rect 191668 436150 191696 436591
rect 191656 436144 191708 436150
rect 191656 436086 191708 436092
rect 191654 435296 191710 435305
rect 191654 435231 191710 435240
rect 191668 434790 191696 435231
rect 191656 434784 191708 434790
rect 191656 434726 191708 434732
rect 191576 434574 191696 434602
rect 191668 434042 191696 434574
rect 191656 434036 191708 434042
rect 191656 433978 191708 433984
rect 191668 433673 191696 433978
rect 191654 433664 191710 433673
rect 191654 433599 191710 433608
rect 191656 432608 191708 432614
rect 191656 432550 191708 432556
rect 191668 432313 191696 432550
rect 191654 432304 191710 432313
rect 191654 432239 191710 432248
rect 191760 431254 191788 549086
rect 191748 431248 191800 431254
rect 191748 431190 191800 431196
rect 191760 430953 191788 431190
rect 191746 430944 191802 430953
rect 191746 430879 191802 430888
rect 191012 430568 191064 430574
rect 191012 430510 191064 430516
rect 191024 429593 191052 430510
rect 191010 429584 191066 429593
rect 191010 429519 191066 429528
rect 190828 429140 190880 429146
rect 190828 429082 190880 429088
rect 190840 428233 190868 429082
rect 190826 428224 190882 428233
rect 190826 428159 190882 428168
rect 191746 426864 191802 426873
rect 191746 426799 191802 426808
rect 191760 426494 191788 426799
rect 191748 426488 191800 426494
rect 191748 426430 191800 426436
rect 191746 425504 191802 425513
rect 191746 425439 191802 425448
rect 191760 425134 191788 425439
rect 191748 425128 191800 425134
rect 191748 425070 191800 425076
rect 191012 425060 191064 425066
rect 191012 425002 191064 425008
rect 191024 423881 191052 425002
rect 191010 423872 191066 423881
rect 191010 423807 191066 423816
rect 191746 422512 191802 422521
rect 191746 422447 191802 422456
rect 191760 422346 191788 422447
rect 191748 422340 191800 422346
rect 191748 422282 191800 422288
rect 191746 417072 191802 417081
rect 191746 417007 191802 417016
rect 191760 416838 191788 417007
rect 191748 416832 191800 416838
rect 191748 416774 191800 416780
rect 191656 416764 191708 416770
rect 191656 416706 191708 416712
rect 191668 415449 191696 416706
rect 191654 415440 191710 415449
rect 191654 415375 191710 415384
rect 191194 414080 191250 414089
rect 191194 414015 191196 414024
rect 191248 414015 191250 414024
rect 191196 413986 191248 413992
rect 191102 412720 191158 412729
rect 191102 412655 191158 412664
rect 191010 407008 191066 407017
rect 191010 406943 191066 406952
rect 191024 405754 191052 406943
rect 191012 405748 191064 405754
rect 191012 405690 191064 405696
rect 191010 402928 191066 402937
rect 191010 402863 191066 402872
rect 191024 401674 191052 402863
rect 191012 401668 191064 401674
rect 191012 401610 191064 401616
rect 191010 400208 191066 400217
rect 191010 400143 191066 400152
rect 191024 398886 191052 400143
rect 191012 398880 191064 398886
rect 191012 398822 191064 398828
rect 190826 398576 190882 398585
rect 190826 398511 190882 398520
rect 190840 397594 190868 398511
rect 190828 397588 190880 397594
rect 190828 397530 190880 397536
rect 191116 387433 191144 412655
rect 191748 411936 191800 411942
rect 191748 411878 191800 411884
rect 191760 411369 191788 411878
rect 191746 411360 191802 411369
rect 191746 411295 191802 411304
rect 191748 410576 191800 410582
rect 191748 410518 191800 410524
rect 191760 410009 191788 410518
rect 191746 410000 191802 410009
rect 191746 409935 191802 409944
rect 191748 405680 191800 405686
rect 191746 405648 191748 405657
rect 191800 405648 191802 405657
rect 191746 405583 191802 405592
rect 191748 404320 191800 404326
rect 191746 404288 191748 404297
rect 191800 404288 191802 404297
rect 191746 404223 191802 404232
rect 191748 401600 191800 401606
rect 191746 401568 191748 401577
rect 191800 401568 191802 401577
rect 191746 401503 191802 401512
rect 191194 397216 191250 397225
rect 191194 397151 191250 397160
rect 191102 387424 191158 387433
rect 191102 387359 191158 387368
rect 191208 385422 191236 397151
rect 191748 396024 191800 396030
rect 191748 395966 191800 395972
rect 191760 395865 191788 395966
rect 191746 395856 191802 395865
rect 191746 395791 191802 395800
rect 191196 385416 191248 385422
rect 191196 385358 191248 385364
rect 190458 370560 190514 370569
rect 190458 370495 190514 370504
rect 190472 334801 190500 370495
rect 190552 366376 190604 366382
rect 190552 366318 190604 366324
rect 190564 338745 190592 366318
rect 191748 338768 191800 338774
rect 190550 338736 190606 338745
rect 190550 338671 190606 338680
rect 191746 338736 191748 338745
rect 191800 338736 191802 338745
rect 191746 338671 191802 338680
rect 191746 336016 191802 336025
rect 191746 335951 191802 335960
rect 190458 334792 190514 334801
rect 190458 334727 190514 334736
rect 190368 333260 190420 333266
rect 190368 333202 190420 333208
rect 191562 330440 191618 330449
rect 191562 330375 191618 330384
rect 190368 327208 190420 327214
rect 190368 327150 190420 327156
rect 189816 303748 189868 303754
rect 189816 303690 189868 303696
rect 189724 253020 189776 253026
rect 189724 252962 189776 252968
rect 189078 252648 189134 252657
rect 189078 252583 189134 252592
rect 188986 245848 189042 245857
rect 188986 245783 189042 245792
rect 189078 245712 189134 245721
rect 189078 245647 189134 245656
rect 188894 234424 188950 234433
rect 188894 234359 188950 234368
rect 188434 234016 188490 234025
rect 188434 233951 188490 233960
rect 188988 203584 189040 203590
rect 188988 203526 189040 203532
rect 188344 200796 188396 200802
rect 188344 200738 188396 200744
rect 186964 198008 187016 198014
rect 186964 197950 187016 197956
rect 187608 192500 187660 192506
rect 187608 192442 187660 192448
rect 186320 186992 186372 186998
rect 186320 186934 186372 186940
rect 187514 154592 187570 154601
rect 187514 154527 187570 154536
rect 186228 153264 186280 153270
rect 186228 153206 186280 153212
rect 186240 148374 186268 153206
rect 186228 148368 186280 148374
rect 186228 148310 186280 148316
rect 186962 146568 187018 146577
rect 186962 146503 187018 146512
rect 186320 140820 186372 140826
rect 186320 140762 186372 140768
rect 186332 133890 186360 140762
rect 186976 135969 187004 146503
rect 186962 135960 187018 135969
rect 186962 135895 187018 135904
rect 186320 133884 186372 133890
rect 186320 133826 186372 133832
rect 187528 129742 187556 154527
rect 187516 129736 187568 129742
rect 187516 129678 187568 129684
rect 187516 126268 187568 126274
rect 187516 126210 187568 126216
rect 187528 125730 187556 126210
rect 187516 125724 187568 125730
rect 187516 125666 187568 125672
rect 185676 117292 185728 117298
rect 185676 117234 185728 117240
rect 185768 116068 185820 116074
rect 185768 116010 185820 116016
rect 185780 111110 185808 116010
rect 185768 111104 185820 111110
rect 185768 111046 185820 111052
rect 187054 106720 187110 106729
rect 187054 106655 187110 106664
rect 186228 104916 186280 104922
rect 186228 104858 186280 104864
rect 185584 100700 185636 100706
rect 185584 100642 185636 100648
rect 185122 93120 185178 93129
rect 185122 93055 185178 93064
rect 185136 86902 185164 93055
rect 185124 86896 185176 86902
rect 185124 86838 185176 86844
rect 186240 78713 186268 104858
rect 186964 102196 187016 102202
rect 186964 102138 187016 102144
rect 185582 78704 185638 78713
rect 185582 78639 185638 78648
rect 186226 78704 186282 78713
rect 186226 78639 186282 78648
rect 184940 72480 184992 72486
rect 184940 72422 184992 72428
rect 185596 70378 185624 78639
rect 186976 74526 187004 102138
rect 187068 84153 187096 106655
rect 187054 84144 187110 84153
rect 187054 84079 187110 84088
rect 186964 74520 187016 74526
rect 186964 74462 187016 74468
rect 185584 70372 185636 70378
rect 185584 70314 185636 70320
rect 184294 60616 184350 60625
rect 184294 60551 184350 60560
rect 184308 54534 184336 60551
rect 184296 54528 184348 54534
rect 184296 54470 184348 54476
rect 187528 47598 187556 125666
rect 187620 107574 187648 192442
rect 188434 154864 188490 154873
rect 188434 154799 188490 154808
rect 188342 144800 188398 144809
rect 188342 144735 188398 144744
rect 188356 143857 188384 144735
rect 188448 144226 188476 154799
rect 188804 148368 188856 148374
rect 188804 148310 188856 148316
rect 188526 146432 188582 146441
rect 188526 146367 188582 146376
rect 188436 144220 188488 144226
rect 188436 144162 188488 144168
rect 188342 143848 188398 143857
rect 188342 143783 188398 143792
rect 188356 132462 188384 143783
rect 188540 139398 188568 146367
rect 188528 139392 188580 139398
rect 188528 139334 188580 139340
rect 188344 132456 188396 132462
rect 188344 132398 188396 132404
rect 188816 124846 188844 148310
rect 189000 135250 189028 203526
rect 189092 152425 189120 245647
rect 189722 242992 189778 243001
rect 189722 242927 189778 242936
rect 189736 237386 189764 242927
rect 189724 237380 189776 237386
rect 189724 237322 189776 237328
rect 189828 215937 189856 303690
rect 189998 299568 190054 299577
rect 189998 299503 190054 299512
rect 190012 296002 190040 299503
rect 190000 295996 190052 296002
rect 190000 295938 190052 295944
rect 189906 295488 189962 295497
rect 189906 295423 189962 295432
rect 189920 285666 189948 295423
rect 189908 285660 189960 285666
rect 189908 285602 189960 285608
rect 189908 281580 189960 281586
rect 189908 281522 189960 281528
rect 189920 239873 189948 281522
rect 190380 246430 190408 327150
rect 191472 302184 191524 302190
rect 191472 302126 191524 302132
rect 191484 300937 191512 302126
rect 191470 300928 191526 300937
rect 191470 300863 191526 300872
rect 191470 298752 191526 298761
rect 191470 298687 191526 298696
rect 191484 298178 191512 298687
rect 191472 298172 191524 298178
rect 191472 298114 191524 298120
rect 191470 297664 191526 297673
rect 191470 297599 191526 297608
rect 191484 296750 191512 297599
rect 191472 296744 191524 296750
rect 191472 296686 191524 296692
rect 191472 294704 191524 294710
rect 191472 294646 191524 294652
rect 191484 294409 191512 294646
rect 191470 294400 191526 294409
rect 191470 294335 191526 294344
rect 191470 293312 191526 293321
rect 191470 293247 191526 293256
rect 191484 292602 191512 293247
rect 191472 292596 191524 292602
rect 191472 292538 191524 292544
rect 191472 292460 191524 292466
rect 191472 292402 191524 292408
rect 191484 292233 191512 292402
rect 191470 292224 191526 292233
rect 191470 292159 191526 292168
rect 191470 291136 191526 291145
rect 191470 291071 191526 291080
rect 190826 290048 190882 290057
rect 190826 289983 190828 289992
rect 190880 289983 190882 289992
rect 190828 289954 190880 289960
rect 191484 289950 191512 291071
rect 191472 289944 191524 289950
rect 191472 289886 191524 289892
rect 191472 289128 191524 289134
rect 191472 289070 191524 289076
rect 191484 288969 191512 289070
rect 191470 288960 191526 288969
rect 191470 288895 191526 288904
rect 191470 287872 191526 287881
rect 191470 287807 191526 287816
rect 191484 287774 191512 287807
rect 191472 287768 191524 287774
rect 191472 287710 191524 287716
rect 191378 286784 191434 286793
rect 191378 286719 191434 286728
rect 191392 285938 191420 286719
rect 191472 286340 191524 286346
rect 191472 286282 191524 286288
rect 191380 285932 191432 285938
rect 191380 285874 191432 285880
rect 191484 285705 191512 286282
rect 191470 285696 191526 285705
rect 191470 285631 191526 285640
rect 191470 284608 191526 284617
rect 191470 284543 191526 284552
rect 191484 284374 191512 284543
rect 191472 284368 191524 284374
rect 191472 284310 191524 284316
rect 191470 282432 191526 282441
rect 191470 282367 191526 282376
rect 191484 281654 191512 282367
rect 191472 281648 191524 281654
rect 191472 281590 191524 281596
rect 191470 281344 191526 281353
rect 191470 281279 191526 281288
rect 191484 280838 191512 281279
rect 191472 280832 191524 280838
rect 191472 280774 191524 280780
rect 191472 280288 191524 280294
rect 191470 280256 191472 280265
rect 191524 280256 191526 280265
rect 191470 280191 191526 280200
rect 191472 279472 191524 279478
rect 191472 279414 191524 279420
rect 191484 279177 191512 279414
rect 191470 279168 191526 279177
rect 191470 279103 191526 279112
rect 191470 278080 191526 278089
rect 191470 278015 191526 278024
rect 191484 277438 191512 278015
rect 191472 277432 191524 277438
rect 191472 277374 191524 277380
rect 190642 276992 190698 277001
rect 190642 276927 190698 276936
rect 190656 276078 190684 276927
rect 190644 276072 190696 276078
rect 190644 276014 190696 276020
rect 191576 275913 191604 330375
rect 191654 322144 191710 322153
rect 191654 322079 191710 322088
rect 191562 275904 191618 275913
rect 191562 275839 191618 275848
rect 191576 275058 191604 275839
rect 191564 275052 191616 275058
rect 191564 274994 191616 275000
rect 190828 274032 190880 274038
rect 190828 273974 190880 273980
rect 190840 273737 190868 273974
rect 190826 273728 190882 273737
rect 190826 273663 190882 273672
rect 191564 273216 191616 273222
rect 191564 273158 191616 273164
rect 191576 272649 191604 273158
rect 191562 272640 191618 272649
rect 191562 272575 191618 272584
rect 191562 271552 191618 271561
rect 191562 271487 191618 271496
rect 191576 270570 191604 271487
rect 191564 270564 191616 270570
rect 191564 270506 191616 270512
rect 191470 270464 191526 270473
rect 191470 270399 191526 270408
rect 191484 269249 191512 270399
rect 191564 269408 191616 269414
rect 191562 269376 191564 269385
rect 191616 269376 191618 269385
rect 191562 269311 191618 269320
rect 191470 269240 191526 269249
rect 191470 269175 191526 269184
rect 191564 269068 191616 269074
rect 191564 269010 191616 269016
rect 191576 268297 191604 269010
rect 191562 268288 191618 268297
rect 191562 268223 191618 268232
rect 191668 267734 191696 322079
rect 191576 267706 191696 267734
rect 190644 265668 190696 265674
rect 190644 265610 190696 265616
rect 190656 265033 190684 265610
rect 190642 265024 190698 265033
rect 190642 264959 190698 264968
rect 191378 260672 191434 260681
rect 191378 260607 191434 260616
rect 191392 260234 191420 260607
rect 191380 260228 191432 260234
rect 191380 260170 191432 260176
rect 190460 258188 190512 258194
rect 190460 258130 190512 258136
rect 190472 258097 190500 258130
rect 190458 258088 190514 258097
rect 190458 258023 190514 258032
rect 190642 257408 190698 257417
rect 190642 257343 190698 257352
rect 190656 257242 190684 257343
rect 190644 257236 190696 257242
rect 190644 257178 190696 257184
rect 191012 255264 191064 255270
rect 191010 255232 191012 255241
rect 191064 255232 191066 255241
rect 191010 255167 191066 255176
rect 191104 252544 191156 252550
rect 191104 252486 191156 252492
rect 191010 251968 191066 251977
rect 191010 251903 191012 251912
rect 191064 251903 191066 251912
rect 191012 251874 191064 251880
rect 191010 249792 191066 249801
rect 191010 249727 191066 249736
rect 191024 248470 191052 249727
rect 191012 248464 191064 248470
rect 191012 248406 191064 248412
rect 190460 247512 190512 247518
rect 190460 247454 190512 247460
rect 190368 246424 190420 246430
rect 190368 246366 190420 246372
rect 189906 239864 189962 239873
rect 189906 239799 189962 239808
rect 189814 215928 189870 215937
rect 189814 215863 189870 215872
rect 190472 184210 190500 247454
rect 191116 204270 191144 252486
rect 191576 248577 191604 267706
rect 191656 266348 191708 266354
rect 191656 266290 191708 266296
rect 191668 266121 191696 266290
rect 191654 266112 191710 266121
rect 191654 266047 191710 266056
rect 191654 262848 191710 262857
rect 191654 262783 191710 262792
rect 191668 262274 191696 262783
rect 191656 262268 191708 262274
rect 191656 262210 191708 262216
rect 191654 261760 191710 261769
rect 191654 261695 191710 261704
rect 191668 260914 191696 261695
rect 191656 260908 191708 260914
rect 191656 260850 191708 260856
rect 191654 259584 191710 259593
rect 191654 259519 191710 259528
rect 191668 259486 191696 259519
rect 191656 259480 191708 259486
rect 191656 259422 191708 259428
rect 191654 256320 191710 256329
rect 191654 256255 191710 256264
rect 191668 256018 191696 256255
rect 191656 256012 191708 256018
rect 191656 255954 191708 255960
rect 191654 250880 191710 250889
rect 191654 250815 191710 250824
rect 191668 250578 191696 250815
rect 191656 250572 191708 250578
rect 191656 250514 191708 250520
rect 191562 248568 191618 248577
rect 191562 248503 191618 248512
rect 191760 248414 191788 335951
rect 191852 267734 191880 567310
rect 193126 553140 193182 553149
rect 193126 553075 193182 553084
rect 193140 529310 193168 553075
rect 253112 539368 253164 539374
rect 253112 539310 253164 539316
rect 193600 536110 193628 539172
rect 193588 536104 193640 536110
rect 193588 536046 193640 536052
rect 194152 535537 194180 539172
rect 194138 535528 194194 535537
rect 194138 535463 194194 535472
rect 194704 532001 194732 539172
rect 195440 536081 195468 539172
rect 195992 536246 196020 539172
rect 196084 539158 196742 539186
rect 196912 539158 197294 539186
rect 197464 539158 198030 539186
rect 198200 539158 198582 539186
rect 198752 539158 199318 539186
rect 199396 539158 199870 539186
rect 195980 536240 196032 536246
rect 195980 536182 196032 536188
rect 195426 536072 195482 536081
rect 195426 536007 195482 536016
rect 195980 533452 196032 533458
rect 195980 533394 196032 533400
rect 194690 531992 194746 532001
rect 194690 531927 194746 531936
rect 193128 529304 193180 529310
rect 193128 529246 193180 529252
rect 195244 518220 195296 518226
rect 195244 518162 195296 518168
rect 193496 514140 193548 514146
rect 193496 514082 193548 514088
rect 191932 510944 191984 510950
rect 191932 510886 191984 510892
rect 191944 465730 191972 510886
rect 191932 465724 191984 465730
rect 191932 465666 191984 465672
rect 193036 465724 193088 465730
rect 193036 465666 193088 465672
rect 192666 450392 192722 450401
rect 192666 450327 192722 450336
rect 192680 447409 192708 450327
rect 192760 449812 192812 449818
rect 192760 449754 192812 449760
rect 192772 448633 192800 449754
rect 192758 448624 192814 448633
rect 192758 448559 192814 448568
rect 192666 447400 192722 447409
rect 192666 447335 192722 447344
rect 193048 443737 193076 465666
rect 193126 461680 193182 461689
rect 193126 461615 193182 461624
rect 193034 443728 193090 443737
rect 193034 443663 193090 443672
rect 193048 443086 193076 443663
rect 193036 443080 193088 443086
rect 193036 443022 193088 443028
rect 192484 420232 192536 420238
rect 192484 420174 192536 420180
rect 192390 419792 192446 419801
rect 192390 419727 192446 419736
rect 192404 419558 192432 419727
rect 192392 419552 192444 419558
rect 192392 419494 192444 419500
rect 192496 408649 192524 420174
rect 193140 419801 193168 461615
rect 193402 454880 193458 454889
rect 193402 454815 193458 454824
rect 193310 452568 193366 452577
rect 193310 452503 193366 452512
rect 193220 450288 193272 450294
rect 193220 450230 193272 450236
rect 193232 449449 193260 450230
rect 193218 449440 193274 449449
rect 193218 449375 193274 449384
rect 193324 440910 193352 452503
rect 193416 449970 193444 454815
rect 193508 450294 193536 514082
rect 195256 498846 195284 518162
rect 195992 504490 196020 533394
rect 196084 526454 196112 539158
rect 196912 533458 196940 539158
rect 197464 538214 197492 539158
rect 197372 538186 197492 538214
rect 197372 535430 197400 538186
rect 197636 536240 197688 536246
rect 197636 536182 197688 536188
rect 197450 535528 197506 535537
rect 197450 535463 197506 535472
rect 197360 535424 197412 535430
rect 197360 535366 197412 535372
rect 196900 533452 196952 533458
rect 196900 533394 196952 533400
rect 197360 533452 197412 533458
rect 197360 533394 197412 533400
rect 196072 526448 196124 526454
rect 196072 526390 196124 526396
rect 196624 523728 196676 523734
rect 196624 523670 196676 523676
rect 195980 504484 196032 504490
rect 195980 504426 196032 504432
rect 195244 498840 195296 498846
rect 195244 498782 195296 498788
rect 195426 498808 195482 498817
rect 195426 498743 195482 498752
rect 195334 491872 195390 491881
rect 195334 491807 195390 491816
rect 195242 478136 195298 478145
rect 195242 478071 195298 478080
rect 194508 453348 194560 453354
rect 194508 453290 194560 453296
rect 193496 450288 193548 450294
rect 193496 450230 193548 450236
rect 193416 449942 193614 449970
rect 194520 449750 194548 453290
rect 195256 452742 195284 478071
rect 195348 476785 195376 491807
rect 195440 483682 195468 498743
rect 195428 483676 195480 483682
rect 195428 483618 195480 483624
rect 195334 476776 195390 476785
rect 195334 476711 195390 476720
rect 196636 468625 196664 523670
rect 197372 491978 197400 533394
rect 197464 528554 197492 535463
rect 197648 528562 197676 536182
rect 198200 533458 198228 539158
rect 198188 533452 198240 533458
rect 198188 533394 198240 533400
rect 198752 529145 198780 539158
rect 199396 536625 199424 539158
rect 199382 536616 199438 536625
rect 199382 536551 199438 536560
rect 199396 535401 199424 536551
rect 199382 535392 199438 535401
rect 199382 535327 199438 535336
rect 198832 529916 198884 529922
rect 198832 529858 198884 529864
rect 198738 529136 198794 529145
rect 198738 529071 198794 529080
rect 197636 528556 197688 528562
rect 197464 528526 197584 528554
rect 197452 523796 197504 523802
rect 197452 523738 197504 523744
rect 197360 491972 197412 491978
rect 197360 491914 197412 491920
rect 196622 468616 196678 468625
rect 195336 468580 195388 468586
rect 196622 468551 196678 468560
rect 195336 468522 195388 468528
rect 195244 452736 195296 452742
rect 195244 452678 195296 452684
rect 195256 451274 195284 452678
rect 195072 451246 195284 451274
rect 195072 450242 195100 451246
rect 194718 450214 195100 450242
rect 195348 449818 195376 468522
rect 197360 467152 197412 467158
rect 197360 467094 197412 467100
rect 197372 464370 197400 467094
rect 197360 464364 197412 464370
rect 197360 464306 197412 464312
rect 197360 458312 197412 458318
rect 197360 458254 197412 458260
rect 196072 456068 196124 456074
rect 196072 456010 196124 456016
rect 195612 451376 195664 451382
rect 195612 451318 195664 451324
rect 195624 450228 195652 451318
rect 196084 450242 196112 456010
rect 197372 450242 197400 458254
rect 197464 452577 197492 523738
rect 197450 452568 197506 452577
rect 197450 452503 197506 452512
rect 197556 450401 197584 528526
rect 197636 528498 197688 528504
rect 198002 490648 198058 490657
rect 198002 490583 198058 490592
rect 198016 458318 198044 490583
rect 198740 478916 198792 478922
rect 198740 478858 198792 478864
rect 198752 478242 198780 478858
rect 198740 478236 198792 478242
rect 198740 478178 198792 478184
rect 198740 476604 198792 476610
rect 198740 476546 198792 476552
rect 198004 458312 198056 458318
rect 198004 458254 198056 458260
rect 197910 454064 197966 454073
rect 197910 453999 197966 454008
rect 197542 450392 197598 450401
rect 197542 450327 197598 450336
rect 197924 450242 197952 453999
rect 198752 451274 198780 476546
rect 198844 453966 198872 529858
rect 199396 478922 199424 535327
rect 200408 533458 200436 539172
rect 200776 539158 201158 539186
rect 201604 539158 201710 539186
rect 202064 539158 202446 539186
rect 200776 538214 200804 539158
rect 200500 538186 200804 538214
rect 200396 533452 200448 533458
rect 200396 533394 200448 533400
rect 200500 533338 200528 538186
rect 200132 533310 200528 533338
rect 201500 533384 201552 533390
rect 201500 533326 201552 533332
rect 200132 519654 200160 533310
rect 200212 530596 200264 530602
rect 200212 530538 200264 530544
rect 200120 519648 200172 519654
rect 200120 519590 200172 519596
rect 199476 485104 199528 485110
rect 199476 485046 199528 485052
rect 199488 478990 199516 485046
rect 199476 478984 199528 478990
rect 199476 478926 199528 478932
rect 199384 478916 199436 478922
rect 199384 478858 199436 478864
rect 199488 476610 199516 478926
rect 199476 476604 199528 476610
rect 199476 476546 199528 476552
rect 200224 456249 200252 530538
rect 201512 465050 201540 533326
rect 201604 527882 201632 539158
rect 202064 533390 202092 539158
rect 202984 538121 203012 539172
rect 203260 539158 203734 539186
rect 204286 539158 204484 539186
rect 202970 538112 203026 538121
rect 202970 538047 203026 538056
rect 202984 536897 203012 538047
rect 202970 536888 203026 536897
rect 202970 536823 203026 536832
rect 202052 533384 202104 533390
rect 202052 533326 202104 533332
rect 203260 528554 203288 539158
rect 203522 536888 203578 536897
rect 203522 536823 203578 536832
rect 202892 528526 203288 528554
rect 201592 527876 201644 527882
rect 201592 527818 201644 527824
rect 202892 514146 202920 528526
rect 203536 521014 203564 536823
rect 204456 530641 204484 539158
rect 204548 539158 205022 539186
rect 205192 539158 205574 539186
rect 205652 539158 206310 539186
rect 204442 530632 204498 530641
rect 204442 530567 204498 530576
rect 204548 529242 204576 539158
rect 205192 538214 205220 539158
rect 204640 538186 205220 538214
rect 204536 529236 204588 529242
rect 204536 529178 204588 529184
rect 204640 528554 204668 538186
rect 205086 530632 205142 530641
rect 205086 530567 205142 530576
rect 204272 528526 204668 528554
rect 203524 521008 203576 521014
rect 203524 520950 203576 520956
rect 204272 520946 204300 528526
rect 204260 520940 204312 520946
rect 204260 520882 204312 520888
rect 204904 515500 204956 515506
rect 204904 515442 204956 515448
rect 202880 514140 202932 514146
rect 202880 514082 202932 514088
rect 203522 512680 203578 512689
rect 203522 512615 203578 512624
rect 202142 509824 202198 509833
rect 202142 509759 202198 509768
rect 201500 465044 201552 465050
rect 201500 464986 201552 464992
rect 201498 462360 201554 462369
rect 201498 462295 201554 462304
rect 201512 460934 201540 462295
rect 201512 460906 201816 460934
rect 201406 458960 201462 458969
rect 201406 458895 201462 458904
rect 200210 456240 200266 456249
rect 200210 456175 200266 456184
rect 198832 453960 198884 453966
rect 198832 453902 198884 453908
rect 200396 453960 200448 453966
rect 200396 453902 200448 453908
rect 198844 453257 198872 453902
rect 198830 453248 198886 453257
rect 198830 453183 198886 453192
rect 198752 451246 198872 451274
rect 198844 450242 198872 451246
rect 196084 450214 196558 450242
rect 197372 450214 197478 450242
rect 197924 450214 198398 450242
rect 198844 450214 199318 450242
rect 200408 450228 200436 453902
rect 201420 452713 201448 458895
rect 200854 452704 200910 452713
rect 200854 452639 200910 452648
rect 201406 452704 201462 452713
rect 201406 452639 201462 452648
rect 200868 450242 200896 452639
rect 201788 450242 201816 460906
rect 202156 454753 202184 509759
rect 203536 489190 203564 512615
rect 203614 489288 203670 489297
rect 203614 489223 203670 489232
rect 203524 489184 203576 489190
rect 203524 489126 203576 489132
rect 202878 483712 202934 483721
rect 202878 483647 202934 483656
rect 202786 465896 202842 465905
rect 202786 465831 202842 465840
rect 202800 462369 202828 465831
rect 202786 462360 202842 462369
rect 202786 462295 202842 462304
rect 202142 454744 202198 454753
rect 202142 454679 202198 454688
rect 202892 450537 202920 483647
rect 203628 467265 203656 489223
rect 203614 467256 203670 467265
rect 203614 467191 203670 467200
rect 204260 466540 204312 466546
rect 204260 466482 204312 466488
rect 204272 463690 204300 466482
rect 204260 463684 204312 463690
rect 204260 463626 204312 463632
rect 204272 460934 204300 463626
rect 204916 461553 204944 515442
rect 204996 509992 205048 509998
rect 204996 509934 205048 509940
rect 205008 463010 205036 509934
rect 205100 509930 205128 530567
rect 205652 527950 205680 539158
rect 206376 535288 206428 535294
rect 206376 535230 206428 535236
rect 206284 533384 206336 533390
rect 206284 533326 206336 533332
rect 205640 527944 205692 527950
rect 205640 527886 205692 527892
rect 205640 511284 205692 511290
rect 205640 511226 205692 511232
rect 205088 509924 205140 509930
rect 205088 509866 205140 509872
rect 204996 463004 205048 463010
rect 204996 462946 205048 462952
rect 204902 461544 204958 461553
rect 204902 461479 204958 461488
rect 204272 460906 204576 460934
rect 202970 457600 203026 457609
rect 202970 457535 203026 457544
rect 202984 454073 203012 457535
rect 202970 454064 203026 454073
rect 202970 453999 203026 454008
rect 202878 450528 202934 450537
rect 202878 450463 202934 450472
rect 202984 450242 203012 453999
rect 204168 452668 204220 452674
rect 204168 452610 204220 452616
rect 204180 450566 204208 452610
rect 204168 450560 204220 450566
rect 204074 450528 204130 450537
rect 204168 450502 204220 450508
rect 204074 450463 204130 450472
rect 200868 450214 201342 450242
rect 201788 450214 202262 450242
rect 202984 450214 203182 450242
rect 204088 449970 204116 450463
rect 204548 450242 204576 460906
rect 204548 450214 205022 450242
rect 205652 450129 205680 511226
rect 206296 469878 206324 533326
rect 206388 518226 206416 535230
rect 206848 532642 206876 539172
rect 207400 538257 207428 539172
rect 207386 538248 207442 538257
rect 207386 538183 207442 538192
rect 208136 535537 208164 539172
rect 208412 539158 208702 539186
rect 208122 535528 208178 535537
rect 208122 535463 208178 535472
rect 206836 532636 206888 532642
rect 206836 532578 206888 532584
rect 207204 529304 207256 529310
rect 207204 529246 207256 529252
rect 206376 518220 206428 518226
rect 206376 518162 206428 518168
rect 206376 507204 206428 507210
rect 206376 507146 206428 507152
rect 206388 471209 206416 507146
rect 206468 475380 206520 475386
rect 206468 475322 206520 475328
rect 206374 471200 206430 471209
rect 206374 471135 206430 471144
rect 206284 469872 206336 469878
rect 206284 469814 206336 469820
rect 206480 457473 206508 475322
rect 207112 465044 207164 465050
rect 207112 464986 207164 464992
rect 206466 457464 206522 457473
rect 206466 457399 206522 457408
rect 207124 454170 207152 464986
rect 207216 460934 207244 529246
rect 208412 512650 208440 539158
rect 209424 534070 209452 539172
rect 209976 535294 210004 539172
rect 210160 539158 210726 539186
rect 209964 535288 210016 535294
rect 209964 535230 210016 535236
rect 209412 534064 209464 534070
rect 209412 534006 209464 534012
rect 209044 532976 209096 532982
rect 209044 532918 209096 532924
rect 208400 512644 208452 512650
rect 208400 512586 208452 512592
rect 209056 489161 209084 532918
rect 210160 528554 210188 539158
rect 211264 532982 211292 539172
rect 212000 538214 212028 539172
rect 212000 538186 212488 538214
rect 212460 536489 212488 538186
rect 212446 536480 212502 536489
rect 212446 536415 212502 536424
rect 211804 533452 211856 533458
rect 211804 533394 211856 533400
rect 211252 532976 211304 532982
rect 211252 532918 211304 532924
rect 209792 528526 210188 528554
rect 209042 489152 209098 489161
rect 209042 489087 209098 489096
rect 209042 483032 209098 483041
rect 209042 482967 209098 482976
rect 209056 471209 209084 482967
rect 209792 472666 209820 528526
rect 210424 500336 210476 500342
rect 210424 500278 210476 500284
rect 210238 492824 210294 492833
rect 210238 492759 210294 492768
rect 210252 492726 210280 492759
rect 210240 492720 210292 492726
rect 210240 492662 210292 492668
rect 209780 472660 209832 472666
rect 209780 472602 209832 472608
rect 209792 472546 209820 472602
rect 209792 472518 209912 472546
rect 209042 471200 209098 471209
rect 209042 471135 209098 471144
rect 209778 470656 209834 470665
rect 209778 470591 209834 470600
rect 209792 460934 209820 470591
rect 209884 464681 209912 472518
rect 209870 464672 209926 464681
rect 209870 464607 209926 464616
rect 207216 460906 207336 460934
rect 209792 460906 210372 460934
rect 207112 454164 207164 454170
rect 207112 454106 207164 454112
rect 207124 450242 207152 454106
rect 207308 450265 207336 460906
rect 208398 460320 208454 460329
rect 208398 460255 208454 460264
rect 207046 450214 207152 450242
rect 207294 450256 207350 450265
rect 207294 450191 207350 450200
rect 207570 450256 207626 450265
rect 208412 450242 208440 460255
rect 209872 454096 209924 454102
rect 209872 454038 209924 454044
rect 209884 450242 209912 454038
rect 207626 450214 207966 450242
rect 208412 450214 208886 450242
rect 209806 450214 209912 450242
rect 210344 450242 210372 460906
rect 210436 454102 210464 500278
rect 210516 492720 210568 492726
rect 210516 492662 210568 492668
rect 210528 486538 210556 492662
rect 210516 486532 210568 486538
rect 210516 486474 210568 486480
rect 211816 459542 211844 533394
rect 212460 509250 212488 536415
rect 212552 533458 212580 539172
rect 212644 539158 213118 539186
rect 213196 539158 213854 539186
rect 214024 539158 214406 539186
rect 214760 539158 215142 539186
rect 215404 539158 215694 539186
rect 212540 533452 212592 533458
rect 212540 533394 212592 533400
rect 212644 533361 212672 539158
rect 213196 538214 213224 539158
rect 212736 538186 213224 538214
rect 212630 533352 212686 533361
rect 212630 533287 212686 533296
rect 212448 509244 212500 509250
rect 212448 509186 212500 509192
rect 212460 508570 212488 509186
rect 212448 508564 212500 508570
rect 212448 508506 212500 508512
rect 212736 465730 212764 538186
rect 213184 533452 213236 533458
rect 213184 533394 213236 533400
rect 213196 515438 213224 533394
rect 213274 533352 213330 533361
rect 213274 533287 213330 533296
rect 213288 523705 213316 533287
rect 213920 529780 213972 529786
rect 213920 529722 213972 529728
rect 213274 523696 213330 523705
rect 213274 523631 213330 523640
rect 213184 515432 213236 515438
rect 213184 515374 213236 515380
rect 213184 511284 213236 511290
rect 213184 511226 213236 511232
rect 213196 468586 213224 511226
rect 213932 479534 213960 529722
rect 214024 494834 214052 539158
rect 214656 535560 214708 535566
rect 214656 535502 214708 535508
rect 214564 529984 214616 529990
rect 214564 529926 214616 529932
rect 214012 494828 214064 494834
rect 214012 494770 214064 494776
rect 213920 479528 213972 479534
rect 213920 479470 213972 479476
rect 213184 468580 213236 468586
rect 213184 468522 213236 468528
rect 212724 465724 212776 465730
rect 212724 465666 212776 465672
rect 214576 464545 214604 529926
rect 214668 522986 214696 535502
rect 214760 529786 214788 539158
rect 215404 536761 215432 539158
rect 215390 536752 215446 536761
rect 215390 536687 215446 536696
rect 214748 529780 214800 529786
rect 214748 529722 214800 529728
rect 214656 522980 214708 522986
rect 214656 522922 214708 522928
rect 214656 496188 214708 496194
rect 214656 496130 214708 496136
rect 214562 464536 214618 464545
rect 214562 464471 214618 464480
rect 213918 464400 213974 464409
rect 213918 464335 213974 464344
rect 213932 463729 213960 464335
rect 213918 463720 213974 463729
rect 213918 463655 213974 463664
rect 213828 461644 213880 461650
rect 213828 461586 213880 461592
rect 211804 459536 211856 459542
rect 211804 459478 211856 459484
rect 213840 456822 213868 461586
rect 213932 460934 213960 463655
rect 213932 460906 214144 460934
rect 213276 456816 213328 456822
rect 213276 456758 213328 456764
rect 213828 456816 213880 456822
rect 213828 456758 213880 456764
rect 211160 455456 211212 455462
rect 211160 455398 211212 455404
rect 210424 454096 210476 454102
rect 210424 454038 210476 454044
rect 211172 450242 211200 455398
rect 212630 454744 212686 454753
rect 212630 454679 212686 454688
rect 212644 450242 212672 454679
rect 213288 450242 213316 456758
rect 214116 450242 214144 460906
rect 214668 455394 214696 496130
rect 215300 478916 215352 478922
rect 215300 478858 215352 478864
rect 215312 460934 215340 478858
rect 215404 461689 215432 536687
rect 216416 535566 216444 539172
rect 216404 535560 216456 535566
rect 216404 535502 216456 535508
rect 216968 535498 216996 539172
rect 217244 539158 217718 539186
rect 218072 539158 218270 539186
rect 215944 535492 215996 535498
rect 215944 535434 215996 535440
rect 216956 535492 217008 535498
rect 216956 535434 217008 535440
rect 215956 518294 215984 535434
rect 217244 528554 217272 539158
rect 217324 534880 217376 534886
rect 217324 534822 217376 534828
rect 216784 528526 217272 528554
rect 215944 518288 215996 518294
rect 215944 518230 215996 518236
rect 216784 498914 216812 528526
rect 217336 500274 217364 534822
rect 217324 500268 217376 500274
rect 217324 500210 217376 500216
rect 216772 498908 216824 498914
rect 216772 498850 216824 498856
rect 217324 496188 217376 496194
rect 217324 496130 217376 496136
rect 217336 482322 217364 496130
rect 217324 482316 217376 482322
rect 217324 482258 217376 482264
rect 218072 479534 218100 539158
rect 218992 533361 219020 539172
rect 218978 533352 219034 533361
rect 218978 533287 219034 533296
rect 219544 530641 219572 539172
rect 219636 539158 220110 539186
rect 220846 539158 220952 539186
rect 219530 530632 219586 530641
rect 219530 530567 219586 530576
rect 219636 529990 219664 539158
rect 220082 533352 220138 533361
rect 220082 533287 220138 533296
rect 219624 529984 219676 529990
rect 219624 529926 219676 529932
rect 219440 526448 219492 526454
rect 219440 526390 219492 526396
rect 218704 525088 218756 525094
rect 218704 525030 218756 525036
rect 218152 486464 218204 486470
rect 218152 486406 218204 486412
rect 218060 479528 218112 479534
rect 218060 479470 218112 479476
rect 217324 472660 217376 472666
rect 217324 472602 217376 472608
rect 216680 465112 216732 465118
rect 216680 465054 216732 465060
rect 216692 461718 216720 465054
rect 216680 461712 216732 461718
rect 215390 461680 215446 461689
rect 216680 461654 216732 461660
rect 215390 461615 215446 461624
rect 217336 461582 217364 472602
rect 216680 461576 216732 461582
rect 216680 461518 216732 461524
rect 217324 461576 217376 461582
rect 217324 461518 217376 461524
rect 216692 461038 216720 461518
rect 216680 461032 216732 461038
rect 216680 460974 216732 460980
rect 216692 460934 216720 460974
rect 215312 460906 216076 460934
rect 216692 460906 216904 460934
rect 215390 460320 215446 460329
rect 215390 460255 215446 460264
rect 215404 455569 215432 460255
rect 215390 455560 215446 455569
rect 215390 455495 215446 455504
rect 214656 455388 214708 455394
rect 214656 455330 214708 455336
rect 215404 450242 215432 455495
rect 216048 450242 216076 460906
rect 216876 450242 216904 460906
rect 218164 456142 218192 486406
rect 218716 485081 218744 525030
rect 218702 485072 218758 485081
rect 218702 485007 218758 485016
rect 218702 482216 218758 482225
rect 218702 482151 218758 482160
rect 218152 456136 218204 456142
rect 218152 456078 218204 456084
rect 218716 452674 218744 482151
rect 219452 456929 219480 526390
rect 220096 487898 220124 533287
rect 220924 494834 220952 539158
rect 221384 538354 221412 539172
rect 221372 538348 221424 538354
rect 221372 538290 221424 538296
rect 222120 537538 222148 539172
rect 222108 537532 222160 537538
rect 222108 537474 222160 537480
rect 222672 533458 222700 539172
rect 222764 539158 223422 539186
rect 222660 533452 222712 533458
rect 222660 533394 222712 533400
rect 222764 528554 222792 539158
rect 223578 538248 223634 538257
rect 223578 538183 223634 538192
rect 222842 535528 222898 535537
rect 222842 535463 222898 535472
rect 222212 528526 222792 528554
rect 222212 523734 222240 528526
rect 222200 523728 222252 523734
rect 222200 523670 222252 523676
rect 222200 508564 222252 508570
rect 222200 508506 222252 508512
rect 220912 494828 220964 494834
rect 220912 494770 220964 494776
rect 222108 489184 222160 489190
rect 222108 489126 222160 489132
rect 220084 487892 220136 487898
rect 220084 487834 220136 487840
rect 219438 456920 219494 456929
rect 219438 456855 219494 456864
rect 219806 456920 219862 456929
rect 219806 456855 219862 456864
rect 218980 456136 219032 456142
rect 218980 456078 219032 456084
rect 218704 452668 218756 452674
rect 218704 452610 218756 452616
rect 218716 450242 218744 452610
rect 210344 450214 210726 450242
rect 211172 450214 211646 450242
rect 212644 450214 212750 450242
rect 213288 450214 213670 450242
rect 214116 450214 214590 450242
rect 215404 450214 215510 450242
rect 216048 450214 216430 450242
rect 216876 450214 217350 450242
rect 218454 450214 218744 450242
rect 218992 450242 219020 456078
rect 219820 450242 219848 456855
rect 222120 455326 222148 489126
rect 221648 455320 221700 455326
rect 221648 455262 221700 455268
rect 222108 455320 222160 455326
rect 222108 455262 222160 455268
rect 221660 454102 221688 455262
rect 222212 454753 222240 508506
rect 222856 475386 222884 535463
rect 222934 534032 222990 534041
rect 222934 533967 222990 533976
rect 222948 494766 222976 533967
rect 223592 531282 223620 538183
rect 223960 533361 223988 539172
rect 224696 538257 224724 539172
rect 224682 538248 224738 538257
rect 224682 538183 224738 538192
rect 225248 536110 225276 539172
rect 225524 539158 225998 539186
rect 225236 536104 225288 536110
rect 225236 536046 225288 536052
rect 223946 533352 224002 533361
rect 223946 533287 224002 533296
rect 223580 531276 223632 531282
rect 223580 531218 223632 531224
rect 222936 494760 222988 494766
rect 222936 494702 222988 494708
rect 223592 484430 223620 531218
rect 225524 528554 225552 539158
rect 226536 535537 226564 539172
rect 226720 539158 227102 539186
rect 226522 535528 226578 535537
rect 226522 535463 226578 535472
rect 226720 528554 226748 539158
rect 226984 536104 227036 536110
rect 226984 536046 227036 536052
rect 224972 528526 225552 528554
rect 226352 528526 226748 528554
rect 223580 484424 223632 484430
rect 223580 484366 223632 484372
rect 223592 480254 223620 484366
rect 223592 480226 223712 480254
rect 222844 475380 222896 475386
rect 222844 475322 222896 475328
rect 223580 468580 223632 468586
rect 223580 468522 223632 468528
rect 223486 456920 223542 456929
rect 223486 456855 223542 456864
rect 222198 454744 222254 454753
rect 222198 454679 222254 454688
rect 221648 454096 221700 454102
rect 221648 454038 221700 454044
rect 222106 454064 222162 454073
rect 221188 454028 221240 454034
rect 221188 453970 221240 453976
rect 218992 450214 219374 450242
rect 219820 450214 220294 450242
rect 221200 450228 221228 453970
rect 221660 450242 221688 454038
rect 223500 454034 223528 456855
rect 222106 453999 222162 454008
rect 223488 454028 223540 454034
rect 222120 453257 222148 453999
rect 223488 453970 223540 453976
rect 222106 453248 222162 453257
rect 222106 453183 222162 453192
rect 223028 452668 223080 452674
rect 223028 452610 223080 452616
rect 221660 450214 222134 450242
rect 223040 450228 223068 452610
rect 223592 451274 223620 468522
rect 223684 457473 223712 480226
rect 224972 476814 225000 528526
rect 226248 526312 226300 526318
rect 226248 526254 226300 526260
rect 224960 476808 225012 476814
rect 224960 476750 225012 476756
rect 226260 466478 226288 526254
rect 226352 474842 226380 528526
rect 226996 522986 227024 536046
rect 227824 533458 227852 539172
rect 227916 539158 228390 539186
rect 229126 539158 229324 539186
rect 227812 533452 227864 533458
rect 227812 533394 227864 533400
rect 227916 528554 227944 539158
rect 228364 530596 228416 530602
rect 228364 530538 228416 530544
rect 227732 528526 227944 528554
rect 226984 522980 227036 522986
rect 226984 522922 227036 522928
rect 227628 491972 227680 491978
rect 227628 491914 227680 491920
rect 226340 474836 226392 474842
rect 226340 474778 226392 474784
rect 226984 474836 227036 474842
rect 226984 474778 227036 474784
rect 224960 466472 225012 466478
rect 224960 466414 225012 466420
rect 226248 466472 226300 466478
rect 226248 466414 226300 466420
rect 224972 460934 225000 466414
rect 226340 463820 226392 463826
rect 226340 463762 226392 463768
rect 226352 460934 226380 463762
rect 224972 460906 225644 460934
rect 226352 460906 226472 460934
rect 223670 457464 223726 457473
rect 223670 457399 223726 457408
rect 223684 456929 223712 457399
rect 223670 456920 223726 456929
rect 223670 456855 223726 456864
rect 225052 455796 225104 455802
rect 225052 455738 225104 455744
rect 223592 451246 223712 451274
rect 223684 450242 223712 451246
rect 223684 450214 224158 450242
rect 225064 450228 225092 455738
rect 225616 450242 225644 460906
rect 226444 450242 226472 460906
rect 226996 455802 227024 474778
rect 227640 463826 227668 491914
rect 227732 490521 227760 528526
rect 227718 490512 227774 490521
rect 227718 490447 227774 490456
rect 228376 469849 228404 530538
rect 229296 526318 229324 539158
rect 229664 534041 229692 539172
rect 230400 534750 230428 539172
rect 230492 539158 230966 539186
rect 230388 534744 230440 534750
rect 230388 534686 230440 534692
rect 229650 534032 229706 534041
rect 229650 533967 229706 533976
rect 229284 526312 229336 526318
rect 229284 526254 229336 526260
rect 229100 522980 229152 522986
rect 229100 522922 229152 522928
rect 228454 493504 228510 493513
rect 228454 493439 228510 493448
rect 228468 469878 228496 493439
rect 229112 472054 229140 522922
rect 230492 511290 230520 539158
rect 231688 535498 231716 539172
rect 231872 539158 232254 539186
rect 232332 539158 232806 539186
rect 233344 539158 233542 539186
rect 233712 539158 234094 539186
rect 234632 539158 234830 539186
rect 231676 535492 231728 535498
rect 231676 535434 231728 535440
rect 231216 534812 231268 534818
rect 231216 534754 231268 534760
rect 231122 522336 231178 522345
rect 231122 522271 231178 522280
rect 230480 511284 230532 511290
rect 230480 511226 230532 511232
rect 229100 472048 229152 472054
rect 229100 471990 229152 471996
rect 228456 469872 228508 469878
rect 228362 469840 228418 469849
rect 228456 469814 228508 469820
rect 228362 469775 228418 469784
rect 227720 468512 227772 468518
rect 227720 468454 227772 468460
rect 227628 463820 227680 463826
rect 227628 463762 227680 463768
rect 226984 455796 227036 455802
rect 226984 455738 227036 455744
rect 227732 451382 227760 468454
rect 227810 464672 227866 464681
rect 227810 464607 227866 464616
rect 227824 454034 227852 464607
rect 229112 460934 229140 471990
rect 229112 460906 229232 460934
rect 227812 454028 227864 454034
rect 227812 453970 227864 453976
rect 228732 454028 228784 454034
rect 228732 453970 228784 453976
rect 227720 451376 227772 451382
rect 227720 451318 227772 451324
rect 227732 450242 227760 451318
rect 225616 450214 225998 450242
rect 226444 450214 226918 450242
rect 227732 450214 227838 450242
rect 207570 450191 207626 450200
rect 205638 450120 205694 450129
rect 228744 450106 228772 453970
rect 229204 450242 229232 460906
rect 231136 459649 231164 522271
rect 231228 496194 231256 534754
rect 231216 496188 231268 496194
rect 231216 496130 231268 496136
rect 231214 491192 231270 491201
rect 231214 491127 231270 491136
rect 231228 467129 231256 491127
rect 231872 479505 231900 539158
rect 232332 528554 232360 539158
rect 233240 533384 233292 533390
rect 232502 533352 232558 533361
rect 233240 533326 233292 533332
rect 232502 533287 232558 533296
rect 231964 528526 232360 528554
rect 231964 480865 231992 528526
rect 232516 504422 232544 533287
rect 232504 504416 232556 504422
rect 232504 504358 232556 504364
rect 232504 486532 232556 486538
rect 232504 486474 232556 486480
rect 231950 480856 232006 480865
rect 231950 480791 232006 480800
rect 231858 479496 231914 479505
rect 231858 479431 231914 479440
rect 231306 474872 231362 474881
rect 231306 474807 231362 474816
rect 231214 467120 231270 467129
rect 231214 467055 231270 467064
rect 231122 459640 231178 459649
rect 231122 459575 231178 459584
rect 230570 455968 230626 455977
rect 230570 455903 230626 455912
rect 230584 450242 230612 455903
rect 231136 451274 231164 459575
rect 231320 455977 231348 474807
rect 231860 461712 231912 461718
rect 231860 461654 231912 461660
rect 231872 460934 231900 461654
rect 231872 460906 232176 460934
rect 232148 458425 232176 460906
rect 232134 458416 232190 458425
rect 232134 458351 232190 458360
rect 231306 455968 231362 455977
rect 231306 455903 231362 455912
rect 231320 455569 231348 455903
rect 231306 455560 231362 455569
rect 231306 455495 231362 455504
rect 231136 451246 231348 451274
rect 231320 450242 231348 451246
rect 232148 450242 232176 458351
rect 232516 453937 232544 486474
rect 233252 483682 233280 533326
rect 233344 515438 233372 539158
rect 233712 533390 233740 539158
rect 233884 535492 233936 535498
rect 233884 535434 233936 535440
rect 233700 533384 233752 533390
rect 233700 533326 233752 533332
rect 233332 515432 233384 515438
rect 233332 515374 233384 515380
rect 233896 497554 233924 535434
rect 234632 500177 234660 539158
rect 235368 533361 235396 539172
rect 236012 539158 236118 539186
rect 235354 533352 235410 533361
rect 235354 533287 235410 533296
rect 234618 500168 234674 500177
rect 234618 500103 234674 500112
rect 233884 497548 233936 497554
rect 233884 497490 233936 497496
rect 235906 496088 235962 496097
rect 235906 496023 235962 496032
rect 233240 483676 233292 483682
rect 233240 483618 233292 483624
rect 233976 455456 234028 455462
rect 233976 455398 234028 455404
rect 232502 453928 232558 453937
rect 232502 453863 232558 453872
rect 233514 453928 233570 453937
rect 233514 453863 233570 453872
rect 233528 451489 233556 453863
rect 233514 451480 233570 451489
rect 233514 451415 233570 451424
rect 229204 450214 229678 450242
rect 230584 450214 230782 450242
rect 231320 450214 231702 450242
rect 232148 450214 232622 450242
rect 233528 450228 233556 451415
rect 233988 450242 234016 455398
rect 235920 454073 235948 496023
rect 236012 486742 236040 539158
rect 236656 533322 236684 539172
rect 236644 533316 236696 533322
rect 236644 533258 236696 533264
rect 237392 504422 237420 539172
rect 237484 539158 237958 539186
rect 237484 525094 237512 539158
rect 238680 538286 238708 539172
rect 238668 538280 238720 538286
rect 238668 538222 238720 538228
rect 238680 533390 238708 538222
rect 239232 536722 239260 539172
rect 239220 536716 239272 536722
rect 239220 536658 239272 536664
rect 239784 534886 239812 539172
rect 240244 539158 240534 539186
rect 240704 539158 241086 539186
rect 241532 539158 241822 539186
rect 241900 539158 242374 539186
rect 242912 539158 243110 539186
rect 239772 534880 239824 534886
rect 239772 534822 239824 534828
rect 239404 533452 239456 533458
rect 239404 533394 239456 533400
rect 238668 533384 238720 533390
rect 238668 533326 238720 533332
rect 238024 529236 238076 529242
rect 238024 529178 238076 529184
rect 237472 525088 237524 525094
rect 237472 525030 237524 525036
rect 237380 504416 237432 504422
rect 237380 504358 237432 504364
rect 236000 486736 236052 486742
rect 236000 486678 236052 486684
rect 238036 465118 238064 529178
rect 238116 486736 238168 486742
rect 238116 486678 238168 486684
rect 237380 465112 237432 465118
rect 237380 465054 237432 465060
rect 238024 465112 238076 465118
rect 238024 465054 238076 465060
rect 235998 462904 236054 462913
rect 235998 462839 236054 462848
rect 234894 454064 234950 454073
rect 234894 453999 234950 454008
rect 235906 454064 235962 454073
rect 235906 453999 235962 454008
rect 234908 450242 234936 453999
rect 236012 450242 236040 462839
rect 237392 460934 237420 465054
rect 237392 460906 237972 460934
rect 237472 456816 237524 456822
rect 237472 456758 237524 456764
rect 237484 450242 237512 456758
rect 233988 450214 234462 450242
rect 234908 450214 235382 450242
rect 236012 450214 236486 450242
rect 237406 450214 237512 450242
rect 237944 450242 237972 460906
rect 238128 456822 238156 486678
rect 239416 482322 239444 533394
rect 240140 532908 240192 532914
rect 240140 532850 240192 532856
rect 239404 482316 239456 482322
rect 239404 482258 239456 482264
rect 239404 469872 239456 469878
rect 239404 469814 239456 469820
rect 238116 456816 238168 456822
rect 238116 456758 238168 456764
rect 239416 453937 239444 469814
rect 240152 456074 240180 532850
rect 240244 515506 240272 539158
rect 240704 532914 240732 539158
rect 240692 532908 240744 532914
rect 240692 532850 240744 532856
rect 240232 515500 240284 515506
rect 240232 515442 240284 515448
rect 240782 481536 240838 481545
rect 240782 481471 240838 481480
rect 240796 480282 240824 481471
rect 240784 480276 240836 480282
rect 240784 480218 240836 480224
rect 240232 470620 240284 470626
rect 240232 470562 240284 470568
rect 240244 468518 240272 470562
rect 240232 468512 240284 468518
rect 240232 468454 240284 468460
rect 240796 460329 240824 480218
rect 241428 469192 241480 469198
rect 241428 469134 241480 469140
rect 241440 468518 241468 469134
rect 241428 468512 241480 468518
rect 241428 468454 241480 468460
rect 241440 460934 241468 468454
rect 241348 460906 241468 460934
rect 240782 460320 240838 460329
rect 240782 460255 240838 460264
rect 240140 456068 240192 456074
rect 240140 456010 240192 456016
rect 239402 453928 239458 453937
rect 239402 453863 239458 453872
rect 239218 451888 239274 451897
rect 239218 451823 239274 451832
rect 239232 451353 239260 451823
rect 239218 451344 239274 451353
rect 241348 451314 241376 460906
rect 241532 458862 241560 539158
rect 241900 528554 241928 539158
rect 242912 529242 242940 539158
rect 243542 538792 243598 538801
rect 243542 538727 243598 538736
rect 242900 529236 242952 529242
rect 242900 529178 242952 529184
rect 241624 528526 241928 528554
rect 241624 485110 241652 528526
rect 241612 485104 241664 485110
rect 241612 485046 241664 485052
rect 243556 483002 243584 538727
rect 243648 535537 243676 539172
rect 244384 538218 244412 539172
rect 244372 538212 244424 538218
rect 244372 538154 244424 538160
rect 244280 537532 244332 537538
rect 244280 537474 244332 537480
rect 244292 536722 244320 537474
rect 244384 536858 244412 538154
rect 244372 536852 244424 536858
rect 244372 536794 244424 536800
rect 244832 536852 244884 536858
rect 244832 536794 244884 536800
rect 244280 536716 244332 536722
rect 244280 536658 244332 536664
rect 243634 535528 243690 535537
rect 243634 535463 243690 535472
rect 244292 528554 244320 536658
rect 244556 533452 244608 533458
rect 244556 533394 244608 533400
rect 244292 528526 244504 528554
rect 244278 518120 244334 518129
rect 244278 518055 244334 518064
rect 242900 482996 242952 483002
rect 242900 482938 242952 482944
rect 243544 482996 243596 483002
rect 243544 482938 243596 482944
rect 242912 481710 242940 482938
rect 242900 481704 242952 481710
rect 242900 481646 242952 481652
rect 242164 469260 242216 469266
rect 242164 469202 242216 469208
rect 241520 458856 241572 458862
rect 241520 458798 241572 458804
rect 241426 456920 241482 456929
rect 241426 456855 241482 456864
rect 241440 453354 241468 456855
rect 241428 453348 241480 453354
rect 241428 453290 241480 453296
rect 242176 452849 242204 469202
rect 242162 452840 242218 452849
rect 242162 452775 242218 452784
rect 239218 451279 239274 451288
rect 240140 451308 240192 451314
rect 237944 450214 238326 450242
rect 239232 450228 239260 451279
rect 240140 451250 240192 451256
rect 241336 451308 241388 451314
rect 241336 451250 241388 451256
rect 240152 450228 240180 451250
rect 240692 451240 240744 451246
rect 240692 451182 240744 451188
rect 240704 450242 240732 451182
rect 240704 450214 241086 450242
rect 242176 450228 242204 452775
rect 242912 450242 242940 481646
rect 244292 462913 244320 518055
rect 244476 502994 244504 528526
rect 244568 522306 244596 533394
rect 244844 528554 244872 536794
rect 244936 536178 244964 539172
rect 245028 539158 245502 539186
rect 244924 536172 244976 536178
rect 244924 536114 244976 536120
rect 245028 533458 245056 539158
rect 245936 536172 245988 536178
rect 245936 536114 245988 536120
rect 245016 533452 245068 533458
rect 245016 533394 245068 533400
rect 244844 528526 244964 528554
rect 244936 527950 244964 528526
rect 244924 527944 244976 527950
rect 244924 527886 244976 527892
rect 244556 522300 244608 522306
rect 244556 522242 244608 522248
rect 244464 502988 244516 502994
rect 244464 502930 244516 502936
rect 244278 462904 244334 462913
rect 244278 462839 244334 462848
rect 242992 462392 243044 462398
rect 242992 462334 243044 462340
rect 243004 455394 243032 462334
rect 245948 460934 245976 536114
rect 246224 532030 246252 539172
rect 246776 536790 246804 539172
rect 246764 536784 246816 536790
rect 246764 536726 246816 536732
rect 247512 535498 247540 539172
rect 247696 539158 248078 539186
rect 248524 539158 248814 539186
rect 248984 539158 249366 539186
rect 247696 538214 247724 539158
rect 247604 538186 247724 538214
rect 246304 535492 246356 535498
rect 246304 535434 246356 535440
rect 247500 535492 247552 535498
rect 247500 535434 247552 535440
rect 246212 532024 246264 532030
rect 246212 531966 246264 531972
rect 246316 489190 246344 535434
rect 247604 530602 247632 538186
rect 248420 533452 248472 533458
rect 248420 533394 248472 533400
rect 247592 530596 247644 530602
rect 247592 530538 247644 530544
rect 247684 530596 247736 530602
rect 247684 530538 247736 530544
rect 247696 507142 247724 530538
rect 247684 507136 247736 507142
rect 247684 507078 247736 507084
rect 248432 491978 248460 533394
rect 248524 525094 248552 539158
rect 248984 533458 249012 539158
rect 249708 536852 249760 536858
rect 249708 536794 249760 536800
rect 248972 533452 249024 533458
rect 248972 533394 249024 533400
rect 248604 527876 248656 527882
rect 248604 527818 248656 527824
rect 248512 525088 248564 525094
rect 248512 525030 248564 525036
rect 248420 491972 248472 491978
rect 248420 491914 248472 491920
rect 246304 489184 246356 489190
rect 246304 489126 246356 489132
rect 247130 485072 247186 485081
rect 247130 485007 247186 485016
rect 246948 471300 247000 471306
rect 246948 471242 247000 471248
rect 246960 468586 246988 471242
rect 246948 468580 247000 468586
rect 246948 468522 247000 468528
rect 245948 460906 246160 460934
rect 244922 460184 244978 460193
rect 244922 460119 244978 460128
rect 242992 455388 243044 455394
rect 242992 455330 243044 455336
rect 243544 455388 243596 455394
rect 243544 455330 243596 455336
rect 243556 450242 243584 455330
rect 244936 452713 244964 460119
rect 244922 452704 244978 452713
rect 244922 452639 244978 452648
rect 242912 450214 243110 450242
rect 243556 450214 244030 450242
rect 244936 450228 244964 452639
rect 245934 450256 245990 450265
rect 245870 450214 245934 450242
rect 245934 450191 245990 450200
rect 228822 450120 228878 450129
rect 205694 450078 205942 450106
rect 228744 450092 228822 450106
rect 228758 450078 228822 450092
rect 205638 450055 205694 450064
rect 228822 450055 228878 450064
rect 204166 449984 204222 449993
rect 204088 449956 204166 449970
rect 204102 449942 204166 449956
rect 204166 449919 204222 449928
rect 195336 449812 195388 449818
rect 195336 449754 195388 449760
rect 194508 449744 194560 449750
rect 246132 449721 246160 460906
rect 246396 457496 246448 457502
rect 246396 457438 246448 457444
rect 246408 450242 246436 457438
rect 246408 450214 246790 450242
rect 247144 449721 247172 485007
rect 248616 463758 248644 527818
rect 249064 473408 249116 473414
rect 249064 473350 249116 473356
rect 248420 463752 248472 463758
rect 248420 463694 248472 463700
rect 248604 463752 248656 463758
rect 248604 463694 248656 463700
rect 247500 457496 247552 457502
rect 247500 457438 247552 457444
rect 247512 450242 247540 457438
rect 248432 450242 248460 463694
rect 249076 456113 249104 473350
rect 249720 471306 249748 536794
rect 250088 533361 250116 539172
rect 250180 539158 250654 539186
rect 251192 539158 251390 539186
rect 250074 533352 250130 533361
rect 250074 533287 250130 533296
rect 250180 528554 250208 539158
rect 250444 533452 250496 533458
rect 250444 533394 250496 533400
rect 249812 528526 250208 528554
rect 249812 527105 249840 528526
rect 249798 527096 249854 527105
rect 249798 527031 249854 527040
rect 250456 497486 250484 533394
rect 250444 497480 250496 497486
rect 250444 497422 250496 497428
rect 250442 485888 250498 485897
rect 250442 485823 250498 485832
rect 249800 483676 249852 483682
rect 249800 483618 249852 483624
rect 249708 471300 249760 471306
rect 249708 471242 249760 471248
rect 249812 460222 249840 483618
rect 249800 460216 249852 460222
rect 249800 460158 249852 460164
rect 249616 459604 249668 459610
rect 249616 459546 249668 459552
rect 249062 456104 249118 456113
rect 249062 456039 249118 456048
rect 249076 451274 249104 456039
rect 249628 454034 249656 459546
rect 249616 454028 249668 454034
rect 249616 453970 249668 453976
rect 250456 452169 250484 485823
rect 251192 471170 251220 539158
rect 251928 534750 251956 539172
rect 252020 539158 252494 539186
rect 251916 534744 251968 534750
rect 251916 534686 251968 534692
rect 252020 533338 252048 539158
rect 252100 538348 252152 538354
rect 252100 538290 252152 538296
rect 251284 533310 252048 533338
rect 251284 514078 251312 533310
rect 252112 528554 252140 538290
rect 251836 528526 252140 528554
rect 253124 528554 253152 539310
rect 253216 536081 253244 539172
rect 253202 536072 253258 536081
rect 253202 536007 253258 536016
rect 253124 528526 253244 528554
rect 251456 515432 251508 515438
rect 251456 515374 251508 515380
rect 251272 514072 251324 514078
rect 251272 514014 251324 514020
rect 251362 492688 251418 492697
rect 251362 492623 251418 492632
rect 251376 474774 251404 492623
rect 251468 478174 251496 515374
rect 251836 487830 251864 528526
rect 253216 509998 253244 528526
rect 253204 509992 253256 509998
rect 253204 509934 253256 509940
rect 253204 504416 253256 504422
rect 253204 504358 253256 504364
rect 251824 487824 251876 487830
rect 251824 487766 251876 487772
rect 251456 478168 251508 478174
rect 251456 478110 251508 478116
rect 251468 477562 251496 478110
rect 251456 477556 251508 477562
rect 251456 477498 251508 477504
rect 251916 477556 251968 477562
rect 251916 477498 251968 477504
rect 251364 474768 251416 474774
rect 251364 474710 251416 474716
rect 251180 471164 251232 471170
rect 251180 471106 251232 471112
rect 251192 470694 251220 471106
rect 251180 470688 251232 470694
rect 251180 470630 251232 470636
rect 251376 470594 251404 474710
rect 251824 471164 251876 471170
rect 251824 471106 251876 471112
rect 251284 470566 251404 470594
rect 251086 466576 251142 466585
rect 251086 466511 251142 466520
rect 251100 465905 251128 466511
rect 251086 465896 251142 465905
rect 251086 465831 251142 465840
rect 251180 462324 251232 462330
rect 251180 462266 251232 462272
rect 251192 460970 251220 462266
rect 251180 460964 251232 460970
rect 251180 460906 251232 460912
rect 250442 452160 250498 452169
rect 250442 452095 250498 452104
rect 249076 451246 249288 451274
rect 249260 450242 249288 451246
rect 251192 450242 251220 460906
rect 251284 456142 251312 470566
rect 251272 456136 251324 456142
rect 251272 456078 251324 456084
rect 251836 451042 251864 471106
rect 251928 462330 251956 477498
rect 251916 462324 251968 462330
rect 251916 462266 251968 462272
rect 253216 458930 253244 504358
rect 253308 500342 253336 586486
rect 253386 556200 253442 556209
rect 253386 556135 253442 556144
rect 253296 500336 253348 500342
rect 253296 500278 253348 500284
rect 253400 481545 253428 556135
rect 253952 538801 253980 587347
rect 254044 582321 254072 611322
rect 254584 603220 254636 603226
rect 254584 603162 254636 603168
rect 254596 589966 254624 603162
rect 255318 603120 255374 603129
rect 255318 603055 255374 603064
rect 255332 594289 255360 603055
rect 255976 598913 256004 702442
rect 267660 697610 267688 703520
rect 274548 703112 274600 703118
rect 274548 703054 274600 703060
rect 269304 702840 269356 702846
rect 269304 702782 269356 702788
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 258080 612808 258132 612814
rect 258080 612750 258132 612756
rect 256700 610020 256752 610026
rect 256700 609962 256752 609968
rect 256056 598936 256108 598942
rect 255962 598904 256018 598913
rect 256056 598878 256108 598884
rect 255962 598839 256018 598848
rect 255410 597680 255466 597689
rect 255410 597615 255412 597624
rect 255464 597615 255466 597624
rect 255412 597586 255464 597592
rect 255410 596592 255466 596601
rect 255410 596527 255466 596536
rect 255424 596222 255452 596527
rect 255412 596216 255464 596222
rect 255412 596158 255464 596164
rect 255318 594280 255374 594289
rect 255318 594215 255374 594224
rect 255332 594114 255360 594215
rect 255320 594108 255372 594114
rect 255320 594050 255372 594056
rect 255410 591016 255466 591025
rect 255410 590951 255466 590960
rect 255424 590714 255452 590951
rect 255412 590708 255464 590714
rect 255412 590650 255464 590656
rect 254584 589960 254636 589966
rect 254584 589902 254636 589908
rect 255410 589928 255466 589937
rect 255410 589863 255466 589872
rect 255424 589354 255452 589863
rect 255412 589348 255464 589354
rect 255412 589290 255464 589296
rect 255410 588160 255466 588169
rect 255410 588095 255466 588104
rect 255424 587926 255452 588095
rect 255412 587920 255464 587926
rect 255412 587862 255464 587868
rect 255410 585168 255466 585177
rect 255410 585103 255466 585112
rect 255320 584452 255372 584458
rect 255320 584394 255372 584400
rect 255332 584225 255360 584394
rect 255318 584216 255374 584225
rect 255318 584151 255374 584160
rect 255424 584066 255452 585103
rect 255332 584038 255452 584066
rect 254030 582312 254086 582321
rect 254030 582247 254086 582256
rect 254030 577552 254086 577561
rect 254030 577487 254086 577496
rect 253938 538792 253994 538801
rect 253938 538727 253994 538736
rect 254044 534818 254072 577487
rect 254122 547904 254178 547913
rect 254122 547839 254178 547848
rect 254136 536858 254164 547839
rect 254214 542464 254270 542473
rect 254214 542399 254270 542408
rect 254124 536852 254176 536858
rect 254124 536794 254176 536800
rect 254032 534812 254084 534818
rect 254032 534754 254084 534760
rect 253938 507920 253994 507929
rect 253938 507855 253994 507864
rect 253952 501634 253980 507855
rect 254228 505782 254256 542399
rect 254216 505776 254268 505782
rect 254216 505718 254268 505724
rect 253940 501628 253992 501634
rect 253940 501570 253992 501576
rect 253386 481536 253442 481545
rect 253386 481471 253442 481480
rect 254124 479528 254176 479534
rect 254124 479470 254176 479476
rect 253480 473476 253532 473482
rect 253480 473418 253532 473424
rect 253204 458924 253256 458930
rect 253204 458866 253256 458872
rect 252100 456136 252152 456142
rect 252100 456078 252152 456084
rect 251914 451480 251970 451489
rect 251914 451415 251970 451424
rect 251824 451036 251876 451042
rect 251824 450978 251876 450984
rect 247512 450214 247894 450242
rect 248432 450214 248814 450242
rect 249260 450214 249734 450242
rect 251192 450214 251574 450242
rect 250654 449954 250944 449970
rect 250654 449948 250956 449954
rect 250654 449942 250904 449948
rect 250904 449890 250956 449896
rect 251928 449750 251956 451415
rect 252112 450242 252140 456078
rect 253388 454028 253440 454034
rect 253388 453970 253440 453976
rect 252112 450214 252494 450242
rect 253400 450228 253428 453970
rect 251916 449744 251968 449750
rect 194508 449686 194560 449692
rect 246118 449712 246174 449721
rect 246118 449647 246174 449656
rect 247130 449712 247186 449721
rect 251916 449686 251968 449692
rect 247130 449647 247186 449656
rect 253492 448066 253520 473418
rect 253938 472152 253994 472161
rect 253938 472087 253994 472096
rect 253952 471209 253980 472087
rect 253938 471200 253994 471209
rect 253938 471135 253994 471144
rect 254032 458856 254084 458862
rect 254032 458798 254084 458804
rect 253572 456816 253624 456822
rect 253572 456758 253624 456764
rect 253584 448610 253612 456758
rect 253584 448582 253980 448610
rect 253570 448080 253626 448089
rect 253492 448038 253570 448066
rect 253570 448015 253626 448024
rect 193312 440904 193364 440910
rect 193312 440846 193364 440852
rect 253572 423428 253624 423434
rect 253572 423370 253624 423376
rect 193126 419792 193182 419801
rect 193126 419727 193182 419736
rect 253584 413681 253612 423370
rect 253570 413672 253626 413681
rect 253570 413607 253626 413616
rect 192574 413264 192630 413273
rect 192574 413199 192630 413208
rect 192482 408640 192538 408649
rect 192482 408575 192538 408584
rect 192496 327214 192524 408575
rect 192588 384946 192616 413199
rect 193312 407788 193364 407794
rect 193312 407730 193364 407736
rect 192668 396092 192720 396098
rect 192668 396034 192720 396040
rect 192680 391105 192708 396034
rect 193220 391332 193272 391338
rect 193220 391274 193272 391280
rect 192666 391096 192722 391105
rect 192666 391031 192722 391040
rect 193232 390998 193260 391274
rect 193220 390992 193272 390998
rect 193126 390960 193182 390969
rect 193220 390934 193272 390940
rect 193126 390895 193182 390904
rect 193140 389473 193168 390895
rect 193126 389464 193182 389473
rect 193126 389399 193182 389408
rect 192576 384940 192628 384946
rect 192576 384882 192628 384888
rect 192484 327208 192536 327214
rect 192484 327150 192536 327156
rect 193324 320929 193352 407730
rect 253572 398200 253624 398206
rect 253572 398142 253624 398148
rect 253584 393314 253612 398142
rect 253492 393286 253612 393314
rect 193402 391096 193458 391105
rect 193458 391054 193614 391082
rect 193402 391031 193458 391040
rect 194140 390992 194192 390998
rect 218336 390992 218388 390998
rect 194192 390940 194534 390946
rect 194140 390934 194534 390940
rect 218336 390934 218388 390940
rect 218796 390992 218848 390998
rect 251732 390992 251784 390998
rect 248878 390960 248934 390969
rect 218848 390940 219190 390946
rect 218796 390934 219190 390940
rect 194152 390918 194534 390934
rect 194612 390374 195454 390402
rect 195992 390374 196374 390402
rect 194138 389872 194194 389881
rect 194138 389807 194194 389816
rect 194152 386374 194180 389807
rect 194140 386368 194192 386374
rect 194140 386310 194192 386316
rect 194612 358698 194640 390374
rect 195992 387818 196020 390374
rect 197280 389162 197308 390388
rect 197268 389156 197320 389162
rect 197268 389098 197320 389104
rect 197280 387870 197308 389098
rect 195900 387790 196020 387818
rect 196072 387864 196124 387870
rect 196072 387806 196124 387812
rect 197268 387864 197320 387870
rect 197268 387806 197320 387812
rect 195900 385694 195928 387790
rect 195888 385688 195940 385694
rect 195888 385630 195940 385636
rect 196084 373994 196112 387806
rect 198200 387705 198228 390388
rect 198752 390374 199134 390402
rect 198186 387696 198242 387705
rect 198186 387631 198242 387640
rect 198752 383625 198780 390374
rect 200224 386073 200252 390388
rect 201144 386345 201172 390388
rect 202064 389298 202092 390388
rect 202052 389292 202104 389298
rect 202052 389234 202104 389240
rect 202984 387734 203012 390388
rect 203168 390374 203918 390402
rect 202972 387728 203024 387734
rect 202972 387670 203024 387676
rect 201130 386336 201186 386345
rect 201130 386271 201186 386280
rect 200210 386064 200266 386073
rect 200210 385999 200266 386008
rect 198830 384432 198886 384441
rect 198830 384367 198886 384376
rect 198738 383616 198794 383625
rect 198738 383551 198794 383560
rect 198752 382945 198780 383551
rect 198738 382936 198794 382945
rect 198738 382871 198794 382880
rect 197452 378888 197504 378894
rect 197452 378830 197504 378836
rect 195992 373966 196112 373994
rect 195992 362273 196020 373966
rect 195978 362264 196034 362273
rect 195978 362199 196034 362208
rect 195992 359514 196020 362199
rect 195980 359508 196032 359514
rect 195980 359450 196032 359456
rect 194600 358692 194652 358698
rect 194600 358634 194652 358640
rect 195242 358048 195298 358057
rect 195242 357983 195298 357992
rect 193310 320920 193366 320929
rect 193310 320855 193366 320864
rect 192484 309596 192536 309602
rect 192484 309538 192536 309544
rect 192022 296032 192078 296041
rect 192022 295967 192078 295976
rect 192036 295361 192064 295967
rect 192022 295352 192078 295361
rect 192022 295287 192078 295296
rect 192496 291825 192524 309538
rect 195256 308446 195284 357983
rect 196622 341456 196678 341465
rect 196622 341391 196678 341400
rect 195978 316704 196034 316713
rect 195978 316639 196034 316648
rect 195426 316160 195482 316169
rect 195426 316095 195482 316104
rect 195334 315344 195390 315353
rect 195334 315279 195390 315288
rect 195244 308440 195296 308446
rect 195244 308382 195296 308388
rect 193864 306468 193916 306474
rect 193864 306410 193916 306416
rect 192942 301880 192998 301889
rect 192942 301815 192998 301824
rect 192956 296993 192984 301815
rect 193770 301744 193826 301753
rect 193770 301679 193826 301688
rect 193128 300960 193180 300966
rect 193128 300902 193180 300908
rect 193140 298897 193168 300902
rect 193494 300792 193550 300801
rect 193494 300727 193550 300736
rect 193508 300121 193536 300727
rect 193494 300112 193550 300121
rect 193494 300047 193550 300056
rect 193678 300112 193734 300121
rect 193678 300047 193734 300056
rect 193692 299674 193720 300047
rect 193680 299668 193732 299674
rect 193680 299610 193732 299616
rect 193126 298888 193182 298897
rect 193126 298823 193182 298832
rect 192942 296984 192998 296993
rect 192942 296919 192998 296928
rect 193678 295216 193734 295225
rect 193784 295202 193812 301679
rect 193876 301580 193904 306410
rect 194416 305040 194468 305046
rect 194416 304982 194468 304988
rect 194428 301580 194456 304982
rect 195348 301889 195376 315279
rect 195440 305658 195468 316095
rect 195992 309369 196020 316639
rect 195978 309360 196034 309369
rect 195978 309295 196034 309304
rect 195428 305652 195480 305658
rect 195428 305594 195480 305600
rect 195612 303748 195664 303754
rect 195612 303690 195664 303696
rect 195334 301880 195390 301889
rect 195334 301815 195390 301824
rect 195058 301744 195114 301753
rect 195058 301679 195114 301688
rect 195072 301580 195100 301679
rect 195624 301580 195652 303690
rect 195992 303618 196020 309295
rect 195980 303612 196032 303618
rect 195980 303554 196032 303560
rect 195978 300928 196034 300937
rect 196636 300914 196664 341391
rect 197464 325694 197492 378830
rect 198740 345160 198792 345166
rect 198740 345102 198792 345108
rect 197464 325666 197584 325694
rect 197358 320784 197414 320793
rect 197358 320719 197414 320728
rect 197372 305250 197400 320719
rect 197556 306374 197584 325666
rect 198752 306374 198780 345102
rect 198844 309602 198872 384367
rect 203168 373994 203196 390374
rect 204824 389201 204852 390388
rect 205744 390374 205942 390402
rect 206480 390374 206862 390402
rect 207032 390374 207782 390402
rect 208504 390374 208702 390402
rect 209240 390374 209622 390402
rect 209792 390374 210542 390402
rect 211172 390374 211646 390402
rect 204810 389192 204866 389201
rect 204810 389127 204866 389136
rect 204824 388793 204852 389127
rect 204810 388784 204866 388793
rect 204810 388719 204866 388728
rect 204824 383654 204852 388719
rect 205640 387048 205692 387054
rect 205640 386990 205692 386996
rect 204824 383626 204944 383654
rect 202984 373966 203196 373994
rect 202984 356046 203012 373966
rect 202972 356040 203024 356046
rect 202972 355982 203024 355988
rect 202144 342372 202196 342378
rect 202144 342314 202196 342320
rect 200762 338736 200818 338745
rect 200762 338671 200818 338680
rect 200776 313313 200804 338671
rect 201682 336288 201738 336297
rect 201682 336223 201738 336232
rect 201498 331800 201554 331809
rect 201498 331735 201554 331744
rect 200210 313304 200266 313313
rect 200210 313239 200266 313248
rect 200762 313304 200818 313313
rect 200762 313239 200818 313248
rect 198832 309596 198884 309602
rect 198832 309538 198884 309544
rect 199384 309596 199436 309602
rect 199384 309538 199436 309544
rect 197556 306346 197676 306374
rect 198752 306346 198872 306374
rect 197360 305244 197412 305250
rect 197360 305186 197412 305192
rect 197360 305108 197412 305114
rect 197360 305050 197412 305056
rect 196716 303612 196768 303618
rect 196716 303554 196768 303560
rect 196728 301594 196756 303554
rect 197372 301594 197400 305050
rect 196728 301566 196834 301594
rect 197372 301566 197478 301594
rect 197648 300966 197676 306346
rect 198738 305688 198794 305697
rect 198738 305623 198794 305632
rect 198372 305244 198424 305250
rect 198372 305186 198424 305192
rect 198384 301594 198412 305186
rect 198752 304337 198780 305623
rect 198738 304328 198794 304337
rect 198738 304263 198794 304272
rect 198752 303754 198780 304263
rect 198740 303748 198792 303754
rect 198740 303690 198792 303696
rect 198844 301594 198872 306346
rect 199396 301594 199424 309538
rect 200224 301594 200252 313239
rect 201040 303748 201092 303754
rect 201040 303690 201092 303696
rect 198384 301566 198674 301594
rect 198844 301566 199226 301594
rect 199396 301566 199870 301594
rect 200224 301566 200422 301594
rect 201052 301580 201080 303690
rect 201512 303618 201540 331735
rect 201592 329928 201644 329934
rect 201592 329870 201644 329876
rect 201604 306374 201632 329870
rect 201696 329225 201724 336223
rect 201682 329216 201738 329225
rect 201682 329151 201738 329160
rect 202050 323640 202106 323649
rect 202050 323575 202106 323584
rect 202064 306374 202092 323575
rect 202156 307766 202184 342314
rect 204258 326360 204314 326369
rect 204258 326295 204314 326304
rect 203062 318880 203118 318889
rect 203062 318815 203118 318824
rect 202144 307760 202196 307766
rect 202144 307702 202196 307708
rect 201604 306346 201724 306374
rect 202064 306346 202368 306374
rect 201500 303612 201552 303618
rect 201500 303554 201552 303560
rect 201696 301594 201724 306346
rect 201868 303612 201920 303618
rect 201868 303554 201920 303560
rect 201618 301566 201724 301594
rect 201880 301594 201908 303554
rect 202340 301594 202368 306346
rect 203076 301594 203104 318815
rect 203984 307760 204036 307766
rect 203984 307702 204036 307708
rect 201880 301566 202262 301594
rect 202340 301566 202814 301594
rect 203076 301566 203458 301594
rect 203996 301580 204024 307702
rect 204272 301594 204300 326295
rect 204916 319433 204944 383626
rect 205652 354686 205680 386990
rect 205744 378078 205772 390374
rect 206480 387054 206508 390374
rect 206468 387048 206520 387054
rect 206468 386990 206520 386996
rect 207032 380186 207060 390374
rect 208400 387048 208452 387054
rect 208400 386990 208452 386996
rect 207020 380180 207072 380186
rect 207020 380122 207072 380128
rect 205732 378072 205784 378078
rect 205732 378014 205784 378020
rect 208412 373289 208440 386990
rect 208504 383042 208532 390374
rect 209240 387054 209268 390374
rect 209228 387048 209280 387054
rect 209228 386990 209280 386996
rect 208492 383036 208544 383042
rect 208492 382978 208544 382984
rect 208398 373280 208454 373289
rect 208398 373215 208454 373224
rect 209044 371884 209096 371890
rect 209044 371826 209096 371832
rect 206374 356688 206430 356697
rect 206374 356623 206430 356632
rect 205640 354680 205692 354686
rect 205640 354622 205692 354628
rect 205652 352646 205680 354622
rect 205640 352640 205692 352646
rect 205640 352582 205692 352588
rect 204996 351212 205048 351218
rect 204996 351154 205048 351160
rect 204718 319424 204774 319433
rect 204718 319359 204774 319368
rect 204902 319424 204958 319433
rect 204902 319359 204958 319368
rect 204732 301594 204760 319359
rect 205008 315353 205036 351154
rect 206282 349752 206338 349761
rect 206282 349687 206338 349696
rect 205640 334008 205692 334014
rect 205640 333950 205692 333956
rect 205652 333334 205680 333950
rect 205640 333328 205692 333334
rect 205640 333270 205692 333276
rect 205638 328400 205694 328409
rect 205638 328335 205694 328344
rect 205652 327457 205680 328335
rect 205638 327448 205694 327457
rect 205638 327383 205694 327392
rect 205652 325694 205680 327383
rect 205652 325666 206048 325694
rect 204994 315344 205050 315353
rect 204994 315279 205050 315288
rect 205822 305144 205878 305153
rect 205822 305079 205878 305088
rect 204272 301566 204654 301594
rect 204732 301566 205206 301594
rect 205836 301580 205864 305079
rect 206020 301594 206048 325666
rect 206296 305153 206324 349687
rect 206388 328409 206416 356623
rect 207294 333432 207350 333441
rect 207294 333367 207350 333376
rect 207110 329896 207166 329905
rect 207110 329831 207166 329840
rect 206374 328400 206430 328409
rect 206374 328335 206430 328344
rect 206282 305144 206338 305153
rect 206282 305079 206338 305088
rect 207124 301594 207152 329831
rect 206020 301566 206402 301594
rect 207046 301566 207152 301594
rect 207308 301594 207336 333367
rect 208398 331256 208454 331265
rect 208398 331191 208454 331200
rect 208214 302560 208270 302569
rect 208214 302495 208270 302504
rect 207308 301566 207598 301594
rect 208228 301580 208256 302495
rect 208412 301594 208440 331191
rect 209056 323649 209084 371826
rect 209792 369073 209820 390374
rect 211172 382226 211200 390374
rect 212552 389473 212580 390388
rect 212538 389464 212594 389473
rect 212538 389399 212594 389408
rect 213182 385656 213238 385665
rect 213182 385591 213238 385600
rect 211160 382220 211212 382226
rect 211160 382162 211212 382168
rect 211172 380934 211200 382162
rect 211160 380928 211212 380934
rect 211160 380870 211212 380876
rect 211804 380928 211856 380934
rect 211804 380870 211856 380876
rect 209778 369064 209834 369073
rect 209778 368999 209834 369008
rect 211816 365022 211844 380870
rect 212630 378720 212686 378729
rect 212630 378655 212686 378664
rect 211804 365016 211856 365022
rect 211804 364958 211856 364964
rect 211802 359408 211858 359417
rect 211802 359343 211858 359352
rect 209136 342916 209188 342922
rect 209136 342858 209188 342864
rect 209042 323640 209098 323649
rect 209042 323575 209098 323584
rect 209148 321609 209176 342858
rect 209780 327752 209832 327758
rect 209780 327694 209832 327700
rect 209792 324426 209820 327694
rect 211816 325694 211844 359343
rect 212538 333296 212594 333305
rect 212538 333231 212594 333240
rect 211816 325666 212120 325694
rect 209780 324420 209832 324426
rect 209780 324362 209832 324368
rect 210240 324420 210292 324426
rect 210240 324362 210292 324368
rect 208490 321600 208546 321609
rect 208490 321535 208546 321544
rect 209134 321600 209190 321609
rect 209134 321535 209190 321544
rect 208504 306374 208532 321535
rect 208582 318200 208638 318209
rect 208582 318135 208638 318144
rect 208596 313993 208624 318135
rect 208582 313984 208638 313993
rect 208582 313919 208638 313928
rect 210056 307828 210108 307834
rect 210056 307770 210108 307776
rect 208504 306346 208992 306374
rect 208964 301594 208992 306346
rect 208412 301566 208886 301594
rect 208964 301566 209438 301594
rect 210068 301580 210096 307770
rect 210252 301594 210280 324362
rect 211342 312080 211398 312089
rect 211342 312015 211398 312024
rect 211250 311128 211306 311137
rect 211250 311063 211306 311072
rect 210252 301566 210634 301594
rect 211264 301580 211292 311063
rect 211356 301594 211384 312015
rect 212092 303686 212120 325666
rect 212552 306374 212580 333231
rect 212644 325694 212672 378655
rect 213196 375358 213224 385591
rect 213472 384305 213500 390388
rect 213932 390374 214406 390402
rect 213458 384296 213514 384305
rect 213458 384231 213514 384240
rect 213184 375352 213236 375358
rect 213184 375294 213236 375300
rect 213932 373930 213960 390374
rect 215312 385014 215340 390388
rect 215956 390374 216246 390402
rect 216692 390374 217350 390402
rect 218072 390374 218270 390402
rect 215956 387802 215984 390374
rect 215944 387796 215996 387802
rect 215944 387738 215996 387744
rect 215300 385008 215352 385014
rect 215300 384950 215352 384956
rect 215312 384334 215340 384950
rect 215300 384328 215352 384334
rect 215300 384270 215352 384276
rect 213920 373924 213972 373930
rect 213920 373866 213972 373872
rect 212816 362228 212868 362234
rect 212816 362170 212868 362176
rect 212828 356726 212856 362170
rect 212816 356720 212868 356726
rect 212816 356662 212868 356668
rect 214562 353968 214618 353977
rect 214562 353903 214618 353912
rect 214378 345808 214434 345817
rect 214378 345743 214434 345752
rect 214392 341601 214420 345743
rect 214378 341592 214434 341601
rect 214378 341527 214434 341536
rect 213918 334792 213974 334801
rect 213918 334727 213974 334736
rect 212644 325666 213132 325694
rect 213104 314809 213132 325666
rect 213090 314800 213146 314809
rect 213090 314735 213146 314744
rect 212552 306346 212672 306374
rect 212080 303680 212132 303686
rect 212080 303622 212132 303628
rect 212092 301594 212120 303622
rect 212644 301594 212672 306346
rect 213104 301594 213132 314735
rect 213182 313440 213238 313449
rect 213182 313375 213238 313384
rect 213196 304298 213224 313375
rect 213826 306776 213882 306785
rect 213826 306711 213882 306720
rect 213184 304292 213236 304298
rect 213184 304234 213236 304240
rect 213840 303890 213868 306711
rect 213828 303884 213880 303890
rect 213828 303826 213880 303832
rect 213932 303686 213960 334727
rect 214576 318753 214604 353903
rect 215956 338842 215984 387738
rect 216036 384328 216088 384334
rect 216036 384270 216088 384276
rect 216048 347138 216076 384270
rect 216692 381546 216720 390374
rect 216680 381540 216732 381546
rect 216680 381482 216732 381488
rect 218072 374066 218100 390374
rect 218348 381721 218376 390934
rect 218808 390918 219190 390934
rect 248630 390932 248878 390946
rect 248616 390918 248878 390932
rect 220096 386209 220124 390388
rect 220832 390374 221030 390402
rect 221568 390374 221950 390402
rect 220832 386322 220860 390374
rect 221568 388929 221596 390374
rect 221554 388920 221610 388929
rect 221554 388855 221610 388864
rect 221464 387864 221516 387870
rect 221464 387806 221516 387812
rect 220740 386294 220860 386322
rect 220082 386200 220138 386209
rect 220082 386135 220138 386144
rect 218794 384296 218850 384305
rect 218794 384231 218850 384240
rect 218334 381712 218390 381721
rect 218334 381647 218390 381656
rect 218060 374060 218112 374066
rect 218060 374002 218112 374008
rect 218072 371142 218100 374002
rect 218060 371136 218112 371142
rect 218060 371078 218112 371084
rect 218704 366376 218756 366382
rect 218704 366318 218756 366324
rect 217414 355328 217470 355337
rect 217414 355263 217470 355272
rect 216036 347132 216088 347138
rect 216036 347074 216088 347080
rect 217322 344312 217378 344321
rect 217322 344247 217378 344256
rect 215944 338836 215996 338842
rect 215944 338778 215996 338784
rect 215300 338156 215352 338162
rect 215300 338098 215352 338104
rect 214010 318744 214066 318753
rect 214010 318679 214066 318688
rect 214562 318744 214618 318753
rect 214562 318679 214618 318688
rect 214024 317529 214052 318679
rect 214010 317520 214066 317529
rect 214010 317455 214066 317464
rect 213920 303680 213972 303686
rect 213920 303622 213972 303628
rect 214024 301594 214052 317455
rect 214564 303680 214616 303686
rect 214564 303622 214616 303628
rect 214576 301594 214604 303622
rect 215312 301594 215340 338098
rect 215576 337408 215628 337414
rect 215576 337350 215628 337356
rect 215484 336048 215536 336054
rect 215484 335990 215536 335996
rect 215496 306374 215524 335990
rect 215588 325694 215616 337350
rect 216678 329760 216734 329769
rect 216678 329695 216734 329704
rect 216692 328681 216720 329695
rect 216678 328672 216734 328681
rect 216678 328607 216734 328616
rect 215588 325666 216168 325694
rect 215496 306346 215616 306374
rect 215588 301594 215616 306346
rect 216140 301594 216168 325666
rect 216692 306374 216720 328607
rect 216692 306346 217272 306374
rect 217138 305280 217194 305289
rect 217138 305215 217194 305224
rect 217152 301594 217180 305215
rect 217244 303498 217272 306346
rect 217336 305289 217364 344247
rect 217428 329769 217456 355263
rect 217414 329760 217470 329769
rect 217414 329695 217470 329704
rect 218716 328438 218744 366318
rect 218808 355978 218836 384231
rect 218796 355972 218848 355978
rect 218796 355914 218848 355920
rect 219438 334656 219494 334665
rect 219438 334591 219494 334600
rect 219346 329080 219402 329089
rect 219346 329015 219402 329024
rect 218152 328432 218204 328438
rect 218152 328374 218204 328380
rect 218704 328432 218756 328438
rect 218704 328374 218756 328380
rect 218164 327146 218192 328374
rect 218152 327140 218204 327146
rect 218152 327082 218204 327088
rect 218164 325694 218192 327082
rect 218164 325666 218560 325694
rect 217322 305280 217378 305289
rect 217322 305215 217378 305224
rect 217244 303470 217456 303498
rect 217428 301594 217456 303470
rect 218428 302320 218480 302326
rect 218428 302262 218480 302268
rect 211356 301566 211830 301594
rect 212092 301566 212474 301594
rect 212644 301566 213026 301594
rect 213104 301566 213670 301594
rect 214024 301566 214222 301594
rect 214576 301566 214866 301594
rect 215312 301566 215418 301594
rect 215588 301566 216062 301594
rect 216140 301566 216614 301594
rect 217152 301566 217258 301594
rect 217428 301566 217810 301594
rect 218440 301580 218468 302262
rect 218532 301594 218560 325666
rect 219360 302326 219388 329015
rect 219452 303686 219480 334591
rect 219530 329216 219586 329225
rect 219530 329151 219586 329160
rect 219440 303680 219492 303686
rect 219440 303622 219492 303628
rect 219348 302320 219400 302326
rect 219348 302262 219400 302268
rect 219544 301594 219572 329151
rect 220096 315353 220124 386135
rect 220740 377913 220768 386294
rect 220726 377904 220782 377913
rect 220726 377839 220782 377848
rect 221476 365634 221504 387806
rect 221568 380186 221596 388855
rect 222856 384946 222884 390388
rect 223960 387870 223988 390388
rect 223948 387864 224000 387870
rect 223948 387806 224000 387812
rect 224880 386306 224908 390388
rect 225800 386345 225828 390388
rect 226352 390374 226734 390402
rect 224958 386336 225014 386345
rect 224868 386300 224920 386306
rect 224958 386271 225014 386280
rect 225786 386336 225842 386345
rect 225786 386271 225842 386280
rect 224868 386242 224920 386248
rect 222844 384940 222896 384946
rect 222844 384882 222896 384888
rect 221556 380180 221608 380186
rect 221556 380122 221608 380128
rect 221464 365628 221516 365634
rect 221464 365570 221516 365576
rect 221476 337414 221504 365570
rect 222856 355366 222884 384882
rect 222934 364984 222990 364993
rect 222934 364919 222990 364928
rect 222844 355360 222896 355366
rect 222844 355302 222896 355308
rect 222948 351218 222976 364919
rect 222936 351212 222988 351218
rect 222936 351154 222988 351160
rect 224222 343088 224278 343097
rect 224222 343023 224278 343032
rect 222200 338768 222252 338774
rect 222200 338710 222252 338716
rect 221464 337408 221516 337414
rect 221464 337350 221516 337356
rect 222106 334656 222162 334665
rect 222106 334591 222162 334600
rect 222120 327185 222148 334591
rect 221002 327176 221058 327185
rect 221002 327111 221058 327120
rect 222106 327176 222162 327185
rect 222106 327111 222162 327120
rect 220082 315344 220138 315353
rect 220082 315279 220138 315288
rect 219900 303680 219952 303686
rect 219900 303622 219952 303628
rect 219912 301594 219940 303622
rect 220820 302932 220872 302938
rect 220820 302874 220872 302880
rect 220832 302297 220860 302874
rect 220818 302288 220874 302297
rect 220818 302223 220874 302232
rect 218532 301566 219006 301594
rect 219544 301566 219650 301594
rect 219912 301566 220202 301594
rect 220832 301580 220860 302223
rect 221016 301594 221044 327111
rect 222016 303884 222068 303890
rect 222016 303826 222068 303832
rect 221016 301566 221398 301594
rect 222028 301580 222056 303826
rect 222212 301594 222240 338710
rect 222292 334688 222344 334694
rect 222292 334630 222344 334636
rect 222304 328545 222332 334630
rect 222290 328536 222346 328545
rect 222290 328471 222346 328480
rect 222304 325694 222332 328471
rect 224236 327049 224264 343023
rect 223578 327040 223634 327049
rect 223578 326975 223634 326984
rect 224222 327040 224278 327049
rect 224222 326975 224278 326984
rect 223592 325825 223620 326975
rect 223578 325816 223634 325825
rect 223578 325751 223634 325760
rect 223592 325694 223620 325751
rect 222304 325666 222792 325694
rect 223592 325666 224080 325694
rect 222764 301594 222792 325666
rect 223854 304328 223910 304337
rect 223854 304263 223910 304272
rect 222212 301566 222594 301594
rect 222764 301566 223238 301594
rect 223762 301200 223818 301209
rect 223868 301186 223896 304263
rect 224052 301594 224080 325666
rect 224224 314764 224276 314770
rect 224224 314706 224276 314712
rect 224236 305726 224264 314706
rect 224880 309806 224908 386242
rect 224972 385665 225000 386271
rect 224958 385656 225014 385665
rect 224958 385591 225014 385600
rect 225602 363624 225658 363633
rect 225602 363559 225658 363568
rect 225616 342961 225644 363559
rect 226352 362914 226380 390374
rect 227640 384402 227668 390388
rect 227732 390374 228574 390402
rect 226432 384396 226484 384402
rect 226432 384338 226484 384344
rect 227628 384396 227680 384402
rect 227628 384338 227680 384344
rect 226444 380254 226472 384338
rect 227640 383722 227668 384338
rect 227628 383716 227680 383722
rect 227628 383658 227680 383664
rect 227628 381540 227680 381546
rect 227628 381482 227680 381488
rect 226432 380248 226484 380254
rect 226432 380190 226484 380196
rect 226340 362908 226392 362914
rect 226340 362850 226392 362856
rect 226352 361622 226380 362850
rect 226340 361616 226392 361622
rect 226340 361558 226392 361564
rect 226984 361616 227036 361622
rect 226984 361558 227036 361564
rect 226996 351801 227024 361558
rect 226982 351792 227038 351801
rect 226982 351727 227038 351736
rect 225602 342952 225658 342961
rect 225602 342887 225658 342896
rect 226982 339552 227038 339561
rect 226982 339487 227038 339496
rect 224958 337376 225014 337385
rect 224958 337311 225014 337320
rect 225142 337376 225198 337385
rect 225142 337311 225198 337320
rect 224868 309800 224920 309806
rect 224868 309742 224920 309748
rect 224224 305720 224276 305726
rect 224224 305662 224276 305668
rect 224972 303686 225000 337311
rect 225156 335481 225184 337311
rect 225142 335472 225198 335481
rect 225142 335407 225198 335416
rect 225156 335354 225184 335407
rect 225064 335326 225184 335354
rect 224960 303680 225012 303686
rect 224960 303622 225012 303628
rect 224052 301566 224434 301594
rect 225064 301580 225092 335326
rect 225878 311264 225934 311273
rect 225878 311199 225934 311208
rect 225236 303680 225288 303686
rect 225236 303622 225288 303628
rect 225248 301594 225276 303622
rect 225892 301594 225920 311199
rect 226430 309496 226486 309505
rect 226430 309431 226486 309440
rect 226444 301594 226472 309431
rect 226890 306640 226946 306649
rect 226890 306575 226946 306584
rect 226904 301753 226932 306575
rect 226996 303657 227024 339487
rect 227640 304774 227668 381482
rect 227732 368422 227760 390374
rect 229664 389337 229692 390388
rect 229650 389328 229706 389337
rect 230584 389298 230612 390388
rect 230768 390374 231518 390402
rect 231872 390374 232438 390402
rect 229650 389263 229706 389272
rect 230572 389292 230624 389298
rect 230572 389234 230624 389240
rect 230584 387818 230612 389234
rect 230492 387790 230612 387818
rect 228364 387116 228416 387122
rect 228364 387058 228416 387064
rect 227810 381576 227866 381585
rect 227810 381511 227866 381520
rect 227824 378146 227852 381511
rect 227812 378140 227864 378146
rect 227812 378082 227864 378088
rect 228376 378078 228404 387058
rect 228364 378072 228416 378078
rect 228364 378014 228416 378020
rect 228454 377360 228510 377369
rect 228454 377295 228510 377304
rect 227720 368416 227772 368422
rect 227720 368358 227772 368364
rect 228364 367804 228416 367810
rect 228364 367746 228416 367752
rect 228376 316034 228404 367746
rect 228468 343738 228496 377295
rect 229742 369200 229798 369209
rect 229742 369135 229798 369144
rect 228548 368416 228600 368422
rect 228548 368358 228600 368364
rect 228560 362273 228588 368358
rect 228546 362264 228602 362273
rect 228546 362199 228602 362208
rect 228456 343732 228508 343738
rect 228456 343674 228508 343680
rect 228284 316006 228404 316034
rect 228284 311953 228312 316006
rect 228270 311944 228326 311953
rect 228270 311879 228326 311888
rect 227628 304768 227680 304774
rect 227628 304710 227680 304716
rect 227640 304201 227668 304710
rect 227626 304192 227682 304201
rect 227626 304127 227682 304136
rect 226982 303648 227038 303657
rect 226982 303583 227038 303592
rect 227994 303648 228050 303657
rect 227994 303583 228050 303592
rect 227444 302252 227496 302258
rect 227444 302194 227496 302200
rect 226890 301744 226946 301753
rect 226890 301679 226946 301688
rect 225248 301566 225630 301594
rect 225892 301566 226274 301594
rect 226444 301566 226826 301594
rect 227456 301580 227484 302194
rect 228008 301580 228036 303583
rect 228284 301594 228312 311879
rect 228468 302190 228496 343674
rect 229282 332616 229338 332625
rect 229282 332551 229338 332560
rect 229296 325694 229324 332551
rect 229296 325666 229416 325694
rect 229192 304768 229244 304774
rect 229192 304710 229244 304716
rect 228456 302184 228508 302190
rect 228456 302126 228508 302132
rect 228284 301566 228666 301594
rect 229204 301580 229232 304710
rect 229388 301594 229416 325666
rect 229756 308145 229784 369135
rect 230386 333296 230442 333305
rect 230386 333231 230442 333240
rect 230400 332625 230428 333231
rect 230386 332616 230442 332625
rect 230386 332551 230442 332560
rect 230492 308446 230520 387790
rect 230768 383654 230796 390374
rect 231216 387932 231268 387938
rect 231216 387874 231268 387880
rect 230768 383626 231164 383654
rect 231136 380934 231164 383626
rect 231124 380928 231176 380934
rect 231124 380870 231176 380876
rect 231136 349110 231164 380870
rect 231228 371210 231256 387874
rect 231872 382974 231900 390374
rect 232596 388000 232648 388006
rect 232596 387942 232648 387948
rect 232608 387569 232636 387942
rect 233344 387870 233372 390388
rect 234264 387938 234292 390388
rect 234252 387932 234304 387938
rect 234252 387874 234304 387880
rect 233332 387864 233384 387870
rect 233332 387806 233384 387812
rect 235264 387864 235316 387870
rect 235264 387806 235316 387812
rect 232594 387560 232650 387569
rect 232594 387495 232650 387504
rect 231860 382968 231912 382974
rect 231860 382910 231912 382916
rect 231216 371204 231268 371210
rect 231216 371146 231268 371152
rect 231228 360874 231256 371146
rect 232504 370524 232556 370530
rect 232504 370466 232556 370472
rect 231216 360868 231268 360874
rect 231216 360810 231268 360816
rect 231124 349104 231176 349110
rect 231124 349046 231176 349052
rect 231124 345092 231176 345098
rect 231124 345034 231176 345040
rect 230570 316840 230626 316849
rect 230570 316775 230626 316784
rect 230480 308440 230532 308446
rect 230480 308382 230532 308388
rect 229742 308136 229798 308145
rect 229742 308071 229798 308080
rect 229756 306374 229784 308071
rect 230584 306374 230612 316775
rect 231136 315314 231164 345034
rect 231124 315308 231176 315314
rect 231124 315250 231176 315256
rect 229756 306346 229968 306374
rect 230584 306346 231256 306374
rect 229940 301594 229968 306346
rect 230388 305652 230440 305658
rect 230388 305594 230440 305600
rect 230400 304366 230428 305594
rect 230388 304360 230440 304366
rect 230388 304302 230440 304308
rect 231032 302184 231084 302190
rect 231032 302126 231084 302132
rect 229388 301566 229862 301594
rect 229940 301566 230414 301594
rect 231044 301580 231072 302126
rect 231228 301594 231256 306346
rect 232228 303680 232280 303686
rect 232228 303622 232280 303628
rect 231228 301566 231610 301594
rect 232240 301580 232268 303622
rect 232516 302938 232544 370466
rect 232608 324970 232636 387495
rect 235276 379506 235304 387806
rect 235368 384441 235396 390388
rect 236288 388006 236316 390388
rect 236380 390374 237222 390402
rect 236276 388000 236328 388006
rect 236276 387942 236328 387948
rect 235354 384432 235410 384441
rect 235354 384367 235410 384376
rect 236380 380866 236408 390374
rect 238128 387802 238156 390388
rect 238116 387796 238168 387802
rect 238116 387738 238168 387744
rect 236368 380860 236420 380866
rect 236368 380802 236420 380808
rect 236644 380860 236696 380866
rect 236644 380802 236696 380808
rect 235264 379500 235316 379506
rect 235264 379442 235316 379448
rect 235908 379500 235960 379506
rect 235908 379442 235960 379448
rect 234528 371884 234580 371890
rect 234528 371826 234580 371832
rect 233884 329860 233936 329866
rect 233884 329802 233936 329808
rect 232596 324964 232648 324970
rect 232596 324906 232648 324912
rect 233608 322312 233660 322318
rect 233608 322254 233660 322260
rect 233146 312080 233202 312089
rect 233146 312015 233202 312024
rect 232780 304292 232832 304298
rect 232780 304234 232832 304240
rect 232504 302932 232556 302938
rect 232504 302874 232556 302880
rect 232792 301580 232820 304234
rect 233160 303686 233188 312015
rect 233422 309088 233478 309097
rect 233422 309023 233478 309032
rect 233436 308009 233464 309023
rect 233422 308000 233478 308009
rect 233422 307935 233478 307944
rect 233148 303680 233200 303686
rect 233148 303622 233200 303628
rect 233436 301580 233464 307935
rect 233620 301594 233648 322254
rect 233896 303686 233924 329802
rect 234540 325145 234568 371826
rect 234620 332580 234672 332586
rect 234620 332522 234672 332528
rect 234632 331294 234660 332522
rect 234620 331288 234672 331294
rect 234620 331230 234672 331236
rect 234632 325694 234660 331230
rect 234632 325666 235488 325694
rect 234526 325136 234582 325145
rect 234526 325071 234582 325080
rect 234540 324442 234568 325071
rect 234540 324414 234660 324442
rect 233974 318064 234030 318073
rect 233974 317999 234030 318008
rect 233988 309097 234016 317999
rect 234632 316034 234660 324414
rect 234632 316006 234752 316034
rect 233974 309088 234030 309097
rect 233974 309023 234030 309032
rect 233884 303680 233936 303686
rect 233884 303622 233936 303628
rect 234620 303680 234672 303686
rect 234620 303622 234672 303628
rect 233620 301566 234002 301594
rect 234632 301580 234660 303622
rect 234724 301594 234752 316006
rect 235460 301594 235488 325666
rect 235920 307086 235948 379442
rect 236656 369850 236684 380802
rect 236644 369844 236696 369850
rect 236644 369786 236696 369792
rect 236656 354006 236684 369786
rect 238022 356824 238078 356833
rect 238022 356759 238078 356768
rect 236644 354000 236696 354006
rect 236644 353942 236696 353948
rect 237286 314120 237342 314129
rect 237286 314055 237342 314064
rect 235998 313984 236054 313993
rect 235998 313919 236054 313928
rect 235908 307080 235960 307086
rect 235908 307022 235960 307028
rect 236012 301594 236040 313919
rect 234724 301566 235198 301594
rect 235460 301566 235842 301594
rect 236012 301566 236394 301594
rect 223818 301172 223896 301186
rect 223818 301158 223882 301172
rect 223762 301135 223818 301144
rect 196034 300886 196664 300914
rect 197636 300960 197688 300966
rect 236734 300928 236790 300937
rect 197688 300908 198030 300914
rect 197636 300902 198030 300908
rect 197648 300886 198030 300902
rect 195978 300863 196034 300872
rect 237300 300914 237328 314055
rect 238036 304337 238064 356759
rect 238128 353326 238156 387738
rect 239048 384305 239076 390388
rect 239416 390374 239982 390402
rect 239416 385014 239444 390374
rect 240782 389872 240838 389881
rect 240782 389807 240838 389816
rect 240140 389224 240192 389230
rect 240140 389166 240192 389172
rect 239404 385008 239456 385014
rect 239404 384950 239456 384956
rect 239034 384296 239090 384305
rect 239034 384231 239090 384240
rect 239416 356114 239444 384950
rect 240152 362302 240180 389166
rect 240140 362296 240192 362302
rect 240140 362238 240192 362244
rect 240140 359508 240192 359514
rect 240140 359450 240192 359456
rect 240046 359136 240102 359145
rect 240046 359071 240102 359080
rect 239404 356108 239456 356114
rect 239404 356050 239456 356056
rect 238116 353320 238168 353326
rect 238116 353262 238168 353268
rect 238128 330585 238156 353262
rect 239416 339454 239444 356050
rect 239404 339448 239456 339454
rect 239404 339390 239456 339396
rect 238114 330576 238170 330585
rect 238114 330511 238170 330520
rect 238666 313984 238722 313993
rect 238666 313919 238722 313928
rect 238022 304328 238078 304337
rect 238022 304263 238078 304272
rect 238206 302424 238262 302433
rect 238206 302359 238262 302368
rect 238220 301580 238248 302359
rect 238680 300966 238708 313919
rect 239404 303680 239456 303686
rect 239404 303622 239456 303628
rect 239126 302832 239182 302841
rect 239126 302767 239182 302776
rect 239140 301594 239168 302767
rect 238878 301566 239168 301594
rect 239416 301580 239444 303622
rect 240060 302258 240088 359071
rect 240152 328574 240180 359450
rect 240796 332586 240824 389807
rect 241072 389230 241100 390388
rect 241532 390374 242006 390402
rect 241532 389230 241560 390374
rect 241060 389224 241112 389230
rect 241060 389166 241112 389172
rect 241520 389224 241572 389230
rect 241520 389166 241572 389172
rect 241428 378820 241480 378826
rect 241428 378762 241480 378768
rect 240784 332580 240836 332586
rect 240784 332522 240836 332528
rect 240140 328568 240192 328574
rect 240140 328510 240192 328516
rect 240152 325694 240180 328510
rect 240152 325666 240732 325694
rect 240600 302320 240652 302326
rect 240600 302262 240652 302268
rect 240048 302252 240100 302258
rect 240048 302194 240100 302200
rect 240060 301580 240088 302194
rect 240612 301580 240640 302262
rect 240704 301594 240732 325666
rect 240784 313404 240836 313410
rect 240784 313346 240836 313352
rect 240796 305833 240824 313346
rect 240782 305824 240838 305833
rect 240782 305759 240838 305768
rect 241440 302326 241468 378762
rect 241532 364410 241560 389166
rect 242912 388657 242940 390388
rect 243096 390374 243846 390402
rect 242898 388648 242954 388657
rect 242898 388583 242954 388592
rect 242912 386209 242940 388583
rect 242898 386200 242954 386209
rect 242898 386135 242954 386144
rect 243096 379409 243124 390374
rect 244752 389065 244780 390388
rect 244738 389056 244794 389065
rect 244738 388991 244794 389000
rect 244370 384432 244426 384441
rect 244370 384367 244426 384376
rect 244278 383072 244334 383081
rect 244278 383007 244334 383016
rect 243082 379400 243138 379409
rect 243082 379335 243138 379344
rect 243096 378078 243124 379335
rect 243084 378072 243136 378078
rect 243084 378014 243136 378020
rect 242348 373312 242400 373318
rect 242348 373254 242400 373260
rect 241520 364404 241572 364410
rect 241520 364346 241572 364352
rect 242254 362264 242310 362273
rect 242254 362199 242310 362208
rect 242164 356720 242216 356726
rect 242164 356662 242216 356668
rect 241520 326392 241572 326398
rect 241520 326334 241572 326340
rect 241428 302320 241480 302326
rect 241428 302262 241480 302268
rect 241532 301594 241560 326334
rect 242176 305697 242204 356662
rect 242268 326398 242296 362199
rect 242360 347070 242388 373254
rect 242348 347064 242400 347070
rect 242348 347006 242400 347012
rect 243544 338836 243596 338842
rect 243544 338778 243596 338784
rect 242900 334620 242952 334626
rect 242900 334562 242952 334568
rect 242256 326392 242308 326398
rect 242256 326334 242308 326340
rect 242808 307828 242860 307834
rect 242808 307770 242860 307776
rect 242162 305688 242218 305697
rect 242162 305623 242218 305632
rect 242440 305652 242492 305658
rect 242440 305594 242492 305600
rect 240704 301566 241270 301594
rect 241532 301566 241822 301594
rect 242452 301580 242480 305594
rect 242820 303686 242848 307770
rect 242912 303686 242940 334562
rect 243176 331900 243228 331906
rect 243176 331842 243228 331848
rect 242990 303784 243046 303793
rect 242990 303719 243046 303728
rect 242808 303680 242860 303686
rect 242808 303622 242860 303628
rect 242900 303680 242952 303686
rect 242900 303622 242952 303628
rect 243004 301580 243032 303719
rect 243188 301594 243216 331842
rect 243556 303793 243584 338778
rect 244292 335850 244320 383007
rect 244384 366897 244412 384367
rect 245672 373969 245700 390388
rect 245764 390374 246606 390402
rect 245764 375426 245792 390374
rect 247696 384985 247724 390388
rect 248616 389065 248644 390918
rect 251732 390934 251784 390940
rect 252558 390960 252614 390969
rect 248878 390895 248934 390904
rect 250718 390824 250774 390833
rect 250718 390759 250774 390768
rect 249536 389065 249564 390388
rect 250456 389162 250484 390388
rect 250444 389156 250496 389162
rect 250444 389098 250496 389104
rect 247774 389056 247830 389065
rect 247774 388991 247830 389000
rect 248602 389056 248658 389065
rect 248602 388991 248658 389000
rect 249246 389056 249302 389065
rect 249246 388991 249302 389000
rect 249522 389056 249578 389065
rect 249522 388991 249578 389000
rect 247682 384976 247738 384985
rect 247682 384911 247738 384920
rect 247696 380905 247724 384911
rect 247682 380896 247738 380905
rect 247682 380831 247738 380840
rect 245752 375420 245804 375426
rect 245752 375362 245804 375368
rect 245658 373960 245714 373969
rect 245658 373895 245714 373904
rect 245672 372745 245700 373895
rect 245658 372736 245714 372745
rect 245658 372671 245714 372680
rect 246302 372736 246358 372745
rect 246302 372671 246358 372680
rect 244370 366888 244426 366897
rect 244370 366823 244426 366832
rect 244924 355360 244976 355366
rect 244924 355302 244976 355308
rect 244280 335844 244332 335850
rect 244280 335786 244332 335792
rect 244292 335374 244320 335786
rect 244280 335368 244332 335374
rect 244280 335310 244332 335316
rect 244830 311944 244886 311953
rect 244830 311879 244886 311888
rect 244740 304088 244792 304094
rect 244740 304030 244792 304036
rect 243542 303784 243598 303793
rect 243542 303719 243598 303728
rect 243820 303680 243872 303686
rect 243820 303622 243872 303628
rect 243832 301594 243860 303622
rect 244752 301594 244780 304030
rect 244844 301730 244872 311879
rect 244936 303657 244964 355302
rect 246316 347041 246344 372671
rect 246394 362264 246450 362273
rect 246394 362199 246450 362208
rect 246302 347032 246358 347041
rect 246302 346967 246358 346976
rect 246408 343097 246436 362199
rect 247696 344350 247724 380831
rect 247788 362234 247816 388991
rect 249156 387864 249208 387870
rect 249156 387806 249208 387812
rect 249064 364404 249116 364410
rect 249064 364346 249116 364352
rect 247776 362228 247828 362234
rect 247776 362170 247828 362176
rect 247776 358080 247828 358086
rect 247776 358022 247828 358028
rect 247684 344344 247736 344350
rect 247684 344286 247736 344292
rect 246488 343664 246540 343670
rect 246488 343606 246540 343612
rect 246394 343088 246450 343097
rect 246394 343023 246450 343032
rect 246396 340196 246448 340202
rect 246396 340138 246448 340144
rect 246304 339448 246356 339454
rect 246304 339390 246356 339396
rect 245016 335844 245068 335850
rect 245016 335786 245068 335792
rect 245028 311953 245056 335786
rect 245752 333328 245804 333334
rect 245752 333270 245804 333276
rect 245014 311944 245070 311953
rect 245014 311879 245070 311888
rect 244922 303648 244978 303657
rect 244922 303583 244978 303592
rect 244844 301702 245056 301730
rect 245028 301594 245056 301702
rect 245764 301594 245792 333270
rect 246316 304706 246344 339390
rect 246408 307193 246436 340138
rect 246500 333334 246528 343606
rect 246948 338768 247000 338774
rect 246948 338710 247000 338716
rect 246488 333328 246540 333334
rect 246488 333270 246540 333276
rect 246394 307184 246450 307193
rect 246394 307119 246450 307128
rect 246960 305017 246988 338710
rect 247788 336802 247816 358022
rect 247776 336796 247828 336802
rect 247776 336738 247828 336744
rect 247788 335354 247816 336738
rect 247696 335326 247816 335354
rect 247040 333260 247092 333266
rect 247040 333202 247092 333208
rect 246946 305008 247002 305017
rect 246946 304943 247002 304952
rect 246304 304700 246356 304706
rect 246304 304642 246356 304648
rect 246580 304360 246632 304366
rect 246580 304302 246632 304308
rect 243188 301566 243662 301594
rect 243832 301566 244214 301594
rect 244752 301566 244858 301594
rect 245028 301566 245410 301594
rect 245764 301566 246054 301594
rect 246592 301580 246620 304302
rect 246960 304094 246988 304943
rect 246948 304088 247000 304094
rect 246948 304030 247000 304036
rect 247052 301594 247080 333202
rect 247130 325816 247186 325825
rect 247130 325751 247186 325760
rect 247144 320142 247172 325751
rect 247132 320136 247184 320142
rect 247132 320078 247184 320084
rect 247696 308009 247724 335326
rect 247682 308000 247738 308009
rect 247682 307935 247738 307944
rect 247696 301594 247724 307935
rect 249076 304201 249104 364346
rect 249168 361554 249196 387806
rect 249260 371929 249288 388991
rect 250456 373998 250484 389098
rect 250444 373992 250496 373998
rect 250732 373994 250760 390759
rect 251284 390374 251390 390402
rect 251284 376718 251312 390374
rect 251744 385014 251772 390934
rect 252558 390895 252614 390904
rect 252296 387870 252324 390388
rect 252284 387864 252336 387870
rect 252284 387806 252336 387812
rect 252572 386374 252600 390895
rect 253400 389094 253428 390388
rect 253388 389088 253440 389094
rect 253388 389030 253440 389036
rect 253400 387122 253428 389030
rect 253388 387116 253440 387122
rect 253388 387058 253440 387064
rect 252560 386368 252612 386374
rect 252560 386310 252612 386316
rect 251732 385008 251784 385014
rect 251732 384950 251784 384956
rect 251824 385008 251876 385014
rect 251824 384950 251876 384956
rect 251272 376712 251324 376718
rect 251272 376654 251324 376660
rect 250444 373934 250496 373940
rect 250548 373966 250760 373994
rect 249246 371920 249302 371929
rect 249246 371855 249302 371864
rect 249614 371920 249670 371929
rect 249614 371855 249670 371864
rect 249628 364993 249656 371855
rect 249708 365152 249760 365158
rect 249708 365094 249760 365100
rect 249614 364984 249670 364993
rect 249614 364919 249670 364928
rect 249156 361548 249208 361554
rect 249156 361490 249208 361496
rect 249616 361548 249668 361554
rect 249616 361490 249668 361496
rect 249628 355366 249656 361490
rect 249616 355360 249668 355366
rect 249616 355302 249668 355308
rect 249156 317552 249208 317558
rect 249156 317494 249208 317500
rect 249168 304298 249196 317494
rect 249614 311264 249670 311273
rect 249614 311199 249670 311208
rect 249156 304292 249208 304298
rect 249156 304234 249208 304240
rect 249062 304192 249118 304201
rect 249062 304127 249118 304136
rect 249628 303686 249656 311199
rect 248420 303680 248472 303686
rect 248420 303622 248472 303628
rect 249616 303680 249668 303686
rect 249616 303622 249668 303628
rect 247052 301566 247250 301594
rect 247696 301566 247802 301594
rect 248432 301580 248460 303622
rect 249720 302433 249748 365094
rect 250444 325712 250496 325718
rect 250548 325694 250576 373966
rect 251836 361593 251864 384950
rect 252468 383036 252520 383042
rect 252468 382978 252520 382984
rect 251822 361584 251878 361593
rect 251822 361519 251878 361528
rect 250496 325666 250576 325694
rect 250444 325654 250496 325660
rect 250168 304700 250220 304706
rect 250168 304642 250220 304648
rect 248970 302424 249026 302433
rect 248970 302359 249026 302368
rect 249706 302424 249762 302433
rect 249706 302359 249762 302368
rect 248984 301580 249012 302359
rect 250180 301580 250208 304642
rect 250456 301578 250484 325654
rect 251836 309369 251864 361519
rect 251916 344344 251968 344350
rect 251916 344286 251968 344292
rect 251928 330721 251956 344286
rect 251914 330712 251970 330721
rect 251914 330647 251970 330656
rect 252376 329792 252428 329798
rect 252376 329734 252428 329740
rect 252388 328506 252416 329734
rect 252376 328500 252428 328506
rect 252376 328442 252428 328448
rect 252284 319456 252336 319462
rect 252284 319398 252336 319404
rect 251916 310548 251968 310554
rect 251916 310490 251968 310496
rect 251822 309360 251878 309369
rect 251822 309295 251878 309304
rect 251362 306504 251418 306513
rect 251362 306439 251418 306448
rect 250810 303784 250866 303793
rect 250810 303719 250866 303728
rect 250824 303686 250852 303719
rect 250812 303680 250864 303686
rect 250812 303622 250864 303628
rect 250824 301580 250852 303622
rect 251376 301580 251404 306439
rect 251836 301594 251864 309295
rect 251928 307057 251956 310490
rect 251914 307048 251970 307057
rect 251914 306983 251970 306992
rect 252296 306921 252324 319398
rect 252282 306912 252338 306921
rect 252282 306847 252338 306856
rect 252296 302297 252324 306847
rect 252282 302288 252338 302297
rect 252282 302223 252338 302232
rect 250444 301572 250496 301578
rect 251836 301566 252034 301594
rect 250444 301514 250496 301520
rect 236790 300886 237328 300914
rect 237380 300960 237432 300966
rect 238668 300960 238720 300966
rect 237432 300908 237590 300914
rect 237380 300902 237590 300908
rect 249706 300928 249762 300937
rect 238668 300902 238720 300908
rect 237392 300886 237590 300902
rect 249642 300886 249706 300914
rect 236734 300863 236790 300872
rect 252388 300898 252416 328442
rect 252480 311273 252508 382978
rect 252572 365158 252600 386310
rect 252560 365152 252612 365158
rect 252560 365094 252612 365100
rect 253204 360868 253256 360874
rect 253204 360810 253256 360816
rect 252836 352640 252888 352646
rect 252836 352582 252888 352588
rect 252848 325694 252876 352582
rect 253216 334665 253244 360810
rect 253492 348430 253520 393286
rect 253952 378826 253980 448582
rect 254044 392873 254072 458798
rect 254136 427938 254164 479470
rect 254216 456068 254268 456074
rect 254216 456010 254268 456016
rect 254228 432041 254256 456010
rect 254214 432032 254270 432041
rect 254214 431967 254216 431976
rect 254268 431967 254270 431976
rect 254216 431938 254268 431944
rect 254214 427952 254270 427961
rect 254136 427910 254214 427938
rect 254214 427887 254270 427896
rect 254122 415168 254178 415177
rect 254122 415103 254178 415112
rect 254030 392864 254086 392873
rect 254030 392799 254086 392808
rect 254044 392154 254072 392799
rect 254032 392148 254084 392154
rect 254032 392090 254084 392096
rect 254030 392048 254086 392057
rect 254030 391983 254086 391992
rect 254044 385014 254072 391983
rect 254136 388226 254164 415103
rect 254228 388521 254256 427887
rect 255332 415177 255360 584038
rect 255412 583704 255464 583710
rect 255412 583646 255464 583652
rect 255424 583273 255452 583646
rect 255410 583264 255466 583273
rect 255410 583199 255466 583208
rect 255976 580310 256004 598839
rect 256068 587178 256096 598878
rect 256330 592784 256386 592793
rect 256330 592719 256386 592728
rect 256344 592686 256372 592719
rect 256712 592686 256740 609962
rect 257344 599072 257396 599078
rect 257344 599014 257396 599020
rect 256332 592680 256384 592686
rect 256332 592622 256384 592628
rect 256700 592680 256752 592686
rect 256700 592622 256752 592628
rect 256056 587172 256108 587178
rect 256056 587114 256108 587120
rect 255964 580304 256016 580310
rect 255964 580246 256016 580252
rect 255410 579728 255466 579737
rect 255410 579663 255466 579672
rect 255424 577522 255452 579663
rect 255412 577516 255464 577522
rect 255412 577458 255464 577464
rect 255410 577008 255466 577017
rect 255410 576943 255466 576952
rect 255424 576910 255452 576943
rect 255412 576904 255464 576910
rect 255412 576846 255464 576852
rect 255410 575920 255466 575929
rect 255410 575855 255466 575864
rect 255424 575550 255452 575855
rect 255412 575544 255464 575550
rect 255412 575486 255464 575492
rect 255410 574696 255466 574705
rect 255410 574631 255466 574640
rect 255424 574122 255452 574631
rect 255594 574152 255650 574161
rect 255412 574116 255464 574122
rect 255594 574087 255650 574096
rect 255412 574058 255464 574064
rect 255502 572928 255558 572937
rect 255502 572863 255558 572872
rect 255412 572756 255464 572762
rect 255412 572698 255464 572704
rect 255424 572665 255452 572698
rect 255410 572656 255466 572665
rect 255410 572591 255466 572600
rect 255410 571568 255466 571577
rect 255410 571503 255466 571512
rect 255424 571402 255452 571503
rect 255412 571396 255464 571402
rect 255412 571338 255464 571344
rect 255412 570648 255464 570654
rect 255410 570616 255412 570625
rect 255464 570616 255466 570625
rect 255410 570551 255466 570560
rect 255410 569392 255466 569401
rect 255410 569327 255466 569336
rect 255424 568954 255452 569327
rect 255412 568948 255464 568954
rect 255412 568890 255464 568896
rect 255410 568712 255466 568721
rect 255410 568647 255466 568656
rect 255424 568614 255452 568647
rect 255412 568608 255464 568614
rect 255412 568550 255464 568556
rect 255516 567866 255544 572863
rect 255504 567860 255556 567866
rect 255504 567802 255556 567808
rect 255608 567304 255636 574087
rect 255688 570648 255740 570654
rect 255688 570590 255740 570596
rect 255424 567276 255636 567304
rect 255424 431254 255452 567276
rect 255700 567194 255728 570590
rect 255778 567624 255834 567633
rect 255778 567559 255834 567568
rect 255792 567322 255820 567559
rect 255780 567316 255832 567322
rect 255780 567258 255832 567264
rect 255516 567166 255728 567194
rect 255516 537985 255544 567166
rect 255686 566400 255742 566409
rect 255686 566335 255742 566344
rect 255700 565962 255728 566335
rect 255688 565956 255740 565962
rect 255688 565898 255740 565904
rect 255596 565888 255648 565894
rect 255594 565856 255596 565865
rect 255648 565856 255650 565865
rect 255594 565791 255650 565800
rect 255594 564768 255650 564777
rect 255594 564703 255650 564712
rect 255608 564466 255636 564703
rect 255596 564460 255648 564466
rect 255596 564402 255648 564408
rect 255594 563136 255650 563145
rect 255594 563071 255596 563080
rect 255648 563071 255650 563080
rect 255596 563042 255648 563048
rect 255594 561912 255650 561921
rect 255594 561847 255650 561856
rect 255608 561746 255636 561847
rect 255596 561740 255648 561746
rect 255596 561682 255648 561688
rect 255594 560824 255650 560833
rect 255594 560759 255650 560768
rect 255608 560318 255636 560759
rect 255596 560312 255648 560318
rect 255596 560254 255648 560260
rect 255594 559600 255650 559609
rect 255594 559535 255650 559544
rect 255608 558958 255636 559535
rect 255596 558952 255648 558958
rect 255596 558894 255648 558900
rect 255594 557968 255650 557977
rect 255594 557903 255650 557912
rect 255608 557598 255636 557903
rect 255596 557592 255648 557598
rect 255596 557534 255648 557540
rect 255594 556880 255650 556889
rect 255594 556815 255650 556824
rect 255608 556238 255636 556815
rect 255596 556232 255648 556238
rect 255596 556174 255648 556180
rect 257356 555490 257384 599014
rect 258092 584458 258120 612750
rect 263692 601792 263744 601798
rect 263692 601734 263744 601740
rect 259460 601724 259512 601730
rect 259460 601666 259512 601672
rect 258080 584452 258132 584458
rect 258080 584394 258132 584400
rect 258080 568948 258132 568954
rect 258080 568890 258132 568896
rect 257344 555484 257396 555490
rect 257344 555426 257396 555432
rect 256606 554976 256662 554985
rect 256662 554934 256740 554962
rect 256606 554911 256662 554920
rect 255686 554160 255742 554169
rect 255686 554095 255742 554104
rect 255594 553616 255650 553625
rect 255594 553551 255650 553560
rect 255608 553518 255636 553551
rect 255596 553512 255648 553518
rect 255596 553454 255648 553460
rect 255700 553450 255728 554095
rect 255688 553444 255740 553450
rect 255688 553386 255740 553392
rect 255594 552800 255650 552809
rect 255594 552735 255650 552744
rect 255608 552702 255636 552735
rect 255596 552696 255648 552702
rect 255596 552638 255648 552644
rect 255594 550896 255650 550905
rect 255594 550831 255650 550840
rect 255608 550730 255636 550831
rect 255596 550724 255648 550730
rect 255596 550666 255648 550672
rect 255596 550588 255648 550594
rect 255596 550530 255648 550536
rect 255608 550225 255636 550530
rect 255594 550216 255650 550225
rect 255594 550151 255650 550160
rect 255594 548448 255650 548457
rect 255594 548383 255650 548392
rect 255608 547942 255636 548383
rect 255596 547936 255648 547942
rect 255596 547878 255648 547884
rect 255594 546816 255650 546825
rect 255594 546751 255650 546760
rect 255608 546514 255636 546751
rect 255596 546508 255648 546514
rect 255596 546450 255648 546456
rect 255594 545864 255650 545873
rect 255594 545799 255650 545808
rect 255608 545290 255636 545799
rect 255596 545284 255648 545290
rect 255596 545226 255648 545232
rect 255686 545184 255742 545193
rect 255686 545119 255742 545128
rect 255594 544096 255650 544105
rect 255594 544031 255650 544040
rect 255608 543794 255636 544031
rect 255596 543788 255648 543794
rect 255596 543730 255648 543736
rect 255594 541240 255650 541249
rect 255594 541175 255650 541184
rect 255608 541006 255636 541175
rect 255596 541000 255648 541006
rect 255596 540942 255648 540948
rect 255700 539374 255728 545119
rect 255688 539368 255740 539374
rect 255688 539310 255740 539316
rect 255594 538928 255650 538937
rect 255594 538863 255650 538872
rect 255608 538286 255636 538863
rect 255596 538280 255648 538286
rect 255596 538222 255648 538228
rect 255502 537976 255558 537985
rect 255502 537911 255558 537920
rect 255516 467158 255544 537911
rect 256712 530602 256740 554934
rect 256790 551168 256846 551177
rect 256790 551103 256846 551112
rect 256804 531321 256832 551103
rect 257066 533352 257122 533361
rect 257066 533287 257122 533296
rect 256790 531312 256846 531321
rect 256790 531247 256846 531256
rect 256700 530596 256752 530602
rect 256700 530538 256752 530544
rect 256792 494828 256844 494834
rect 256792 494770 256844 494776
rect 255504 467152 255556 467158
rect 255504 467094 255556 467100
rect 255516 466721 255544 467094
rect 255502 466712 255558 466721
rect 255502 466647 255558 466656
rect 255502 465760 255558 465769
rect 255502 465695 255558 465704
rect 255516 444825 255544 465695
rect 255594 460320 255650 460329
rect 255594 460255 255650 460264
rect 255608 448905 255636 460255
rect 255594 448896 255650 448905
rect 255594 448831 255650 448840
rect 255608 447817 255636 448831
rect 255594 447808 255650 447817
rect 255594 447743 255650 447752
rect 255594 447536 255650 447545
rect 255594 447471 255650 447480
rect 255608 446418 255636 447471
rect 255596 446412 255648 446418
rect 255596 446354 255648 446360
rect 255962 446176 256018 446185
rect 255962 446111 256018 446120
rect 255502 444816 255558 444825
rect 255502 444751 255558 444760
rect 255504 443896 255556 443902
rect 255504 443838 255556 443844
rect 255516 443465 255544 443838
rect 255502 443456 255558 443465
rect 255502 443391 255558 443400
rect 255504 442264 255556 442270
rect 255504 442206 255556 442212
rect 255516 442105 255544 442206
rect 255502 442096 255558 442105
rect 255502 442031 255558 442040
rect 255504 439544 255556 439550
rect 255504 439486 255556 439492
rect 255516 439113 255544 439486
rect 255502 439104 255558 439113
rect 255502 439039 255558 439048
rect 255504 438864 255556 438870
rect 255504 438806 255556 438812
rect 255516 437753 255544 438806
rect 255976 438802 256004 446111
rect 255964 438796 256016 438802
rect 255964 438738 256016 438744
rect 255502 437744 255558 437753
rect 255502 437679 255558 437688
rect 255870 437608 255926 437617
rect 255870 437543 255926 437552
rect 255884 436393 255912 437543
rect 255870 436384 255926 436393
rect 255870 436319 255926 436328
rect 255504 436076 255556 436082
rect 255504 436018 255556 436024
rect 255516 435033 255544 436018
rect 255502 435024 255558 435033
rect 255502 434959 255558 434968
rect 255504 434036 255556 434042
rect 255504 433978 255556 433984
rect 255516 433673 255544 433978
rect 255502 433664 255558 433673
rect 255502 433599 255558 433608
rect 255412 431248 255464 431254
rect 255412 431190 255464 431196
rect 255424 430681 255452 431190
rect 255410 430672 255466 430681
rect 255410 430607 255466 430616
rect 255412 429548 255464 429554
rect 255412 429490 255464 429496
rect 255424 429321 255452 429490
rect 255410 429312 255466 429321
rect 255410 429247 255466 429256
rect 255410 426592 255466 426601
rect 255410 426527 255466 426536
rect 255424 426494 255452 426527
rect 255412 426488 255464 426494
rect 255412 426430 255464 426436
rect 256608 425740 256660 425746
rect 256608 425682 256660 425688
rect 256620 425241 256648 425682
rect 256606 425232 256662 425241
rect 256606 425167 256662 425176
rect 256620 424386 256648 425167
rect 256608 424380 256660 424386
rect 256608 424322 256660 424328
rect 255502 423600 255558 423609
rect 255502 423535 255558 423544
rect 255516 422346 255544 423535
rect 255504 422340 255556 422346
rect 255504 422282 255556 422288
rect 255502 422240 255558 422249
rect 255502 422175 255558 422184
rect 255516 420986 255544 422175
rect 255504 420980 255556 420986
rect 255504 420922 255556 420928
rect 255502 420880 255558 420889
rect 255502 420815 255558 420824
rect 255516 419558 255544 420815
rect 255504 419552 255556 419558
rect 255410 419520 255466 419529
rect 255504 419494 255556 419500
rect 255410 419455 255412 419464
rect 255464 419455 255466 419464
rect 255412 419426 255464 419432
rect 255502 418160 255558 418169
rect 255502 418095 255558 418104
rect 255516 416838 255544 418095
rect 255504 416832 255556 416838
rect 255410 416800 255466 416809
rect 255504 416774 255556 416780
rect 255410 416735 255412 416744
rect 255464 416735 255466 416744
rect 255412 416706 255464 416712
rect 255318 415168 255374 415177
rect 255318 415103 255374 415112
rect 255504 412616 255556 412622
rect 255504 412558 255556 412564
rect 255516 412457 255544 412558
rect 255502 412448 255558 412457
rect 255502 412383 255558 412392
rect 255502 411088 255558 411097
rect 255502 411023 255558 411032
rect 255410 409728 255466 409737
rect 255410 409663 255466 409672
rect 255424 408542 255452 409663
rect 255412 408536 255464 408542
rect 255412 408478 255464 408484
rect 255410 408368 255466 408377
rect 255410 408303 255466 408312
rect 255424 407862 255452 408303
rect 255412 407856 255464 407862
rect 255412 407798 255464 407804
rect 255424 406450 255452 407798
rect 255516 407794 255544 411023
rect 255504 407788 255556 407794
rect 255504 407730 255556 407736
rect 255502 407008 255558 407017
rect 255502 406943 255558 406952
rect 255332 406422 255452 406450
rect 254214 388512 254270 388521
rect 254214 388447 254270 388456
rect 254136 388198 254348 388226
rect 254214 388104 254270 388113
rect 254214 388039 254270 388048
rect 254032 385008 254084 385014
rect 254032 384950 254084 384956
rect 254228 384690 254256 388039
rect 254044 384662 254256 384690
rect 253940 378820 253992 378826
rect 253940 378762 253992 378768
rect 253938 375320 253994 375329
rect 253938 375255 253994 375264
rect 253952 358086 253980 375255
rect 253940 358080 253992 358086
rect 253940 358022 253992 358028
rect 253480 348424 253532 348430
rect 253480 348366 253532 348372
rect 253296 341624 253348 341630
rect 253296 341566 253348 341572
rect 253202 334656 253258 334665
rect 253202 334591 253258 334600
rect 253308 329225 253336 341566
rect 254044 329798 254072 384662
rect 254320 383738 254348 388198
rect 254136 383710 254348 383738
rect 254136 375329 254164 383710
rect 255332 383654 255360 406422
rect 255516 405754 255544 406943
rect 255504 405748 255556 405754
rect 255504 405690 255556 405696
rect 255410 404016 255466 404025
rect 255410 403951 255466 403960
rect 255424 403034 255452 403951
rect 255412 403028 255464 403034
rect 255412 402970 255464 402976
rect 255410 402656 255466 402665
rect 255410 402591 255466 402600
rect 255424 401674 255452 402591
rect 255412 401668 255464 401674
rect 255412 401610 255464 401616
rect 255410 401296 255466 401305
rect 255410 401231 255466 401240
rect 255424 400246 255452 401231
rect 255412 400240 255464 400246
rect 255412 400182 255464 400188
rect 255410 399936 255466 399945
rect 255410 399871 255466 399880
rect 255424 398138 255452 399871
rect 255412 398132 255464 398138
rect 255412 398074 255464 398080
rect 255410 395584 255466 395593
rect 255410 395519 255466 395528
rect 255424 394738 255452 395519
rect 255412 394732 255464 394738
rect 255412 394674 255464 394680
rect 255410 394224 255466 394233
rect 255410 394159 255466 394168
rect 255424 393378 255452 394159
rect 256700 393984 256752 393990
rect 256700 393926 256752 393932
rect 255412 393372 255464 393378
rect 255412 393314 255464 393320
rect 255504 392148 255556 392154
rect 255504 392090 255556 392096
rect 255332 383626 255452 383654
rect 254122 375320 254178 375329
rect 254122 375255 254178 375264
rect 255424 369782 255452 383626
rect 255412 369776 255464 369782
rect 255412 369718 255464 369724
rect 254584 349920 254636 349926
rect 254584 349862 254636 349868
rect 254032 329792 254084 329798
rect 254032 329734 254084 329740
rect 253294 329216 253350 329225
rect 253294 329151 253350 329160
rect 252848 325666 253336 325694
rect 252466 311264 252522 311273
rect 252466 311199 252522 311208
rect 252744 308440 252796 308446
rect 252744 308382 252796 308388
rect 252560 307080 252612 307086
rect 252560 307022 252612 307028
rect 249706 300863 249762 300872
rect 252376 300892 252428 300898
rect 252376 300834 252428 300840
rect 193734 295174 193812 295202
rect 193678 295151 193734 295160
rect 192482 291816 192538 291825
rect 192482 291751 192538 291760
rect 193128 284300 193180 284306
rect 193128 284242 193180 284248
rect 193140 283529 193168 284242
rect 193126 283520 193182 283529
rect 193126 283455 193182 283464
rect 191852 267706 192064 267734
rect 192036 263945 192064 267706
rect 192576 267028 192628 267034
rect 192576 266970 192628 266976
rect 192022 263936 192078 263945
rect 192022 263871 192078 263880
rect 192036 263634 192064 263871
rect 192024 263628 192076 263634
rect 192024 263570 192076 263576
rect 191668 248386 191788 248414
rect 191196 246356 191248 246362
rect 191196 246298 191248 246304
rect 191208 229022 191236 246298
rect 191668 244361 191696 248386
rect 191746 247616 191802 247625
rect 191746 247551 191802 247560
rect 191760 247110 191788 247551
rect 191748 247104 191800 247110
rect 191748 247046 191800 247052
rect 191286 244352 191342 244361
rect 191286 244287 191342 244296
rect 191654 244352 191710 244361
rect 191654 244287 191710 244296
rect 191300 235249 191328 244287
rect 192484 243568 192536 243574
rect 192484 243510 192536 243516
rect 191838 242856 191894 242865
rect 191838 242791 191894 242800
rect 191746 242176 191802 242185
rect 191746 242111 191802 242120
rect 191760 241602 191788 242111
rect 191852 241602 191880 242791
rect 191748 241596 191800 241602
rect 191748 241538 191800 241544
rect 191840 241596 191892 241602
rect 191840 241538 191892 241544
rect 191286 235240 191342 235249
rect 191286 235175 191342 235184
rect 191196 229016 191248 229022
rect 191196 228958 191248 228964
rect 191104 204264 191156 204270
rect 191104 204206 191156 204212
rect 190460 184204 190512 184210
rect 190460 184146 190512 184152
rect 190368 177336 190420 177342
rect 190368 177278 190420 177284
rect 189908 156052 189960 156058
rect 189908 155994 189960 156000
rect 189172 153876 189224 153882
rect 189172 153818 189224 153824
rect 189078 152416 189134 152425
rect 189078 152351 189134 152360
rect 189184 151094 189212 153818
rect 189172 151088 189224 151094
rect 189172 151030 189224 151036
rect 189184 150482 189212 151030
rect 189172 150476 189224 150482
rect 189172 150418 189224 150424
rect 189816 150476 189868 150482
rect 189816 150418 189868 150424
rect 189080 142248 189132 142254
rect 189080 142190 189132 142196
rect 189092 137290 189120 142190
rect 189080 137284 189132 137290
rect 189080 137226 189132 137232
rect 188988 135244 189040 135250
rect 188988 135186 189040 135192
rect 189724 135244 189776 135250
rect 189724 135186 189776 135192
rect 188896 134020 188948 134026
rect 188896 133962 188948 133968
rect 188804 124840 188856 124846
rect 188804 124782 188856 124788
rect 188344 122120 188396 122126
rect 188344 122062 188396 122068
rect 187700 117972 187752 117978
rect 187700 117914 187752 117920
rect 187712 117434 187740 117914
rect 187700 117428 187752 117434
rect 187700 117370 187752 117376
rect 188252 113280 188304 113286
rect 188252 113222 188304 113228
rect 188264 109750 188292 113222
rect 188252 109744 188304 109750
rect 188252 109686 188304 109692
rect 187608 107568 187660 107574
rect 187608 107510 187660 107516
rect 188356 105942 188384 122062
rect 188344 105936 188396 105942
rect 188344 105878 188396 105884
rect 188344 102808 188396 102814
rect 188344 102750 188396 102756
rect 188356 82822 188384 102750
rect 188436 96688 188488 96694
rect 188436 96630 188488 96636
rect 188448 92313 188476 96630
rect 188434 92304 188490 92313
rect 188434 92239 188490 92248
rect 188526 91216 188582 91225
rect 188526 91151 188582 91160
rect 188540 88262 188568 91151
rect 188528 88256 188580 88262
rect 188528 88198 188580 88204
rect 188344 82816 188396 82822
rect 188344 82758 188396 82764
rect 188908 65550 188936 133962
rect 188988 117428 189040 117434
rect 188988 117370 189040 117376
rect 188896 65544 188948 65550
rect 188896 65486 188948 65492
rect 187516 47592 187568 47598
rect 187516 47534 187568 47540
rect 189000 11762 189028 117370
rect 189080 107772 189132 107778
rect 189080 107714 189132 107720
rect 189092 107574 189120 107714
rect 189080 107568 189132 107574
rect 189080 107510 189132 107516
rect 189092 83745 189120 107510
rect 189736 95305 189764 135186
rect 189828 122398 189856 150418
rect 189920 133929 189948 155994
rect 190380 142154 190408 177278
rect 190460 166320 190512 166326
rect 190460 166262 190512 166268
rect 190288 142126 190408 142154
rect 190288 138553 190316 142126
rect 190366 138680 190422 138689
rect 190366 138615 190422 138624
rect 190274 138544 190330 138553
rect 190274 138479 190330 138488
rect 189998 136776 190054 136785
rect 189998 136711 190054 136720
rect 189906 133920 189962 133929
rect 189906 133855 189962 133864
rect 190012 131102 190040 136711
rect 190000 131096 190052 131102
rect 190000 131038 190052 131044
rect 190274 129840 190330 129849
rect 190274 129775 190330 129784
rect 190288 125594 190316 129775
rect 190380 125746 190408 138615
rect 190472 134745 190500 166262
rect 192496 158001 192524 243510
rect 192588 235958 192616 266970
rect 192668 249960 192720 249966
rect 192668 249902 192720 249908
rect 192680 240786 192708 249902
rect 192668 240780 192720 240786
rect 192668 240722 192720 240728
rect 192576 235952 192628 235958
rect 192576 235894 192628 235900
rect 193140 235346 193168 283455
rect 193404 246424 193456 246430
rect 193404 246366 193456 246372
rect 193416 238754 193444 246366
rect 193496 244928 193548 244934
rect 193496 244870 193548 244876
rect 193508 241074 193536 244870
rect 193678 244216 193734 244225
rect 193678 244151 193734 244160
rect 193586 242448 193642 242457
rect 193586 242383 193642 242392
rect 193600 241210 193628 242383
rect 193692 241369 193720 244151
rect 249156 242072 249208 242078
rect 194506 242040 194562 242049
rect 249156 242014 249208 242020
rect 249800 242072 249852 242078
rect 250166 242040 250222 242049
rect 249800 242014 249852 242020
rect 194506 241975 194562 241984
rect 193678 241360 193734 241369
rect 193678 241295 193734 241304
rect 193600 241182 193812 241210
rect 193508 241046 193720 241074
rect 193416 238726 193628 238754
rect 193600 238678 193628 238726
rect 193588 238672 193640 238678
rect 193588 238614 193640 238620
rect 193692 237386 193720 241046
rect 193680 237380 193732 237386
rect 193680 237322 193732 237328
rect 193128 235340 193180 235346
rect 193128 235282 193180 235288
rect 193312 204264 193364 204270
rect 193312 204206 193364 204212
rect 193128 187060 193180 187066
rect 193128 187002 193180 187008
rect 192576 167136 192628 167142
rect 192576 167078 192628 167084
rect 192482 157992 192538 158001
rect 192482 157927 192538 157936
rect 192588 153134 192616 167078
rect 192576 153128 192628 153134
rect 192576 153070 192628 153076
rect 192588 151814 192616 153070
rect 192588 151786 192984 151814
rect 191104 149864 191156 149870
rect 191104 149806 191156 149812
rect 190458 134736 190514 134745
rect 190458 134671 190514 134680
rect 190472 134026 190500 134671
rect 190460 134020 190512 134026
rect 190460 133962 190512 133968
rect 191116 132394 191144 149806
rect 192482 149152 192538 149161
rect 192482 149087 192538 149096
rect 191748 136604 191800 136610
rect 191748 136546 191800 136552
rect 191760 136377 191788 136546
rect 191746 136368 191802 136377
rect 191746 136303 191802 136312
rect 191746 135552 191802 135561
rect 191746 135487 191802 135496
rect 191760 135318 191788 135487
rect 191748 135312 191800 135318
rect 191748 135254 191800 135260
rect 192496 134473 192524 149087
rect 192956 139913 192984 151786
rect 193036 140480 193088 140486
rect 193036 140422 193088 140428
rect 192942 139904 192998 139913
rect 192942 139839 192998 139848
rect 191746 134464 191802 134473
rect 191746 134399 191802 134408
rect 192482 134464 192538 134473
rect 192482 134399 192538 134408
rect 191656 132456 191708 132462
rect 191656 132398 191708 132404
rect 191104 132388 191156 132394
rect 191104 132330 191156 132336
rect 190458 125760 190514 125769
rect 190380 125730 190458 125746
rect 190368 125724 190458 125730
rect 190420 125718 190458 125724
rect 190458 125695 190514 125704
rect 190368 125666 190420 125672
rect 190380 125635 190408 125666
rect 190276 125588 190328 125594
rect 190276 125530 190328 125536
rect 189816 122392 189868 122398
rect 189816 122334 189868 122340
rect 190368 122392 190420 122398
rect 190368 122334 190420 122340
rect 190380 121666 190408 122334
rect 190458 121680 190514 121689
rect 190380 121638 190458 121666
rect 190274 110800 190330 110809
rect 190274 110735 190330 110744
rect 190288 109002 190316 110735
rect 190276 108996 190328 109002
rect 190276 108938 190328 108944
rect 189816 98048 189868 98054
rect 189816 97990 189868 97996
rect 189722 95296 189778 95305
rect 189722 95231 189778 95240
rect 189828 89593 189856 97990
rect 189814 89584 189870 89593
rect 189814 89519 189870 89528
rect 189078 83736 189134 83745
rect 189078 83671 189134 83680
rect 189092 82929 189120 83671
rect 189078 82920 189134 82929
rect 189078 82855 189134 82864
rect 189722 82920 189778 82929
rect 189722 82855 189778 82864
rect 189736 49026 189764 82855
rect 190380 62830 190408 121638
rect 190458 121615 190514 121624
rect 191116 117609 191144 132330
rect 191668 131209 191696 132398
rect 191654 131200 191710 131209
rect 191654 131135 191710 131144
rect 191760 130914 191788 134399
rect 193048 132025 193076 140422
rect 193034 132016 193090 132025
rect 193034 131951 193090 131960
rect 191668 130886 191788 130914
rect 191668 129305 191696 130886
rect 191748 129736 191800 129742
rect 191748 129678 191800 129684
rect 191654 129296 191710 129305
rect 191654 129231 191710 129240
rect 191760 128489 191788 129678
rect 191746 128480 191802 128489
rect 191746 128415 191802 128424
rect 192298 127664 192354 127673
rect 192298 127599 192354 127608
rect 192312 127022 192340 127599
rect 192300 127016 192352 127022
rect 192300 126958 192352 126964
rect 192852 127016 192904 127022
rect 192852 126958 192904 126964
rect 192392 126880 192444 126886
rect 192392 126822 192444 126828
rect 192404 126585 192432 126822
rect 192390 126576 192446 126585
rect 192390 126511 192446 126520
rect 191746 123040 191802 123049
rect 191746 122975 191802 122984
rect 191760 122874 191788 122975
rect 191748 122868 191800 122874
rect 191748 122810 191800 122816
rect 191196 121440 191248 121446
rect 191194 121408 191196 121417
rect 191248 121408 191250 121417
rect 191194 121343 191250 121352
rect 191748 120692 191800 120698
rect 191748 120634 191800 120640
rect 191760 120329 191788 120634
rect 191746 120320 191802 120329
rect 191746 120255 191802 120264
rect 191748 120080 191800 120086
rect 191748 120022 191800 120028
rect 191760 119513 191788 120022
rect 191746 119504 191802 119513
rect 191746 119439 191802 119448
rect 191746 118688 191802 118697
rect 191746 118623 191802 118632
rect 191102 117600 191158 117609
rect 191102 117535 191158 117544
rect 191760 117434 191788 118623
rect 191748 117428 191800 117434
rect 191748 117370 191800 117376
rect 191748 117292 191800 117298
rect 191748 117234 191800 117240
rect 191286 116784 191342 116793
rect 191286 116719 191342 116728
rect 191300 116074 191328 116719
rect 191288 116068 191340 116074
rect 191288 116010 191340 116016
rect 191760 115977 191788 117234
rect 191746 115968 191802 115977
rect 191012 115932 191064 115938
rect 191746 115903 191802 115912
rect 191012 115874 191064 115880
rect 191024 115161 191052 115874
rect 191010 115152 191066 115161
rect 191010 115087 191066 115096
rect 191746 114064 191802 114073
rect 191746 113999 191802 114008
rect 191196 113280 191248 113286
rect 191194 113248 191196 113257
rect 191248 113248 191250 113257
rect 191760 113218 191788 113999
rect 191194 113183 191250 113192
rect 191748 113212 191800 113218
rect 191748 113154 191800 113160
rect 191564 112464 191616 112470
rect 191564 112406 191616 112412
rect 191380 111784 191432 111790
rect 191380 111726 191432 111732
rect 191392 110537 191420 111726
rect 191378 110528 191434 110537
rect 191378 110463 191434 110472
rect 191576 109721 191604 112406
rect 191562 109712 191618 109721
rect 191562 109647 191618 109656
rect 191196 108928 191248 108934
rect 191194 108896 191196 108905
rect 191248 108896 191250 108905
rect 191194 108831 191250 108840
rect 191194 107808 191250 107817
rect 191194 107743 191196 107752
rect 191248 107743 191250 107752
rect 191196 107714 191248 107720
rect 191748 107636 191800 107642
rect 191748 107578 191800 107584
rect 191760 107001 191788 107578
rect 191746 106992 191802 107001
rect 191746 106927 191802 106936
rect 191746 106176 191802 106185
rect 191746 106111 191802 106120
rect 191760 105942 191788 106111
rect 191748 105936 191800 105942
rect 191748 105878 191800 105884
rect 191746 105088 191802 105097
rect 191746 105023 191802 105032
rect 191760 104922 191788 105023
rect 191748 104916 191800 104922
rect 191748 104858 191800 104864
rect 191746 104272 191802 104281
rect 191746 104207 191802 104216
rect 191654 103456 191710 103465
rect 191654 103391 191710 103400
rect 191102 102640 191158 102649
rect 191102 102575 191158 102584
rect 190644 100700 190696 100706
rect 190644 100642 190696 100648
rect 190656 99929 190684 100642
rect 190642 99920 190698 99929
rect 190642 99855 190698 99864
rect 190644 97980 190696 97986
rect 190644 97922 190696 97928
rect 190656 97209 190684 97922
rect 190642 97200 190698 97209
rect 190642 97135 190698 97144
rect 191116 93945 191144 102575
rect 191668 102202 191696 103391
rect 191656 102196 191708 102202
rect 191656 102138 191708 102144
rect 191654 101552 191710 101561
rect 191654 101487 191710 101496
rect 191668 100774 191696 101487
rect 191656 100768 191708 100774
rect 191562 100736 191618 100745
rect 191656 100710 191708 100716
rect 191562 100671 191618 100680
rect 191576 99521 191604 100671
rect 191562 99512 191618 99521
rect 191562 99447 191618 99456
rect 191102 93936 191158 93945
rect 191102 93871 191158 93880
rect 191116 85377 191144 93871
rect 191102 85368 191158 85377
rect 191102 85303 191158 85312
rect 191576 83473 191604 99447
rect 191656 98116 191708 98122
rect 191656 98058 191708 98064
rect 191668 98025 191696 98058
rect 191654 98016 191710 98025
rect 191654 97951 191710 97960
rect 191654 94480 191710 94489
rect 191654 94415 191710 94424
rect 191562 83464 191618 83473
rect 191562 83399 191618 83408
rect 191668 77217 191696 94415
rect 191760 93786 191788 104207
rect 191760 93758 191880 93786
rect 191746 93664 191802 93673
rect 191746 93599 191802 93608
rect 191760 93158 191788 93599
rect 191748 93152 191800 93158
rect 191748 93094 191800 93100
rect 191852 92970 191880 93758
rect 191760 92942 191880 92970
rect 191760 84862 191788 92942
rect 191748 84856 191800 84862
rect 191748 84798 191800 84804
rect 191102 77208 191158 77217
rect 191102 77143 191158 77152
rect 191654 77208 191710 77217
rect 191654 77143 191710 77152
rect 190368 62824 190420 62830
rect 190368 62766 190420 62772
rect 191116 62121 191144 77143
rect 192864 71058 192892 126958
rect 193034 126576 193090 126585
rect 193034 126511 193090 126520
rect 192942 124944 192998 124953
rect 192942 124879 192998 124888
rect 192956 124846 192984 124879
rect 192944 124840 192996 124846
rect 192944 124782 192996 124788
rect 192852 71052 192904 71058
rect 192852 70994 192904 71000
rect 191102 62112 191158 62121
rect 191102 62047 191158 62056
rect 192956 53106 192984 124782
rect 192944 53100 192996 53106
rect 192944 53042 192996 53048
rect 189724 49020 189776 49026
rect 189724 48962 189776 48968
rect 193048 44878 193076 126511
rect 193140 96393 193168 187002
rect 193218 157448 193274 157457
rect 193218 157383 193274 157392
rect 193232 141114 193260 157383
rect 193324 142905 193352 204206
rect 193784 182889 193812 241182
rect 194520 238105 194548 241975
rect 194810 241590 195284 241618
rect 195256 240106 195284 241590
rect 197188 241534 197216 241604
rect 199594 241590 200068 241618
rect 197176 241528 197228 241534
rect 197176 241470 197228 241476
rect 196622 241088 196678 241097
rect 196622 241023 196678 241032
rect 195244 240100 195296 240106
rect 195244 240042 195296 240048
rect 194506 238096 194562 238105
rect 194506 238031 194562 238040
rect 195256 189786 195284 240042
rect 196636 234569 196664 241023
rect 197358 237960 197414 237969
rect 197358 237895 197414 237904
rect 196714 236056 196770 236065
rect 196714 235991 196770 236000
rect 196622 234560 196678 234569
rect 196622 234495 196678 234504
rect 196636 214577 196664 234495
rect 196728 223582 196756 235991
rect 197372 233209 197400 237895
rect 197358 233200 197414 233209
rect 197358 233135 197414 233144
rect 198646 233200 198702 233209
rect 198646 233135 198702 233144
rect 196716 223576 196768 223582
rect 196716 223518 196768 223524
rect 197268 223576 197320 223582
rect 197268 223518 197320 223524
rect 195978 214568 196034 214577
rect 195978 214503 196034 214512
rect 196622 214568 196678 214577
rect 196622 214503 196678 214512
rect 195992 203590 196020 214503
rect 195980 203584 196032 203590
rect 195980 203526 196032 203532
rect 196624 202224 196676 202230
rect 196624 202166 196676 202172
rect 195888 202156 195940 202162
rect 195888 202098 195940 202104
rect 195244 189780 195296 189786
rect 195244 189722 195296 189728
rect 195796 188352 195848 188358
rect 195796 188294 195848 188300
rect 193770 182880 193826 182889
rect 193770 182815 193826 182824
rect 195808 164966 195836 188294
rect 195796 164960 195848 164966
rect 195796 164902 195848 164908
rect 193864 164892 193916 164898
rect 193864 164834 193916 164840
rect 193876 157457 193904 164834
rect 195900 160138 195928 202098
rect 195980 175364 196032 175370
rect 195980 175306 196032 175312
rect 195992 175234 196020 175306
rect 195980 175228 196032 175234
rect 195980 175170 196032 175176
rect 194600 160132 194652 160138
rect 194600 160074 194652 160080
rect 195888 160132 195940 160138
rect 195888 160074 195940 160080
rect 193862 157448 193918 157457
rect 193862 157383 193918 157392
rect 194612 151814 194640 160074
rect 196636 157457 196664 202166
rect 196716 184204 196768 184210
rect 196716 184146 196768 184152
rect 196070 157448 196126 157457
rect 196070 157383 196126 157392
rect 196622 157448 196678 157457
rect 196622 157383 196678 157392
rect 194612 151786 195008 151814
rect 193310 142896 193366 142905
rect 193310 142831 193366 142840
rect 194690 142760 194746 142769
rect 194690 142695 194746 142704
rect 194704 142225 194732 142695
rect 194690 142216 194746 142225
rect 194690 142151 194746 142160
rect 193232 141086 193720 141114
rect 193692 140978 193720 141086
rect 193692 140950 194166 140978
rect 194704 140964 194732 142151
rect 194980 140978 195008 151786
rect 196084 140978 196112 157383
rect 196624 156664 196676 156670
rect 196624 156606 196676 156612
rect 196532 144220 196584 144226
rect 196532 144162 196584 144168
rect 194980 140950 195454 140978
rect 196006 140950 196112 140978
rect 196544 140964 196572 144162
rect 196636 142361 196664 156606
rect 196728 148374 196756 184146
rect 196808 163532 196860 163538
rect 196808 163474 196860 163480
rect 196716 148368 196768 148374
rect 196716 148310 196768 148316
rect 196820 143614 196848 163474
rect 197280 163441 197308 223518
rect 197360 195288 197412 195294
rect 197360 195230 197412 195236
rect 197266 163432 197322 163441
rect 197266 163367 197322 163376
rect 197372 150006 197400 195230
rect 197544 164960 197596 164966
rect 197544 164902 197596 164908
rect 197360 150000 197412 150006
rect 197360 149942 197412 149948
rect 196808 143608 196860 143614
rect 196808 143550 196860 143556
rect 196622 142352 196678 142361
rect 196622 142287 196678 142296
rect 193232 140826 193614 140842
rect 193220 140820 193614 140826
rect 193272 140814 193614 140820
rect 193220 140762 193272 140768
rect 193312 140752 193364 140758
rect 193312 140694 193364 140700
rect 193324 137970 193352 140694
rect 196636 140434 196664 142287
rect 197556 141250 197584 164902
rect 198660 158137 198688 233135
rect 200040 200802 200068 241590
rect 201972 237318 202000 241604
rect 201500 237312 201552 237318
rect 201500 237254 201552 237260
rect 201960 237312 202012 237318
rect 201960 237254 202012 237260
rect 200762 236600 200818 236609
rect 200762 236535 200818 236544
rect 200028 200796 200080 200802
rect 200028 200738 200080 200744
rect 200304 168360 200356 168366
rect 200304 168302 200356 168308
rect 198740 166320 198792 166326
rect 198740 166262 198792 166268
rect 198752 161498 198780 166262
rect 198740 161492 198792 161498
rect 198740 161434 198792 161440
rect 198646 158128 198702 158137
rect 198646 158063 198702 158072
rect 198752 151814 198780 161434
rect 198752 151786 199332 151814
rect 197636 150000 197688 150006
rect 197636 149942 197688 149948
rect 197372 141222 197584 141250
rect 197372 140486 197400 141222
rect 197648 140978 197676 149942
rect 198004 145580 198056 145586
rect 198004 145522 198056 145528
rect 198832 145580 198884 145586
rect 198832 145522 198884 145528
rect 198016 140978 198044 145522
rect 198844 140978 198872 145522
rect 199304 140978 199332 151786
rect 200212 144492 200264 144498
rect 200212 144434 200264 144440
rect 197648 140950 197846 140978
rect 198016 140950 198398 140978
rect 198844 140950 198950 140978
rect 199304 140950 199686 140978
rect 200224 140964 200252 144434
rect 200316 140978 200344 168302
rect 200776 153785 200804 236535
rect 201512 153882 201540 237254
rect 203614 232520 203670 232529
rect 203614 232455 203670 232464
rect 203524 229764 203576 229770
rect 203524 229706 203576 229712
rect 202144 185632 202196 185638
rect 202144 185574 202196 185580
rect 202156 173194 202184 185574
rect 203536 180130 203564 229706
rect 203628 227633 203656 232455
rect 204364 227662 204392 241604
rect 205732 235952 205784 235958
rect 205732 235894 205784 235900
rect 205744 235482 205772 235894
rect 206756 235482 206784 241604
rect 209044 240780 209096 240786
rect 209044 240722 209096 240728
rect 207664 236700 207716 236706
rect 207664 236642 207716 236648
rect 205732 235476 205784 235482
rect 205732 235418 205784 235424
rect 206744 235476 206796 235482
rect 206744 235418 206796 235424
rect 204352 227656 204404 227662
rect 203614 227624 203670 227633
rect 204352 227598 204404 227604
rect 203614 227559 203670 227568
rect 204904 222896 204956 222902
rect 204904 222838 204956 222844
rect 204916 216617 204944 222838
rect 204902 216608 204958 216617
rect 204902 216543 204958 216552
rect 204916 215393 204944 216543
rect 204902 215384 204958 215393
rect 204902 215319 204958 215328
rect 205546 215384 205602 215393
rect 205546 215319 205602 215328
rect 204260 184952 204312 184958
rect 204260 184894 204312 184900
rect 203524 180124 203576 180130
rect 203524 180066 203576 180072
rect 202880 179444 202932 179450
rect 202880 179386 202932 179392
rect 201592 173188 201644 173194
rect 201592 173130 201644 173136
rect 202144 173188 202196 173194
rect 202144 173130 202196 173136
rect 201500 153876 201552 153882
rect 201500 153818 201552 153824
rect 200762 153776 200818 153785
rect 200762 153711 200818 153720
rect 201604 148345 201632 173130
rect 202788 158024 202840 158030
rect 202788 157966 202840 157972
rect 202800 154630 202828 157966
rect 201684 154624 201736 154630
rect 201684 154566 201736 154572
rect 202788 154624 202840 154630
rect 202788 154566 202840 154572
rect 201696 151814 201724 154566
rect 201696 151786 202184 151814
rect 201590 148336 201646 148345
rect 201590 148271 201646 148280
rect 202052 143676 202104 143682
rect 202052 143618 202104 143624
rect 201316 143608 201368 143614
rect 201316 143550 201368 143556
rect 200316 140950 200790 140978
rect 201328 140964 201356 143550
rect 202064 140964 202092 143618
rect 202156 140978 202184 151786
rect 202156 140950 202630 140978
rect 197360 140480 197412 140486
rect 196806 140448 196862 140457
rect 196636 140406 196806 140434
rect 196862 140406 197110 140434
rect 202892 140457 202920 179386
rect 203156 141432 203208 141438
rect 203156 141374 203208 141380
rect 203168 140842 203196 141374
rect 204272 141137 204300 184894
rect 204904 175296 204956 175302
rect 204904 175238 204956 175244
rect 204916 154970 204944 175238
rect 205560 155961 205588 215319
rect 205744 156670 205772 235418
rect 207018 177304 207074 177313
rect 207018 177239 207074 177248
rect 207032 176769 207060 177239
rect 207676 176769 207704 236642
rect 207756 181484 207808 181490
rect 207756 181426 207808 181432
rect 205822 176760 205878 176769
rect 205822 176695 205878 176704
rect 207018 176760 207074 176769
rect 207018 176695 207074 176704
rect 207662 176760 207718 176769
rect 207662 176695 207718 176704
rect 205836 172514 205864 176695
rect 205824 172508 205876 172514
rect 205824 172450 205876 172456
rect 205732 156664 205784 156670
rect 205732 156606 205784 156612
rect 205546 155952 205602 155961
rect 205546 155887 205602 155896
rect 204352 154964 204404 154970
rect 204352 154906 204404 154912
rect 204904 154964 204956 154970
rect 204904 154906 204956 154912
rect 204364 151814 204392 154906
rect 204916 154630 204944 154906
rect 204904 154624 204956 154630
rect 204904 154566 204956 154572
rect 204364 151786 204668 151814
rect 204442 149696 204498 149705
rect 204442 149631 204498 149640
rect 204258 141128 204314 141137
rect 204258 141063 204314 141072
rect 204456 140964 204484 149631
rect 204640 140978 204668 151786
rect 205454 140992 205510 141001
rect 204640 140950 205022 140978
rect 205836 140978 205864 172450
rect 206836 144220 206888 144226
rect 206836 144162 206888 144168
rect 206848 142254 206876 144162
rect 207032 143313 207060 176695
rect 207112 156052 207164 156058
rect 207112 155994 207164 156000
rect 207124 152522 207152 155994
rect 207112 152516 207164 152522
rect 207112 152458 207164 152464
rect 207110 145072 207166 145081
rect 207110 145007 207166 145016
rect 207018 143304 207074 143313
rect 207018 143239 207074 143248
rect 206836 142248 206888 142254
rect 206836 142190 206888 142196
rect 205510 140950 205574 140978
rect 205836 140950 206310 140978
rect 206848 140964 206876 142190
rect 207124 140978 207152 145007
rect 207768 144498 207796 181426
rect 208400 165640 208452 165646
rect 208400 165582 208452 165588
rect 208412 162858 208440 165582
rect 208400 162852 208452 162858
rect 208400 162794 208452 162800
rect 208412 151814 208440 162794
rect 209056 151814 209084 240722
rect 209148 239426 209176 241604
rect 211554 241590 211844 241618
rect 211816 240009 211844 241590
rect 213276 241596 213328 241602
rect 213276 241538 213328 241544
rect 213288 240106 213316 241538
rect 213276 240100 213328 240106
rect 213276 240042 213328 240048
rect 211802 240000 211858 240009
rect 211802 239935 211858 239944
rect 209136 239420 209188 239426
rect 209136 239362 209188 239368
rect 210424 232552 210476 232558
rect 210424 232494 210476 232500
rect 210436 222193 210464 232494
rect 211816 224233 211844 239935
rect 213932 238746 213960 241604
rect 213920 238740 213972 238746
rect 213920 238682 213972 238688
rect 213932 237454 213960 238682
rect 215300 238672 215352 238678
rect 215300 238614 215352 238620
rect 215312 238406 215340 238614
rect 216324 238406 216352 241604
rect 215300 238400 215352 238406
rect 215300 238342 215352 238348
rect 216312 238400 216364 238406
rect 216312 238342 216364 238348
rect 213920 237448 213972 237454
rect 213920 237390 213972 237396
rect 214656 237448 214708 237454
rect 214656 237390 214708 237396
rect 213184 235272 213236 235278
rect 213184 235214 213236 235220
rect 211802 224224 211858 224233
rect 211802 224159 211858 224168
rect 210422 222184 210478 222193
rect 210422 222119 210478 222128
rect 211066 222184 211122 222193
rect 211066 222119 211122 222128
rect 210422 171184 210478 171193
rect 210422 171119 210478 171128
rect 210436 164218 210464 171119
rect 210424 164212 210476 164218
rect 210424 164154 210476 164160
rect 210436 161474 210464 164154
rect 210068 161446 210464 161474
rect 210068 151814 210096 161446
rect 208412 151786 208900 151814
rect 209056 151786 209544 151814
rect 210068 151786 210648 151814
rect 208490 151192 208546 151201
rect 208490 151127 208546 151136
rect 208504 146334 208532 151127
rect 208492 146328 208544 146334
rect 208492 146270 208544 146276
rect 207756 144492 207808 144498
rect 207756 144434 207808 144440
rect 208122 143304 208178 143313
rect 208122 143239 208178 143248
rect 207124 140950 207414 140978
rect 205454 140927 205510 140936
rect 203168 140828 203472 140842
rect 203182 140826 203472 140828
rect 203182 140820 203484 140826
rect 203182 140814 203432 140820
rect 203432 140762 203484 140768
rect 197360 140422 197412 140428
rect 202878 140448 202934 140457
rect 196806 140383 196862 140392
rect 202878 140383 202934 140392
rect 203522 140448 203578 140457
rect 208136 140434 208164 143239
rect 208504 140978 208532 146270
rect 208872 140978 208900 151786
rect 208504 140950 208702 140978
rect 208872 140950 209254 140978
rect 209516 140593 209544 151786
rect 209872 144968 209924 144974
rect 209872 144910 209924 144916
rect 209502 140584 209558 140593
rect 209884 140570 209912 144910
rect 210514 144120 210570 144129
rect 210514 144055 210570 144064
rect 210528 140964 210556 144055
rect 210620 140978 210648 151786
rect 211080 151065 211108 222119
rect 213196 218754 213224 235214
rect 214564 222896 214616 222902
rect 214564 222838 214616 222844
rect 213274 222320 213330 222329
rect 213274 222255 213330 222264
rect 213288 219366 213316 222255
rect 213276 219360 213328 219366
rect 213276 219302 213328 219308
rect 213184 218748 213236 218754
rect 213184 218690 213236 218696
rect 211802 189680 211858 189689
rect 211802 189615 211858 189624
rect 211158 156088 211214 156097
rect 211158 156023 211214 156032
rect 211172 153202 211200 156023
rect 211160 153196 211212 153202
rect 211160 153138 211212 153144
rect 211066 151056 211122 151065
rect 211066 150991 211122 151000
rect 211172 140978 211200 153138
rect 211816 149705 211844 189615
rect 213184 175364 213236 175370
rect 213184 175306 213236 175312
rect 211802 149696 211858 149705
rect 211802 149631 211858 149640
rect 211896 147688 211948 147694
rect 211896 147630 211948 147636
rect 211804 142180 211856 142186
rect 211804 142122 211856 142128
rect 210620 140950 211094 140978
rect 211172 140950 211646 140978
rect 211816 140706 211844 142122
rect 211908 140978 211936 147630
rect 213196 146266 213224 175306
rect 214576 169794 214604 222838
rect 214668 192545 214696 237390
rect 214654 192536 214710 192545
rect 214654 192471 214710 192480
rect 213920 169788 213972 169794
rect 213920 169730 213972 169736
rect 214564 169788 214616 169794
rect 214564 169730 214616 169736
rect 213274 159352 213330 159361
rect 213274 159287 213330 159296
rect 213184 146260 213236 146266
rect 213184 146202 213236 146208
rect 212814 142488 212870 142497
rect 212814 142423 212870 142432
rect 212828 142186 212856 142423
rect 213288 142322 213316 159287
rect 213932 148374 213960 169730
rect 215312 153921 215340 238342
rect 216678 238096 216734 238105
rect 216678 238031 216734 238040
rect 215390 237960 215446 237969
rect 215390 237895 215446 237904
rect 215404 230450 215432 237895
rect 216692 237289 216720 238031
rect 216678 237280 216734 237289
rect 216678 237215 216734 237224
rect 217966 237280 218022 237289
rect 217966 237215 218022 237224
rect 215944 231192 215996 231198
rect 215944 231134 215996 231140
rect 215392 230444 215444 230450
rect 215392 230386 215444 230392
rect 215956 220794 215984 231134
rect 215944 220788 215996 220794
rect 215944 220730 215996 220736
rect 215956 164393 215984 220730
rect 217980 169794 218008 237215
rect 218716 184210 218744 241604
rect 221108 238746 221136 241604
rect 223500 240038 223528 241604
rect 222200 240032 222252 240038
rect 222200 239974 222252 239980
rect 223488 240032 223540 240038
rect 223488 239974 223540 239980
rect 221096 238740 221148 238746
rect 221096 238682 221148 238688
rect 221108 236706 221136 238682
rect 221096 236700 221148 236706
rect 221096 236642 221148 236648
rect 220820 235340 220872 235346
rect 220820 235282 220872 235288
rect 219440 224256 219492 224262
rect 219440 224198 219492 224204
rect 218704 184204 218756 184210
rect 218704 184146 218756 184152
rect 216864 169788 216916 169794
rect 216864 169730 216916 169736
rect 217968 169788 218020 169794
rect 217968 169730 218020 169736
rect 215942 164384 215998 164393
rect 215942 164319 215998 164328
rect 215956 161474 215984 164319
rect 215496 161446 215984 161474
rect 215392 155236 215444 155242
rect 215392 155178 215444 155184
rect 215298 153912 215354 153921
rect 215298 153847 215354 153856
rect 213920 148368 213972 148374
rect 213920 148310 213972 148316
rect 213932 147694 213960 148310
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 215404 147014 215432 155178
rect 215392 147008 215444 147014
rect 215392 146950 215444 146956
rect 214564 146328 214616 146334
rect 214564 146270 214616 146276
rect 214012 143540 214064 143546
rect 214012 143482 214064 143488
rect 213276 142316 213328 142322
rect 213276 142258 213328 142264
rect 212816 142180 212868 142186
rect 212816 142122 212868 142128
rect 212828 140978 212856 142122
rect 213288 140978 213316 142258
rect 211908 140950 212382 140978
rect 212828 140950 212934 140978
rect 213288 140950 213486 140978
rect 214024 140964 214052 143482
rect 214380 140888 214432 140894
rect 214576 140842 214604 146270
rect 215300 142248 215352 142254
rect 215300 142190 215352 142196
rect 214432 140836 214774 140842
rect 214380 140830 214774 140836
rect 214392 140814 214774 140830
rect 211894 140720 211950 140729
rect 211816 140678 211894 140706
rect 211894 140655 211950 140664
rect 209806 140554 210096 140570
rect 209806 140548 210108 140554
rect 209806 140542 210056 140548
rect 209502 140519 209558 140528
rect 210056 140490 210108 140496
rect 208214 140448 208270 140457
rect 203578 140406 203918 140434
rect 208136 140420 208214 140434
rect 208150 140406 208214 140420
rect 203522 140383 203578 140392
rect 215312 140434 215340 142190
rect 215496 140978 215524 161446
rect 216680 149728 216732 149734
rect 216680 149670 216732 149676
rect 216220 147008 216272 147014
rect 216220 146950 216272 146956
rect 216232 140978 216260 146950
rect 216692 140978 216720 149670
rect 216772 146260 216824 146266
rect 216772 146202 216824 146208
rect 216784 141250 216812 146202
rect 216876 143546 216904 169730
rect 218244 150476 218296 150482
rect 218244 150418 218296 150424
rect 216864 143540 216916 143546
rect 216864 143482 216916 143488
rect 218256 143449 218284 150418
rect 218336 149796 218388 149802
rect 218336 149738 218388 149744
rect 218348 147801 218376 149738
rect 219452 149569 219480 224198
rect 220084 216028 220136 216034
rect 220084 215970 220136 215976
rect 220096 210905 220124 215970
rect 220082 210896 220138 210905
rect 220082 210831 220138 210840
rect 220096 167113 220124 210831
rect 220832 173942 220860 235282
rect 222212 230489 222240 239974
rect 225984 239630 226012 241604
rect 227732 241590 228390 241618
rect 224868 239624 224920 239630
rect 224868 239566 224920 239572
rect 225972 239624 226024 239630
rect 225972 239566 226024 239572
rect 222844 235340 222896 235346
rect 222844 235282 222896 235288
rect 222198 230480 222254 230489
rect 222198 230415 222254 230424
rect 220820 173936 220872 173942
rect 220820 173878 220872 173884
rect 221464 173936 221516 173942
rect 221464 173878 221516 173884
rect 220082 167104 220138 167113
rect 220082 167039 220138 167048
rect 219438 149560 219494 149569
rect 219438 149495 219494 149504
rect 218334 147792 218390 147801
rect 218334 147727 218390 147736
rect 218242 143440 218298 143449
rect 218242 143375 218298 143384
rect 216784 141222 217272 141250
rect 217244 140978 217272 141222
rect 215496 140950 215878 140978
rect 216232 140950 216614 140978
rect 216692 140950 217166 140978
rect 217244 140950 217718 140978
rect 218256 140964 218284 143375
rect 218348 142154 218376 147727
rect 220096 146441 220124 167039
rect 220820 158772 220872 158778
rect 220820 158714 220872 158720
rect 220174 149560 220230 149569
rect 220174 149495 220230 149504
rect 218794 146432 218850 146441
rect 218794 146367 218850 146376
rect 220082 146432 220138 146441
rect 220082 146367 220138 146376
rect 218348 142126 218560 142154
rect 218532 140978 218560 142126
rect 218808 141438 218836 146367
rect 220096 143546 220124 146367
rect 219532 143540 219584 143546
rect 219532 143482 219584 143488
rect 220084 143540 220136 143546
rect 220084 143482 220136 143488
rect 218796 141432 218848 141438
rect 218796 141374 218848 141380
rect 218532 140950 219006 140978
rect 219544 140964 219572 143482
rect 219992 142180 220044 142186
rect 219992 142122 220044 142128
rect 220004 140978 220032 142122
rect 220188 141137 220216 149495
rect 220174 141128 220230 141137
rect 220174 141063 220230 141072
rect 220004 140950 220110 140978
rect 220832 140964 220860 158714
rect 221476 151814 221504 173878
rect 222212 161906 222240 230415
rect 222292 173868 222344 173874
rect 222292 173810 222344 173816
rect 222304 172582 222332 173810
rect 222292 172576 222344 172582
rect 222292 172518 222344 172524
rect 222200 161900 222252 161906
rect 222200 161842 222252 161848
rect 222212 161566 222240 161842
rect 222200 161560 222252 161566
rect 222200 161502 222252 161508
rect 222304 155242 222332 172518
rect 222856 171154 222884 235282
rect 222936 191140 222988 191146
rect 222936 191082 222988 191088
rect 222948 173874 222976 191082
rect 222936 173868 222988 173874
rect 222936 173810 222988 173816
rect 222844 171148 222896 171154
rect 222844 171090 222896 171096
rect 222292 155236 222344 155242
rect 222292 155178 222344 155184
rect 222198 154728 222254 154737
rect 222198 154663 222254 154672
rect 222212 154562 222240 154663
rect 222200 154556 222252 154562
rect 222200 154498 222252 154504
rect 221476 151786 221964 151814
rect 220912 148436 220964 148442
rect 220912 148378 220964 148384
rect 220924 140978 220952 148378
rect 221936 142361 221964 151786
rect 221922 142352 221978 142361
rect 221922 142287 221978 142296
rect 221464 142248 221516 142254
rect 221464 142190 221516 142196
rect 220924 140950 221398 140978
rect 220004 140865 220032 140950
rect 219990 140856 220046 140865
rect 219990 140791 220046 140800
rect 221476 140758 221504 142190
rect 221936 140964 221964 142287
rect 222212 140978 222240 154498
rect 222856 142154 222884 171090
rect 222936 161900 222988 161906
rect 222936 161842 222988 161848
rect 222948 144906 222976 161842
rect 224224 160200 224276 160206
rect 224224 160142 224276 160148
rect 223580 153332 223632 153338
rect 223580 153274 223632 153280
rect 222936 144900 222988 144906
rect 222936 144842 222988 144848
rect 223212 142248 223264 142254
rect 223212 142190 223264 142196
rect 223224 142154 223252 142190
rect 222856 142126 223252 142154
rect 222212 140950 222502 140978
rect 223224 140964 223252 142126
rect 223592 141234 223620 153274
rect 223762 141400 223818 141409
rect 223762 141335 223818 141344
rect 223580 141228 223632 141234
rect 223580 141170 223632 141176
rect 223776 140964 223804 141335
rect 221464 140752 221516 140758
rect 221464 140694 221516 140700
rect 215392 140480 215444 140486
rect 215312 140428 215392 140434
rect 215312 140422 215444 140428
rect 224236 140434 224264 160142
rect 224880 149870 224908 239566
rect 226616 189780 226668 189786
rect 226616 189722 226668 189728
rect 225052 157412 225104 157418
rect 225052 157354 225104 157360
rect 225064 151814 225092 157354
rect 226432 155984 226484 155990
rect 226432 155926 226484 155932
rect 225064 151786 225276 151814
rect 224960 150544 225012 150550
rect 224960 150486 225012 150492
rect 224868 149864 224920 149870
rect 224868 149806 224920 149812
rect 224880 149734 224908 149806
rect 224868 149728 224920 149734
rect 224868 149670 224920 149676
rect 224500 141228 224552 141234
rect 224500 141170 224552 141176
rect 224512 140978 224540 141170
rect 224512 140950 224894 140978
rect 224592 140480 224644 140486
rect 224236 140428 224592 140434
rect 224236 140422 224644 140428
rect 215312 140420 215432 140422
rect 215326 140406 215432 140420
rect 224236 140406 224632 140422
rect 208214 140383 208270 140392
rect 193312 137964 193364 137970
rect 193312 137906 193364 137912
rect 224972 136626 225000 150486
rect 225050 136640 225106 136649
rect 224972 136598 225050 136626
rect 225050 136575 225106 136584
rect 193218 124128 193274 124137
rect 193218 124063 193274 124072
rect 193232 104281 193260 124063
rect 225248 123865 225276 151786
rect 225604 142180 225656 142186
rect 225604 142122 225656 142128
rect 225234 123856 225290 123865
rect 225234 123791 225290 123800
rect 225616 112538 225644 142122
rect 225696 140480 225748 140486
rect 225696 140422 225748 140428
rect 225708 122126 225736 140422
rect 226340 139392 226392 139398
rect 226340 139334 226392 139340
rect 226352 139097 226380 139334
rect 226338 139088 226394 139097
rect 226338 139023 226394 139032
rect 226338 136368 226394 136377
rect 226338 136303 226394 136312
rect 226352 135250 226380 136303
rect 226340 135244 226392 135250
rect 226340 135186 226392 135192
rect 226340 133884 226392 133890
rect 226340 133826 226392 133832
rect 226352 133385 226380 133826
rect 226444 133550 226472 155926
rect 226524 144900 226576 144906
rect 226524 144842 226576 144848
rect 226432 133544 226484 133550
rect 226432 133486 226484 133492
rect 226338 133376 226394 133385
rect 226338 133311 226394 133320
rect 226340 132456 226392 132462
rect 226340 132398 226392 132404
rect 226352 132025 226380 132398
rect 226338 132016 226394 132025
rect 226338 131951 226394 131960
rect 226536 129062 226564 144842
rect 226524 129056 226576 129062
rect 226524 128998 226576 129004
rect 226340 126948 226392 126954
rect 226340 126890 226392 126896
rect 226352 126585 226380 126890
rect 226338 126576 226394 126585
rect 226338 126511 226394 126520
rect 226524 124772 226576 124778
rect 226524 124714 226576 124720
rect 226536 124681 226564 124714
rect 226522 124672 226578 124681
rect 226522 124607 226578 124616
rect 226340 124160 226392 124166
rect 226340 124102 226392 124108
rect 226352 123049 226380 124102
rect 226338 123040 226394 123049
rect 226338 122975 226394 122984
rect 226340 122800 226392 122806
rect 226340 122742 226392 122748
rect 226352 122233 226380 122742
rect 226338 122224 226394 122233
rect 226338 122159 226394 122168
rect 225696 122120 225748 122126
rect 225696 122062 225748 122068
rect 226432 121440 226484 121446
rect 226432 121382 226484 121388
rect 226444 120329 226472 121382
rect 226430 120320 226486 120329
rect 226430 120255 226486 120264
rect 226522 118416 226578 118425
rect 226522 118351 226578 118360
rect 226536 117434 226564 118351
rect 226524 117428 226576 117434
rect 226524 117370 226576 117376
rect 226338 114880 226394 114889
rect 226338 114815 226394 114824
rect 226352 114578 226380 114815
rect 226340 114572 226392 114578
rect 226340 114514 226392 114520
rect 225604 112532 225656 112538
rect 225604 112474 225656 112480
rect 226338 111344 226394 111353
rect 226338 111279 226394 111288
rect 226352 111178 226380 111279
rect 226340 111172 226392 111178
rect 226340 111114 226392 111120
rect 226524 111104 226576 111110
rect 226524 111046 226576 111052
rect 226536 110537 226564 111046
rect 226522 110528 226578 110537
rect 226522 110463 226578 110472
rect 225604 109744 225656 109750
rect 225142 109712 225198 109721
rect 225604 109686 225656 109692
rect 225142 109647 225198 109656
rect 225050 104952 225106 104961
rect 224972 104910 225050 104938
rect 193218 104272 193274 104281
rect 193218 104207 193274 104216
rect 193126 96384 193182 96393
rect 193126 96319 193182 96328
rect 193140 95266 193168 96319
rect 193128 95260 193180 95266
rect 193128 95202 193180 95208
rect 193140 91798 193168 95202
rect 193404 94512 193456 94518
rect 193404 94454 193456 94460
rect 193128 91792 193180 91798
rect 193128 91734 193180 91740
rect 193416 89622 193444 94454
rect 199106 93392 199162 93401
rect 198950 93364 199106 93378
rect 198936 93350 199106 93364
rect 198936 92834 198964 93350
rect 199106 93327 199162 93336
rect 205730 93392 205786 93401
rect 208950 93392 209006 93401
rect 205786 93350 206126 93378
rect 208702 93364 208950 93378
rect 208688 93350 208950 93364
rect 205730 93327 205786 93336
rect 200394 92848 200450 92857
rect 193508 92806 193614 92834
rect 193784 92806 194166 92834
rect 193404 89616 193456 89622
rect 193404 89558 193456 89564
rect 193508 88482 193536 92806
rect 193232 88454 193536 88482
rect 193232 75818 193260 88454
rect 193784 84194 193812 92806
rect 194704 85513 194732 92820
rect 194888 92806 195270 92834
rect 194690 85504 194746 85513
rect 194690 85439 194746 85448
rect 194888 84194 194916 92806
rect 195886 85504 195942 85513
rect 195886 85439 195942 85448
rect 193324 84182 193812 84194
rect 193312 84176 193812 84182
rect 193364 84166 193812 84176
rect 194612 84166 194916 84194
rect 193312 84118 193364 84124
rect 193324 82890 193352 84118
rect 193312 82884 193364 82890
rect 193312 82826 193364 82832
rect 193956 82884 194008 82890
rect 193956 82826 194008 82832
rect 193220 75812 193272 75818
rect 193220 75754 193272 75760
rect 193864 75812 193916 75818
rect 193864 75754 193916 75760
rect 193876 63510 193904 75754
rect 193864 63504 193916 63510
rect 193864 63446 193916 63452
rect 193036 44872 193088 44878
rect 193036 44814 193088 44820
rect 193876 25566 193904 63446
rect 193968 58682 193996 82826
rect 194612 74458 194640 84166
rect 195900 78577 195928 85439
rect 195992 81258 196020 92820
rect 196544 92721 196572 92820
rect 196530 92712 196586 92721
rect 196530 92647 196586 92656
rect 196072 88256 196124 88262
rect 196070 88224 196072 88233
rect 196124 88224 196126 88233
rect 196070 88159 196126 88168
rect 197096 87961 197124 92820
rect 197464 92806 197662 92834
rect 198016 92806 198398 92834
rect 198752 92820 198964 92834
rect 198752 92806 198950 92820
rect 199396 92806 199502 92834
rect 197082 87952 197138 87961
rect 197082 87887 197138 87896
rect 197360 85604 197412 85610
rect 197360 85546 197412 85552
rect 195980 81252 196032 81258
rect 195980 81194 196032 81200
rect 195992 80102 196020 81194
rect 195980 80096 196032 80102
rect 195980 80038 196032 80044
rect 196624 80096 196676 80102
rect 196624 80038 196676 80044
rect 195886 78568 195942 78577
rect 195886 78503 195942 78512
rect 194600 74452 194652 74458
rect 194600 74394 194652 74400
rect 194612 73234 194640 74394
rect 194600 73228 194652 73234
rect 194600 73170 194652 73176
rect 195244 73228 195296 73234
rect 195244 73170 195296 73176
rect 193956 58676 194008 58682
rect 193956 58618 194008 58624
rect 195256 35222 195284 73170
rect 195244 35216 195296 35222
rect 195244 35158 195296 35164
rect 193864 25560 193916 25566
rect 193864 25502 193916 25508
rect 188988 11756 189040 11762
rect 188988 11698 189040 11704
rect 196636 8974 196664 80038
rect 197372 73098 197400 85546
rect 197464 78606 197492 92806
rect 198016 85610 198044 92806
rect 198004 85604 198056 85610
rect 198004 85546 198056 85552
rect 197452 78600 197504 78606
rect 197452 78542 197504 78548
rect 198004 78600 198056 78606
rect 198004 78542 198056 78548
rect 197360 73092 197412 73098
rect 197360 73034 197412 73040
rect 198016 10334 198044 78542
rect 198752 77994 198780 92806
rect 199396 89622 199424 92806
rect 200224 92449 200252 92820
rect 203338 92848 203394 92857
rect 200450 92806 200790 92834
rect 200868 92806 201342 92834
rect 201512 92806 201894 92834
rect 200394 92783 200450 92792
rect 200210 92440 200266 92449
rect 200210 92375 200266 92384
rect 199384 89616 199436 89622
rect 199384 89558 199436 89564
rect 198740 77988 198792 77994
rect 198740 77930 198792 77936
rect 199396 57254 199424 89558
rect 200868 88482 200896 92806
rect 200946 92440 201002 92449
rect 200946 92375 201002 92384
rect 200132 88454 200896 88482
rect 200132 82754 200160 88454
rect 200960 84194 200988 92375
rect 200776 84166 200988 84194
rect 200120 82748 200172 82754
rect 200120 82690 200172 82696
rect 200776 71777 200804 84166
rect 201408 82748 201460 82754
rect 201408 82690 201460 82696
rect 201420 82142 201448 82690
rect 201408 82136 201460 82142
rect 201408 82078 201460 82084
rect 201512 74526 201540 92806
rect 202616 92177 202644 92820
rect 202984 92806 203338 92834
rect 202602 92168 202658 92177
rect 202602 92103 202658 92112
rect 202144 91792 202196 91798
rect 202144 91734 202196 91740
rect 201500 74520 201552 74526
rect 201500 74462 201552 74468
rect 200762 71768 200818 71777
rect 200762 71703 200818 71712
rect 199384 57248 199436 57254
rect 199384 57190 199436 57196
rect 200776 13122 200804 71703
rect 201512 67590 201540 74462
rect 201500 67584 201552 67590
rect 201500 67526 201552 67532
rect 202156 50386 202184 91734
rect 202984 63578 203012 92806
rect 208688 92834 208716 93350
rect 211710 93392 211766 93401
rect 211646 93350 211710 93378
rect 208950 93327 209006 93336
rect 211710 93327 211766 93336
rect 224774 93392 224830 93401
rect 224830 93350 224894 93378
rect 224774 93327 224830 93336
rect 212446 92984 212502 92993
rect 212446 92919 212502 92928
rect 212460 92834 212488 92919
rect 224038 92848 224094 92857
rect 203338 92783 203394 92792
rect 203720 90545 203748 92820
rect 203706 90536 203762 90545
rect 203706 90471 203762 90480
rect 203720 89622 203748 90471
rect 204456 90409 204484 92820
rect 204442 90400 204498 90409
rect 204442 90335 204498 90344
rect 203708 89616 203760 89622
rect 203708 89558 203760 89564
rect 204456 86873 204484 90335
rect 205008 89729 205036 92820
rect 205100 92806 205574 92834
rect 206296 92806 206862 92834
rect 205100 91089 205128 92806
rect 205086 91080 205142 91089
rect 205086 91015 205142 91024
rect 204994 89720 205050 89729
rect 204994 89655 205050 89664
rect 204442 86864 204498 86873
rect 204442 86799 204498 86808
rect 205100 84194 205128 91015
rect 206296 84194 206324 92806
rect 207400 88262 207428 92820
rect 207492 92806 207966 92834
rect 208412 92820 208716 92834
rect 208412 92806 208702 92820
rect 206376 88256 206428 88262
rect 206376 88198 206428 88204
rect 207388 88256 207440 88262
rect 207388 88198 207440 88204
rect 204916 84166 205128 84194
rect 205652 84166 206324 84194
rect 202972 63572 203024 63578
rect 202972 63514 203024 63520
rect 202984 57934 203012 63514
rect 202972 57928 203024 57934
rect 202972 57870 203024 57876
rect 202144 50380 202196 50386
rect 202144 50322 202196 50328
rect 204916 37262 204944 84166
rect 205652 79966 205680 84166
rect 205640 79960 205692 79966
rect 205640 79902 205692 79908
rect 205652 79558 205680 79902
rect 205640 79552 205692 79558
rect 205640 79494 205692 79500
rect 206284 79552 206336 79558
rect 206284 79494 206336 79500
rect 205546 79384 205602 79393
rect 205546 79319 205602 79328
rect 205560 78713 205588 79319
rect 205546 78704 205602 78713
rect 205546 78639 205602 78648
rect 204904 37256 204956 37262
rect 204904 37198 204956 37204
rect 205560 19990 205588 78639
rect 205548 19984 205600 19990
rect 205548 19926 205600 19932
rect 206296 17270 206324 79494
rect 206388 56506 206416 88198
rect 207492 84194 207520 92806
rect 207032 84166 207520 84194
rect 207032 73166 207060 84166
rect 207020 73160 207072 73166
rect 207020 73102 207072 73108
rect 207032 72486 207060 73102
rect 207020 72480 207072 72486
rect 207020 72422 207072 72428
rect 206376 56500 206428 56506
rect 206376 56442 206428 56448
rect 206284 17264 206336 17270
rect 206284 17206 206336 17212
rect 200764 13116 200816 13122
rect 200764 13058 200816 13064
rect 198004 10328 198056 10334
rect 198004 10270 198056 10276
rect 196624 8968 196676 8974
rect 196624 8910 196676 8916
rect 206388 6186 206416 56442
rect 208412 32434 208440 92806
rect 209240 88097 209268 92820
rect 209806 92806 210280 92834
rect 209226 88088 209282 88097
rect 209226 88023 209282 88032
rect 210252 85377 210280 92806
rect 210344 86737 210372 92820
rect 211080 89457 211108 92820
rect 212198 92806 212488 92834
rect 212934 92806 213224 92834
rect 212460 91050 212488 92806
rect 213196 92410 213224 92806
rect 213184 92404 213236 92410
rect 213184 92346 213236 92352
rect 212448 91044 212500 91050
rect 212448 90986 212500 90992
rect 210514 89448 210570 89457
rect 210514 89383 210570 89392
rect 211066 89448 211122 89457
rect 211066 89383 211122 89392
rect 210330 86728 210386 86737
rect 210330 86663 210386 86672
rect 210238 85368 210294 85377
rect 210238 85303 210294 85312
rect 210252 84194 210280 85303
rect 210252 84166 210464 84194
rect 210436 56574 210464 84166
rect 210528 80714 210556 89383
rect 212460 82113 212488 90986
rect 212446 82104 212502 82113
rect 212446 82039 212502 82048
rect 210516 80708 210568 80714
rect 210516 80650 210568 80656
rect 213196 59362 213224 92346
rect 213472 90370 213500 92820
rect 213932 92806 214038 92834
rect 213460 90364 213512 90370
rect 213460 90306 213512 90312
rect 213472 88330 213500 90306
rect 213460 88324 213512 88330
rect 213460 88266 213512 88272
rect 213932 84114 213960 92806
rect 214576 88330 214604 92820
rect 215326 92806 215432 92834
rect 215298 90264 215354 90273
rect 215298 90199 215354 90208
rect 214564 88324 214616 88330
rect 214564 88266 214616 88272
rect 213920 84108 213972 84114
rect 213920 84050 213972 84056
rect 215312 66162 215340 90199
rect 215404 85542 215432 92806
rect 215864 88262 215892 92820
rect 216416 90273 216444 92820
rect 216692 92806 217166 92834
rect 216402 90264 216458 90273
rect 216402 90199 216458 90208
rect 215852 88256 215904 88262
rect 215852 88198 215904 88204
rect 216036 88256 216088 88262
rect 216036 88198 216088 88204
rect 215392 85536 215444 85542
rect 215392 85478 215444 85484
rect 215300 66156 215352 66162
rect 215300 66098 215352 66104
rect 215944 66156 215996 66162
rect 215944 66098 215996 66104
rect 215206 62792 215262 62801
rect 215206 62727 215262 62736
rect 215220 62558 215248 62727
rect 215208 62552 215260 62558
rect 215208 62494 215260 62500
rect 213184 59356 213236 59362
rect 213184 59298 213236 59304
rect 210424 56568 210476 56574
rect 210424 56510 210476 56516
rect 210436 43450 210464 56510
rect 210424 43444 210476 43450
rect 210424 43386 210476 43392
rect 213196 40730 213224 59298
rect 213184 40724 213236 40730
rect 213184 40666 213236 40672
rect 208400 32428 208452 32434
rect 208400 32370 208452 32376
rect 215220 18630 215248 62494
rect 215956 31074 215984 66098
rect 216048 62558 216076 88198
rect 216692 84182 216720 92806
rect 217704 89690 217732 92820
rect 217692 89684 217744 89690
rect 217692 89626 217744 89632
rect 218256 86970 218284 92820
rect 218808 92546 218836 92820
rect 218796 92540 218848 92546
rect 218796 92482 218848 92488
rect 218808 90953 218836 92482
rect 218794 90944 218850 90953
rect 218794 90879 218850 90888
rect 219544 86970 219572 92820
rect 219636 92806 220110 92834
rect 218244 86964 218296 86970
rect 218244 86906 218296 86912
rect 219532 86964 219584 86970
rect 219532 86906 219584 86912
rect 216680 84176 216732 84182
rect 216680 84118 216732 84124
rect 216692 82890 216720 84118
rect 216680 82884 216732 82890
rect 216680 82826 216732 82832
rect 217324 82884 217376 82890
rect 217324 82826 217376 82832
rect 216036 62552 216088 62558
rect 216036 62494 216088 62500
rect 217336 60722 217364 82826
rect 219636 81433 219664 92806
rect 220648 89690 220676 92820
rect 221384 91050 221412 92820
rect 221936 92546 221964 92820
rect 222212 92806 222502 92834
rect 222580 92806 223054 92834
rect 223790 92820 224038 92834
rect 223776 92806 224038 92820
rect 221924 92540 221976 92546
rect 221924 92482 221976 92488
rect 221372 91044 221424 91050
rect 221372 90986 221424 90992
rect 220636 89684 220688 89690
rect 220636 89626 220688 89632
rect 220084 86964 220136 86970
rect 220084 86906 220136 86912
rect 219622 81424 219678 81433
rect 219622 81359 219678 81368
rect 220096 75857 220124 86906
rect 220082 75848 220138 75857
rect 220082 75783 220138 75792
rect 220084 65544 220136 65550
rect 220084 65486 220136 65492
rect 217324 60716 217376 60722
rect 217324 60658 217376 60664
rect 217336 46238 217364 60658
rect 217324 46232 217376 46238
rect 217324 46174 217376 46180
rect 215944 31068 215996 31074
rect 215944 31010 215996 31016
rect 215208 18624 215260 18630
rect 215208 18566 215260 18572
rect 206376 6180 206428 6186
rect 206376 6122 206428 6128
rect 220096 4826 220124 65486
rect 222212 62082 222240 92806
rect 222580 84194 222608 92806
rect 223776 90302 223804 92806
rect 224038 92783 224094 92792
rect 224328 90681 224356 92820
rect 224314 90672 224370 90681
rect 224314 90607 224370 90616
rect 223764 90296 223816 90302
rect 223764 90238 223816 90244
rect 224868 90296 224920 90302
rect 224868 90238 224920 90244
rect 222304 84166 222608 84194
rect 222304 83094 222332 84166
rect 222292 83088 222344 83094
rect 222292 83030 222344 83036
rect 222844 83088 222896 83094
rect 222844 83030 222896 83036
rect 222856 82890 222884 83030
rect 222844 82884 222896 82890
rect 222844 82826 222896 82832
rect 222856 69018 222884 82826
rect 222844 69012 222896 69018
rect 222844 68954 222896 68960
rect 222200 62076 222252 62082
rect 222200 62018 222252 62024
rect 222212 60790 222240 62018
rect 222200 60784 222252 60790
rect 222200 60726 222252 60732
rect 222844 60784 222896 60790
rect 222844 60726 222896 60732
rect 222856 14550 222884 60726
rect 222844 14544 222896 14550
rect 222844 14486 222896 14492
rect 224880 7614 224908 90238
rect 224972 80034 225000 104910
rect 225050 104887 225106 104896
rect 225156 103514 225184 109647
rect 225064 103486 225184 103514
rect 224960 80028 225012 80034
rect 224960 79970 225012 79976
rect 225064 78674 225092 103486
rect 225142 97200 225198 97209
rect 225142 97135 225198 97144
rect 225156 92313 225184 97135
rect 225142 92304 225198 92313
rect 225142 92239 225198 92248
rect 225616 90953 225644 109686
rect 226524 108996 226576 109002
rect 226524 108938 226576 108944
rect 226536 107817 226564 108938
rect 226522 107808 226578 107817
rect 226522 107743 226578 107752
rect 226522 104272 226578 104281
rect 226522 104207 226578 104216
rect 226536 103562 226564 104207
rect 226524 103556 226576 103562
rect 226524 103498 226576 103504
rect 226340 102128 226392 102134
rect 226340 102070 226392 102076
rect 226352 101561 226380 102070
rect 226338 101552 226394 101561
rect 226338 101487 226394 101496
rect 226338 100736 226394 100745
rect 226338 100671 226394 100680
rect 226352 99226 226380 100671
rect 226430 99648 226486 99657
rect 226430 99583 226486 99592
rect 226444 99414 226472 99583
rect 226432 99408 226484 99414
rect 226432 99350 226484 99356
rect 226352 99198 226472 99226
rect 226338 98832 226394 98841
rect 226338 98767 226394 98776
rect 225602 90944 225658 90953
rect 225602 90879 225658 90888
rect 226352 82793 226380 98767
rect 226338 82784 226394 82793
rect 226338 82719 226394 82728
rect 225052 78668 225104 78674
rect 225052 78610 225104 78616
rect 226444 71738 226472 99198
rect 226524 98660 226576 98666
rect 226524 98602 226576 98608
rect 226536 96121 226564 98602
rect 226522 96112 226578 96121
rect 226522 96047 226578 96056
rect 226524 96008 226576 96014
rect 226524 95950 226576 95956
rect 226536 95305 226564 95950
rect 226522 95296 226578 95305
rect 226522 95231 226578 95240
rect 226536 88233 226564 95231
rect 226628 94489 226656 189722
rect 227732 178702 227760 241590
rect 230768 240106 230796 241604
rect 230756 240100 230808 240106
rect 230756 240042 230808 240048
rect 231122 236736 231178 236745
rect 231122 236671 231178 236680
rect 228362 230072 228418 230081
rect 228362 230007 228418 230016
rect 228376 192506 228404 230007
rect 228364 192500 228416 192506
rect 228364 192442 228416 192448
rect 228364 186992 228416 186998
rect 228364 186934 228416 186940
rect 227720 178696 227772 178702
rect 227720 178638 227772 178644
rect 227996 173188 228048 173194
rect 227996 173130 228048 173136
rect 228008 168502 228036 173130
rect 227996 168496 228048 168502
rect 227996 168438 228048 168444
rect 227718 160168 227774 160177
rect 227718 160103 227774 160112
rect 226708 137964 226760 137970
rect 226708 137906 226760 137912
rect 226720 137193 226748 137906
rect 226706 137184 226762 137193
rect 226706 137119 226762 137128
rect 226708 136332 226760 136338
rect 226708 136274 226760 136280
rect 226720 135561 226748 136274
rect 226706 135552 226762 135561
rect 226706 135487 226762 135496
rect 226706 134736 226762 134745
rect 226706 134671 226762 134680
rect 226720 133958 226748 134671
rect 226708 133952 226760 133958
rect 226708 133894 226760 133900
rect 226708 133816 226760 133822
rect 226708 133758 226760 133764
rect 226720 133657 226748 133758
rect 226706 133648 226762 133657
rect 226706 133583 226762 133592
rect 226708 133544 226760 133550
rect 226708 133486 226760 133492
rect 226720 132494 226748 133486
rect 226720 132466 226932 132494
rect 226708 131096 226760 131102
rect 226708 131038 226760 131044
rect 226720 130937 226748 131038
rect 226800 131028 226852 131034
rect 226800 130970 226852 130976
rect 226706 130928 226762 130937
rect 226706 130863 226762 130872
rect 226812 130121 226840 130970
rect 226798 130112 226854 130121
rect 226798 130047 226854 130056
rect 226708 129056 226760 129062
rect 226708 128998 226760 129004
rect 226720 128489 226748 128998
rect 226706 128480 226762 128489
rect 226706 128415 226762 128424
rect 226904 127702 226932 132466
rect 226708 127696 226760 127702
rect 226708 127638 226760 127644
rect 226892 127696 226944 127702
rect 226892 127638 226944 127644
rect 226720 127401 226748 127638
rect 226706 127392 226762 127401
rect 226706 127327 226762 127336
rect 227732 125769 227760 160103
rect 227812 146396 227864 146402
rect 227812 146338 227864 146344
rect 227718 125760 227774 125769
rect 227718 125695 227774 125704
rect 226706 117600 226762 117609
rect 226706 117535 226762 117544
rect 226720 117366 226748 117535
rect 226708 117360 226760 117366
rect 226708 117302 226760 117308
rect 226708 116000 226760 116006
rect 226706 115968 226708 115977
rect 226760 115968 226762 115977
rect 226706 115903 226762 115912
rect 227626 113792 227682 113801
rect 227824 113778 227852 146338
rect 227904 141432 227956 141438
rect 227904 141374 227956 141380
rect 227916 116793 227944 141374
rect 228008 139913 228036 168438
rect 228376 160177 228404 186934
rect 229098 165744 229154 165753
rect 229098 165679 229154 165688
rect 228362 160168 228418 160177
rect 228362 160103 228418 160112
rect 227994 139904 228050 139913
rect 227994 139839 228050 139848
rect 227994 129296 228050 129305
rect 227994 129231 228050 129240
rect 228008 127634 228036 129231
rect 227996 127628 228048 127634
rect 227996 127570 228048 127576
rect 229112 124166 229140 165679
rect 230018 150512 230074 150521
rect 230018 150447 230074 150456
rect 230032 149054 230060 150447
rect 230020 149048 230072 149054
rect 230020 148990 230072 148996
rect 229742 144936 229798 144945
rect 229742 144871 229798 144880
rect 229756 129742 229784 144871
rect 230032 142154 230060 148990
rect 230478 146568 230534 146577
rect 230478 146503 230534 146512
rect 229848 142126 230060 142154
rect 229848 136338 229876 142126
rect 229836 136332 229888 136338
rect 229836 136274 229888 136280
rect 230492 131102 230520 146503
rect 230480 131096 230532 131102
rect 230480 131038 230532 131044
rect 229744 129736 229796 129742
rect 229744 129678 229796 129684
rect 229756 124778 229784 129678
rect 229744 124772 229796 124778
rect 229744 124714 229796 124720
rect 229100 124160 229152 124166
rect 229100 124102 229152 124108
rect 228364 123480 228416 123486
rect 228364 123422 228416 123428
rect 227902 116784 227958 116793
rect 227902 116719 227958 116728
rect 227682 113750 227852 113778
rect 227626 113727 227682 113736
rect 226708 113144 226760 113150
rect 226708 113086 226760 113092
rect 226720 112169 226748 113086
rect 226706 112160 226762 112169
rect 226706 112095 226762 112104
rect 226984 109812 227036 109818
rect 226984 109754 227036 109760
rect 226708 107636 226760 107642
rect 226708 107578 226760 107584
rect 226720 107001 226748 107578
rect 226706 106992 226762 107001
rect 226706 106927 226762 106936
rect 226706 105904 226762 105913
rect 226706 105839 226762 105848
rect 226720 104922 226748 105839
rect 226708 104916 226760 104922
rect 226708 104858 226760 104864
rect 226706 103456 226762 103465
rect 226706 103391 226762 103400
rect 226720 102814 226748 103391
rect 226708 102808 226760 102814
rect 226708 102750 226760 102756
rect 226706 102368 226762 102377
rect 226706 102303 226762 102312
rect 226720 102202 226748 102303
rect 226708 102196 226760 102202
rect 226708 102138 226760 102144
rect 226996 98841 227024 109754
rect 227074 108624 227130 108633
rect 227074 108559 227130 108568
rect 227088 108322 227116 108559
rect 227076 108316 227128 108322
rect 227076 108258 227128 108264
rect 227720 108316 227772 108322
rect 227720 108258 227772 108264
rect 226982 98832 227038 98841
rect 226982 98767 227038 98776
rect 227628 94512 227680 94518
rect 226614 94480 226670 94489
rect 227628 94454 227680 94460
rect 226614 94415 226616 94424
rect 226668 94415 226670 94424
rect 226616 94386 226668 94392
rect 226628 94355 226656 94386
rect 227640 93673 227668 94454
rect 227626 93664 227682 93673
rect 227626 93599 227682 93608
rect 226522 88224 226578 88233
rect 226522 88159 226578 88168
rect 227732 86902 227760 108258
rect 227812 102808 227864 102814
rect 227812 102750 227864 102756
rect 227720 86896 227772 86902
rect 227720 86838 227772 86844
rect 227824 82822 227852 102750
rect 227902 98696 227958 98705
rect 227902 98631 227958 98640
rect 227916 98025 227944 98631
rect 227902 98016 227958 98025
rect 227902 97951 227958 97960
rect 227916 89593 227944 97951
rect 228376 96014 228404 123422
rect 230480 116000 230532 116006
rect 230480 115942 230532 115948
rect 229100 111172 229152 111178
rect 229100 111114 229152 111120
rect 228364 96008 228416 96014
rect 228364 95950 228416 95956
rect 228364 94444 228416 94450
rect 228364 94386 228416 94392
rect 227902 89584 227958 89593
rect 227902 89519 227958 89528
rect 228376 86290 228404 94386
rect 228364 86284 228416 86290
rect 228364 86226 228416 86232
rect 228362 83464 228418 83473
rect 228362 83399 228418 83408
rect 227812 82816 227864 82822
rect 227812 82758 227864 82764
rect 226432 71732 226484 71738
rect 226432 71674 226484 71680
rect 226444 70446 226472 71674
rect 226432 70440 226484 70446
rect 226432 70382 226484 70388
rect 226984 70440 227036 70446
rect 226984 70382 227036 70388
rect 226996 28286 227024 70382
rect 226984 28280 227036 28286
rect 226984 28222 227036 28228
rect 224868 7608 224920 7614
rect 224868 7550 224920 7556
rect 220084 4820 220136 4826
rect 220084 4762 220136 4768
rect 228376 4146 228404 83399
rect 229112 75886 229140 111114
rect 229192 99408 229244 99414
rect 229192 99350 229244 99356
rect 229204 92478 229232 99350
rect 229192 92472 229244 92478
rect 229192 92414 229244 92420
rect 229100 75880 229152 75886
rect 229100 75822 229152 75828
rect 230492 67522 230520 115942
rect 230480 67516 230532 67522
rect 230480 67458 230532 67464
rect 231136 14482 231164 236671
rect 231950 229800 232006 229809
rect 231950 229735 232006 229744
rect 231858 222048 231914 222057
rect 231858 221983 231914 221992
rect 231214 142352 231270 142361
rect 231214 142287 231270 142296
rect 231228 131782 231256 142287
rect 231216 131776 231268 131782
rect 231216 131718 231268 131724
rect 231768 116612 231820 116618
rect 231768 116554 231820 116560
rect 231780 116006 231808 116554
rect 231768 116000 231820 116006
rect 231768 115942 231820 115948
rect 231308 93152 231360 93158
rect 231308 93094 231360 93100
rect 231320 85377 231348 93094
rect 231872 92857 231900 221983
rect 231964 162897 231992 229735
rect 233160 222057 233188 241604
rect 235552 241369 235580 241604
rect 234618 241360 234674 241369
rect 234618 241295 234674 241304
rect 235538 241360 235594 241369
rect 235538 241295 235594 241304
rect 233146 222048 233202 222057
rect 233146 221983 233202 221992
rect 233882 213208 233938 213217
rect 233882 213143 233938 213152
rect 233240 167068 233292 167074
rect 233240 167010 233292 167016
rect 231950 162888 232006 162897
rect 231950 162823 232006 162832
rect 231964 132462 231992 162823
rect 231952 132456 232004 132462
rect 231952 132398 232004 132404
rect 232504 124908 232556 124914
rect 232504 124850 232556 124856
rect 231952 103556 232004 103562
rect 231952 103498 232004 103504
rect 231858 92848 231914 92857
rect 231858 92783 231914 92792
rect 231306 85368 231362 85377
rect 231306 85303 231362 85312
rect 231964 81394 231992 103498
rect 232516 92546 232544 124850
rect 233252 113150 233280 167010
rect 233330 153776 233386 153785
rect 233330 153711 233386 153720
rect 233344 138961 233372 153711
rect 233330 138952 233386 138961
rect 233330 138887 233386 138896
rect 233344 138689 233372 138887
rect 233330 138680 233386 138689
rect 233330 138615 233386 138624
rect 233896 133822 233924 213143
rect 234632 187066 234660 241295
rect 237656 240100 237708 240106
rect 237656 240042 237708 240048
rect 237380 239420 237432 239426
rect 237380 239362 237432 239368
rect 237392 235793 237420 239362
rect 237472 236020 237524 236026
rect 237472 235962 237524 235968
rect 237378 235784 237434 235793
rect 237378 235719 237434 235728
rect 235264 231124 235316 231130
rect 235264 231066 235316 231072
rect 234620 187060 234672 187066
rect 234620 187002 234672 187008
rect 234620 160744 234672 160750
rect 234620 160686 234672 160692
rect 234632 158817 234660 160686
rect 234618 158808 234674 158817
rect 234618 158743 234674 158752
rect 234632 141409 234660 158743
rect 234618 141400 234674 141409
rect 234618 141335 234674 141344
rect 233884 133816 233936 133822
rect 233884 133758 233936 133764
rect 233884 117428 233936 117434
rect 233884 117370 233936 117376
rect 233896 117201 233924 117370
rect 233882 117192 233938 117201
rect 233882 117127 233938 117136
rect 233332 115252 233384 115258
rect 233332 115194 233384 115200
rect 233344 114578 233372 115194
rect 233332 114572 233384 114578
rect 233332 114514 233384 114520
rect 233240 113144 233292 113150
rect 233240 113086 233292 113092
rect 233252 112470 233280 113086
rect 233240 112464 233292 112470
rect 233240 112406 233292 112412
rect 232504 92540 232556 92546
rect 232504 92482 232556 92488
rect 231952 81388 232004 81394
rect 231952 81330 232004 81336
rect 233344 70310 233372 114514
rect 233332 70304 233384 70310
rect 233332 70246 233384 70252
rect 233896 68950 233924 117127
rect 235276 90370 235304 231066
rect 235998 228304 236054 228313
rect 235998 228239 236054 228248
rect 236012 111178 236040 228239
rect 236642 226944 236698 226953
rect 236642 226879 236698 226888
rect 236656 206961 236684 226879
rect 236642 206952 236698 206961
rect 236642 206887 236698 206896
rect 236656 162761 236684 206887
rect 236090 162752 236146 162761
rect 236090 162687 236146 162696
rect 236642 162752 236698 162761
rect 236642 162687 236698 162696
rect 236104 161537 236132 162687
rect 236090 161528 236146 161537
rect 236090 161463 236146 161472
rect 236104 139398 236132 161463
rect 237380 153876 237432 153882
rect 237380 153818 237432 153824
rect 237392 153134 237420 153818
rect 237380 153128 237432 153134
rect 237380 153070 237432 153076
rect 236092 139392 236144 139398
rect 236092 139334 236144 139340
rect 236000 111172 236052 111178
rect 236000 111114 236052 111120
rect 237484 103514 237512 235962
rect 237392 103486 237512 103514
rect 237392 98734 237420 103486
rect 237564 102196 237616 102202
rect 237564 102138 237616 102144
rect 237380 98728 237432 98734
rect 237378 98696 237380 98705
rect 237432 98696 237434 98705
rect 237378 98631 237434 98640
rect 235264 90364 235316 90370
rect 235264 90306 235316 90312
rect 233884 68944 233936 68950
rect 233884 68886 233936 68892
rect 235276 68338 235304 90306
rect 237576 77246 237604 102138
rect 237668 85513 237696 240042
rect 237944 237386 237972 241604
rect 240152 241590 240350 241618
rect 237932 237380 237984 237386
rect 237932 237322 237984 237328
rect 237944 236026 237972 237322
rect 237932 236020 237984 236026
rect 237932 235962 237984 235968
rect 239404 232552 239456 232558
rect 239404 232494 239456 232500
rect 239416 213926 239444 232494
rect 239404 213920 239456 213926
rect 239404 213862 239456 213868
rect 240046 149152 240102 149161
rect 240152 149138 240180 241590
rect 242728 238678 242756 241604
rect 243542 240952 243598 240961
rect 243542 240887 243598 240896
rect 242716 238672 242768 238678
rect 242716 238614 242768 238620
rect 242728 237454 242756 238614
rect 242256 237448 242308 237454
rect 242256 237390 242308 237396
rect 242716 237448 242768 237454
rect 242716 237390 242768 237396
rect 242164 236700 242216 236706
rect 242164 236642 242216 236648
rect 240232 180124 240284 180130
rect 240232 180066 240284 180072
rect 240102 149110 240180 149138
rect 240046 149087 240102 149096
rect 239402 148336 239458 148345
rect 239402 148271 239458 148280
rect 237654 85504 237710 85513
rect 237654 85439 237710 85448
rect 238482 85504 238538 85513
rect 238482 85439 238538 85448
rect 238496 84930 238524 85439
rect 238484 84924 238536 84930
rect 238484 84866 238536 84872
rect 237564 77240 237616 77246
rect 237564 77182 237616 77188
rect 238024 77240 238076 77246
rect 238024 77182 238076 77188
rect 235264 68332 235316 68338
rect 235264 68274 235316 68280
rect 233884 60036 233936 60042
rect 233884 59978 233936 59984
rect 233896 17338 233924 59978
rect 233884 17332 233936 17338
rect 233884 17274 233936 17280
rect 233976 17264 234028 17270
rect 233976 17206 234028 17212
rect 231124 14476 231176 14482
rect 231124 14418 231176 14424
rect 228364 4140 228416 4146
rect 228364 4082 228416 4088
rect 233988 3466 234016 17206
rect 238036 4418 238064 77182
rect 239416 51746 239444 148271
rect 240060 135930 240088 149087
rect 240244 142154 240272 180066
rect 240322 156632 240378 156641
rect 240322 156567 240378 156576
rect 240152 142126 240272 142154
rect 240152 137970 240180 142126
rect 240140 137964 240192 137970
rect 240140 137906 240192 137912
rect 240048 135924 240100 135930
rect 240048 135866 240100 135872
rect 240336 131034 240364 156567
rect 240784 142180 240836 142186
rect 240784 142122 240836 142128
rect 240324 131028 240376 131034
rect 240324 130970 240376 130976
rect 240140 77988 240192 77994
rect 240140 77930 240192 77936
rect 239404 51740 239456 51746
rect 239404 51682 239456 51688
rect 238024 4412 238076 4418
rect 238024 4354 238076 4360
rect 239312 4412 239364 4418
rect 239312 4354 239364 4360
rect 184204 3460 184256 3466
rect 184204 3402 184256 3408
rect 233976 3460 234028 3466
rect 233976 3402 234028 3408
rect 239324 480 239352 4354
rect 240152 490 240180 77930
rect 240796 61402 240824 142122
rect 241428 137964 241480 137970
rect 241428 137906 241480 137912
rect 241440 137290 241468 137906
rect 241428 137284 241480 137290
rect 241428 137226 241480 137232
rect 240876 120760 240928 120766
rect 240876 120702 240928 120708
rect 240888 90681 240916 120702
rect 240874 90672 240930 90681
rect 240874 90607 240930 90616
rect 242176 88262 242204 236642
rect 242268 92410 242296 237390
rect 243556 185638 243584 240887
rect 244924 240780 244976 240786
rect 244924 240722 244976 240728
rect 244280 225684 244332 225690
rect 244280 225626 244332 225632
rect 244292 224942 244320 225626
rect 244280 224936 244332 224942
rect 244280 224878 244332 224884
rect 243544 185632 243596 185638
rect 243544 185574 243596 185580
rect 243544 178356 243596 178362
rect 243544 178298 243596 178304
rect 243556 159526 243584 178298
rect 242900 159520 242952 159526
rect 242900 159462 242952 159468
rect 243544 159520 243596 159526
rect 243544 159462 243596 159468
rect 242912 159390 242940 159462
rect 242900 159384 242952 159390
rect 242900 159326 242952 159332
rect 242912 126954 242940 159326
rect 244370 153096 244426 153105
rect 244370 153031 244426 153040
rect 244384 151881 244412 153031
rect 244370 151872 244426 151881
rect 244370 151807 244426 151816
rect 242900 126948 242952 126954
rect 242900 126890 242952 126896
rect 243360 126948 243412 126954
rect 243360 126890 243412 126896
rect 243372 126274 243400 126890
rect 243360 126268 243412 126274
rect 243360 126210 243412 126216
rect 244384 121446 244412 151807
rect 244372 121440 244424 121446
rect 244372 121382 244424 121388
rect 244280 117360 244332 117366
rect 244280 117302 244332 117308
rect 242256 92404 242308 92410
rect 242256 92346 242308 92352
rect 242164 88256 242216 88262
rect 242164 88198 242216 88204
rect 241520 86284 241572 86290
rect 241520 86226 241572 86232
rect 241532 64870 241560 86226
rect 244292 77178 244320 117302
rect 244280 77172 244332 77178
rect 244280 77114 244332 77120
rect 244292 76362 244320 77114
rect 244280 76356 244332 76362
rect 244280 76298 244332 76304
rect 244936 75818 244964 240722
rect 245016 224936 245068 224942
rect 245016 224878 245068 224884
rect 245028 153105 245056 224878
rect 245014 153096 245070 153105
rect 245014 153031 245070 153040
rect 245120 146305 245148 241604
rect 246302 239592 246358 239601
rect 246302 239527 246358 239536
rect 245660 225616 245712 225622
rect 245660 225558 245712 225564
rect 245106 146296 245162 146305
rect 245106 146231 245162 146240
rect 245672 109002 245700 225558
rect 246316 218006 246344 239527
rect 247512 239465 247540 241604
rect 247498 239456 247554 239465
rect 247498 239391 247554 239400
rect 247040 238808 247092 238814
rect 247040 238750 247092 238756
rect 247052 234433 247080 238750
rect 247038 234424 247094 234433
rect 247038 234359 247094 234368
rect 248326 228440 248382 228449
rect 248326 228375 248382 228384
rect 248340 224913 248368 228375
rect 248326 224904 248382 224913
rect 248326 224839 248382 224848
rect 249062 224904 249118 224913
rect 249062 224839 249118 224848
rect 246304 218000 246356 218006
rect 246304 217942 246356 217948
rect 245660 108996 245712 109002
rect 245660 108938 245712 108944
rect 246316 89758 246344 217942
rect 247040 217320 247092 217326
rect 247038 217288 247040 217297
rect 247092 217288 247094 217297
rect 247038 217223 247094 217232
rect 248326 217288 248382 217297
rect 248326 217223 248382 217232
rect 248340 178702 248368 217223
rect 249076 180794 249104 224839
rect 248984 180766 249104 180794
rect 247684 178696 247736 178702
rect 247684 178638 247736 178644
rect 248328 178696 248380 178702
rect 248328 178638 248380 178644
rect 247696 156466 247724 178638
rect 248984 175302 249012 180766
rect 248972 175296 249024 175302
rect 248972 175238 249024 175244
rect 248984 174593 249012 175238
rect 248970 174584 249026 174593
rect 248970 174519 249026 174528
rect 249064 159384 249116 159390
rect 249064 159326 249116 159332
rect 247040 156460 247092 156466
rect 247040 156402 247092 156408
rect 247684 156460 247736 156466
rect 247684 156402 247736 156408
rect 247052 156058 247080 156402
rect 247040 156052 247092 156058
rect 247040 155994 247092 156000
rect 247052 122806 247080 155994
rect 247040 122800 247092 122806
rect 247040 122742 247092 122748
rect 245660 89752 245712 89758
rect 245660 89694 245712 89700
rect 246304 89752 246356 89758
rect 246304 89694 246356 89700
rect 245672 86970 245700 89694
rect 245660 86964 245712 86970
rect 245660 86906 245712 86912
rect 245660 82136 245712 82142
rect 245660 82078 245712 82084
rect 245016 76356 245068 76362
rect 245016 76298 245068 76304
rect 244924 75812 244976 75818
rect 244924 75754 244976 75760
rect 241520 64864 241572 64870
rect 241520 64806 241572 64812
rect 240784 61396 240836 61402
rect 240784 61338 240836 61344
rect 241532 16574 241560 64806
rect 244280 57248 244332 57254
rect 244280 57190 244332 57196
rect 241532 16546 241744 16574
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 16546
rect 244292 6914 244320 57190
rect 245028 15910 245056 76298
rect 245672 16574 245700 82078
rect 245672 16546 245976 16574
rect 245016 15904 245068 15910
rect 245016 15846 245068 15852
rect 244292 6886 245240 6914
rect 244096 4820 244148 4826
rect 244096 4762 244148 4768
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244108 480 244136 4762
rect 245212 480 245240 6886
rect 245948 490 245976 16546
rect 247592 6180 247644 6186
rect 247592 6122 247644 6128
rect 246224 598 246436 626
rect 246224 490 246252 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 462 246252 490
rect 246408 480 246436 598
rect 247604 480 247632 6122
rect 249076 4146 249104 159326
rect 249168 93158 249196 242014
rect 249812 211138 249840 242014
rect 249918 242012 250166 242026
rect 249904 241998 250166 242012
rect 249800 211132 249852 211138
rect 249800 211074 249852 211080
rect 249156 93152 249208 93158
rect 249156 93094 249208 93100
rect 249812 73166 249840 211074
rect 249904 178362 249932 241998
rect 250166 241975 250222 241984
rect 252296 240106 252324 241604
rect 251824 240100 251876 240106
rect 251824 240042 251876 240048
rect 252284 240100 252336 240106
rect 252284 240042 252336 240048
rect 251836 239873 251864 240042
rect 251822 239864 251878 239873
rect 251822 239799 251878 239808
rect 250534 239456 250590 239465
rect 250534 239391 250590 239400
rect 250442 235240 250498 235249
rect 250442 235175 250498 235184
rect 249892 178356 249944 178362
rect 249892 178298 249944 178304
rect 250456 92449 250484 235175
rect 250548 211041 250576 239391
rect 250534 211032 250590 211041
rect 250534 210967 250590 210976
rect 251836 173194 251864 239799
rect 252466 239728 252522 239737
rect 252466 239663 252522 239672
rect 252480 238814 252508 239663
rect 252468 238808 252520 238814
rect 252468 238750 252520 238756
rect 251916 192568 251968 192574
rect 251916 192510 251968 192516
rect 251824 173188 251876 173194
rect 251824 173130 251876 173136
rect 251928 140758 251956 192510
rect 251916 140752 251968 140758
rect 251916 140694 251968 140700
rect 251928 139466 251956 140694
rect 251180 139460 251232 139466
rect 251180 139402 251232 139408
rect 251916 139460 251968 139466
rect 251916 139402 251968 139408
rect 250536 98728 250588 98734
rect 250536 98670 250588 98676
rect 250548 93158 250576 98670
rect 250536 93152 250588 93158
rect 250536 93094 250588 93100
rect 250442 92440 250498 92449
rect 250442 92375 250498 92384
rect 249800 73160 249852 73166
rect 249800 73102 249852 73108
rect 249800 62824 249852 62830
rect 249800 62766 249852 62772
rect 249812 16574 249840 62766
rect 249812 16546 250024 16574
rect 248788 4140 248840 4146
rect 248788 4082 248840 4088
rect 249064 4140 249116 4146
rect 249064 4082 249116 4088
rect 248800 480 248828 4082
rect 249996 480 250024 16546
rect 251192 3602 251220 139402
rect 252572 109750 252600 307022
rect 252756 298058 252784 308382
rect 253202 303648 253258 303657
rect 253202 303583 253258 303592
rect 252926 301608 252982 301617
rect 253216 301594 253244 303583
rect 252982 301580 253244 301594
rect 252982 301566 253230 301580
rect 252926 301543 252982 301552
rect 252836 300892 252888 300898
rect 252836 300834 252888 300840
rect 252848 299033 252876 300834
rect 253308 299849 253336 325666
rect 254030 319424 254086 319433
rect 254030 319359 254086 319368
rect 253018 299840 253074 299849
rect 253018 299775 253074 299784
rect 253294 299840 253350 299849
rect 253294 299775 253350 299784
rect 252834 299024 252890 299033
rect 252834 298959 252890 298968
rect 252834 298072 252890 298081
rect 252756 298030 252834 298058
rect 252834 298007 252890 298016
rect 252834 293448 252890 293457
rect 252756 293406 252834 293434
rect 252756 235346 252784 293406
rect 252834 293383 252890 293392
rect 253032 291938 253060 299775
rect 253952 295662 253980 295693
rect 253940 295656 253992 295662
rect 253938 295624 253940 295633
rect 253992 295624 253994 295633
rect 253938 295559 253994 295568
rect 253202 292904 253258 292913
rect 253202 292839 253258 292848
rect 252848 291910 253060 291938
rect 252744 235340 252796 235346
rect 252744 235282 252796 235288
rect 252744 227792 252796 227798
rect 252744 227734 252796 227740
rect 252756 114481 252784 227734
rect 252848 154601 252876 291910
rect 253018 244488 253074 244497
rect 253018 244423 253074 244432
rect 252926 242856 252982 242865
rect 252926 242791 252982 242800
rect 252940 242049 252968 242791
rect 253032 242078 253060 244423
rect 253020 242072 253072 242078
rect 252926 242040 252982 242049
rect 253020 242014 253072 242020
rect 252926 241975 252982 241984
rect 253216 229022 253244 292839
rect 253204 229016 253256 229022
rect 253204 228958 253256 228964
rect 253216 227798 253244 228958
rect 253204 227792 253256 227798
rect 253204 227734 253256 227740
rect 253952 202162 253980 295559
rect 254044 254017 254072 319359
rect 254596 317393 254624 349862
rect 254582 317384 254638 317393
rect 254582 317319 254638 317328
rect 254122 315344 254178 315353
rect 254122 315279 254178 315288
rect 254030 254008 254086 254017
rect 254030 253943 254086 253952
rect 254030 251560 254086 251569
rect 254030 251495 254086 251504
rect 253940 202156 253992 202162
rect 253940 202098 253992 202104
rect 254044 168366 254072 251495
rect 254136 246401 254164 315279
rect 255320 309800 255372 309806
rect 255320 309742 255372 309748
rect 254214 302288 254270 302297
rect 254214 302223 254270 302232
rect 254228 249801 254256 302223
rect 255332 296177 255360 309742
rect 255318 296168 255374 296177
rect 255318 296103 255374 296112
rect 255332 295497 255360 296103
rect 255318 295488 255374 295497
rect 255318 295423 255374 295432
rect 255320 295316 255372 295322
rect 255320 295258 255372 295264
rect 255332 294409 255360 295258
rect 255318 294400 255374 294409
rect 255318 294335 255374 294344
rect 255424 294114 255452 369718
rect 255516 360194 255544 392090
rect 256712 389298 256740 393926
rect 256700 389292 256752 389298
rect 256700 389234 256752 389240
rect 256804 381546 256832 494770
rect 256976 451036 257028 451042
rect 256976 450978 257028 450984
rect 256882 440464 256938 440473
rect 256882 440399 256938 440408
rect 256896 394641 256924 440399
rect 256988 423434 257016 450978
rect 256976 423428 257028 423434
rect 256976 423370 257028 423376
rect 256882 394632 256938 394641
rect 256882 394567 256938 394576
rect 256792 381540 256844 381546
rect 256792 381482 256844 381488
rect 256792 365016 256844 365022
rect 256792 364958 256844 364964
rect 255504 360188 255556 360194
rect 255504 360130 255556 360136
rect 255516 359718 255544 360130
rect 255504 359712 255556 359718
rect 255504 359654 255556 359660
rect 255964 359712 256016 359718
rect 255964 359654 256016 359660
rect 255976 300898 256004 359654
rect 256700 326392 256752 326398
rect 256700 326334 256752 326340
rect 255596 300892 255648 300898
rect 255596 300834 255648 300840
rect 255964 300892 256016 300898
rect 255964 300834 256016 300840
rect 255502 300792 255558 300801
rect 255502 300727 255558 300736
rect 255516 300082 255544 300727
rect 255608 300393 255636 300834
rect 255594 300384 255650 300393
rect 255594 300319 255650 300328
rect 255504 300076 255556 300082
rect 255504 300018 255556 300024
rect 255504 299464 255556 299470
rect 255504 299406 255556 299412
rect 255516 299169 255544 299406
rect 255502 299160 255558 299169
rect 255502 299095 255558 299104
rect 255870 298752 255926 298761
rect 255870 298687 255926 298696
rect 255594 298616 255650 298625
rect 255594 298551 255650 298560
rect 255502 298208 255558 298217
rect 255502 298143 255504 298152
rect 255556 298143 255558 298152
rect 255504 298114 255556 298120
rect 255502 296984 255558 296993
rect 255502 296919 255558 296928
rect 255516 296818 255544 296919
rect 255504 296812 255556 296818
rect 255504 296754 255556 296760
rect 255504 296608 255556 296614
rect 255502 296576 255504 296585
rect 255556 296576 255558 296585
rect 255502 296511 255558 296520
rect 255332 294086 255452 294114
rect 255332 293185 255360 294086
rect 255412 294024 255464 294030
rect 255410 293992 255412 294001
rect 255464 293992 255466 294001
rect 255410 293927 255466 293936
rect 255412 293276 255464 293282
rect 255412 293218 255464 293224
rect 255318 293176 255374 293185
rect 255318 293111 255374 293120
rect 255424 292641 255452 293218
rect 255410 292632 255466 292641
rect 255410 292567 255466 292576
rect 255504 282872 255556 282878
rect 255504 282814 255556 282820
rect 255412 282804 255464 282810
rect 255412 282746 255464 282752
rect 255424 282033 255452 282746
rect 255516 282441 255544 282814
rect 255502 282432 255558 282441
rect 255502 282367 255558 282376
rect 255410 282024 255466 282033
rect 255410 281959 255466 281968
rect 255412 281512 255464 281518
rect 255410 281480 255412 281489
rect 255464 281480 255466 281489
rect 255410 281415 255466 281424
rect 255504 281444 255556 281450
rect 255504 281386 255556 281392
rect 255516 280265 255544 281386
rect 255502 280256 255558 280265
rect 255502 280191 255558 280200
rect 255412 279472 255464 279478
rect 255412 279414 255464 279420
rect 255424 279041 255452 279414
rect 255410 279032 255466 279041
rect 255410 278967 255466 278976
rect 255504 278724 255556 278730
rect 255504 278666 255556 278672
rect 255410 278488 255466 278497
rect 255410 278423 255466 278432
rect 255424 278050 255452 278423
rect 255412 278044 255464 278050
rect 255412 277986 255464 277992
rect 255516 277681 255544 278666
rect 255502 277672 255558 277681
rect 255502 277607 255558 277616
rect 255412 277364 255464 277370
rect 255412 277306 255464 277312
rect 255424 276457 255452 277306
rect 255502 277264 255558 277273
rect 255502 277199 255558 277208
rect 255410 276448 255466 276457
rect 255410 276383 255466 276392
rect 255516 276078 255544 277199
rect 255504 276072 255556 276078
rect 255504 276014 255556 276020
rect 255412 276004 255464 276010
rect 255412 275946 255464 275952
rect 255424 275097 255452 275946
rect 255504 275664 255556 275670
rect 255504 275606 255556 275612
rect 255516 275505 255544 275606
rect 255502 275496 255558 275505
rect 255502 275431 255558 275440
rect 255410 275088 255466 275097
rect 255410 275023 255466 275032
rect 255504 274644 255556 274650
rect 255504 274586 255556 274592
rect 255410 274272 255466 274281
rect 255410 274207 255466 274216
rect 255424 273970 255452 274207
rect 255412 273964 255464 273970
rect 255412 273906 255464 273912
rect 255516 273873 255544 274586
rect 255502 273864 255558 273873
rect 255502 273799 255558 273808
rect 255504 273216 255556 273222
rect 255410 273184 255466 273193
rect 255504 273158 255556 273164
rect 255410 273119 255466 273128
rect 255424 272105 255452 273119
rect 255516 272513 255544 273158
rect 255502 272504 255558 272513
rect 255502 272439 255558 272448
rect 255410 272096 255466 272105
rect 255410 272031 255466 272040
rect 255502 271824 255558 271833
rect 255502 271759 255558 271768
rect 255318 271688 255374 271697
rect 255318 271623 255374 271632
rect 255332 270609 255360 271623
rect 255410 271280 255466 271289
rect 255410 271215 255466 271224
rect 255424 270842 255452 271215
rect 255516 270881 255544 271759
rect 255502 270872 255558 270881
rect 255412 270836 255464 270842
rect 255502 270807 255558 270816
rect 255412 270778 255464 270784
rect 255318 270600 255374 270609
rect 255318 270535 255374 270544
rect 255412 270496 255464 270502
rect 255412 270438 255464 270444
rect 255424 269929 255452 270438
rect 255410 269920 255466 269929
rect 255410 269855 255466 269864
rect 255502 269104 255558 269113
rect 255502 269039 255558 269048
rect 255410 267880 255466 267889
rect 255410 267815 255412 267824
rect 255464 267815 255466 267824
rect 255412 267786 255464 267792
rect 255516 267782 255544 269039
rect 255504 267776 255556 267782
rect 255504 267718 255556 267724
rect 255412 267708 255464 267714
rect 255412 267650 255464 267656
rect 255424 267481 255452 267650
rect 255410 267472 255466 267481
rect 255410 267407 255466 267416
rect 255412 266212 255464 266218
rect 255412 266154 255464 266160
rect 255318 266112 255374 266121
rect 255318 266047 255374 266056
rect 255332 264994 255360 266047
rect 255424 265713 255452 266154
rect 255410 265704 255466 265713
rect 255410 265639 255466 265648
rect 255320 264988 255372 264994
rect 255320 264930 255372 264936
rect 255502 264344 255558 264353
rect 255502 264279 255558 264288
rect 255412 264172 255464 264178
rect 255412 264114 255464 264120
rect 255424 263945 255452 264114
rect 255410 263936 255466 263945
rect 255410 263871 255466 263880
rect 255516 263770 255544 264279
rect 255504 263764 255556 263770
rect 255504 263706 255556 263712
rect 255502 263120 255558 263129
rect 255502 263055 255558 263064
rect 255516 262342 255544 263055
rect 255504 262336 255556 262342
rect 255410 262304 255466 262313
rect 255504 262278 255556 262284
rect 255410 262239 255412 262248
rect 255464 262239 255466 262248
rect 255412 262210 255464 262216
rect 255410 261896 255466 261905
rect 255410 261831 255466 261840
rect 255424 261390 255452 261831
rect 255504 261520 255556 261526
rect 255504 261462 255556 261468
rect 255412 261384 255464 261390
rect 255412 261326 255464 261332
rect 255318 261080 255374 261089
rect 255318 261015 255374 261024
rect 255332 259729 255360 261015
rect 255516 260953 255544 261462
rect 255502 260944 255558 260953
rect 255502 260879 255558 260888
rect 255410 260536 255466 260545
rect 255410 260471 255412 260480
rect 255464 260471 255466 260480
rect 255412 260442 255464 260448
rect 255318 259720 255374 259729
rect 255318 259655 255374 259664
rect 255412 259412 255464 259418
rect 255412 259354 255464 259360
rect 255424 258369 255452 259354
rect 255410 258360 255466 258369
rect 255410 258295 255466 258304
rect 255412 258052 255464 258058
rect 255412 257994 255464 258000
rect 255318 257544 255374 257553
rect 255318 257479 255374 257488
rect 255332 257378 255360 257479
rect 255320 257372 255372 257378
rect 255320 257314 255372 257320
rect 255424 257145 255452 257994
rect 255410 257136 255466 257145
rect 255410 257071 255466 257080
rect 255502 256320 255558 256329
rect 255502 256255 255558 256264
rect 255516 255406 255544 256255
rect 255504 255400 255556 255406
rect 255410 255368 255466 255377
rect 255504 255342 255556 255348
rect 255410 255303 255412 255312
rect 255464 255303 255466 255312
rect 255412 255274 255464 255280
rect 255502 254960 255558 254969
rect 255502 254895 255558 254904
rect 255412 254584 255464 254590
rect 255410 254552 255412 254561
rect 255464 254552 255466 254561
rect 255410 254487 255466 254496
rect 255516 253978 255544 254895
rect 255504 253972 255556 253978
rect 255504 253914 255556 253920
rect 255502 253328 255558 253337
rect 255502 253263 255558 253272
rect 255410 252784 255466 252793
rect 255410 252719 255412 252728
rect 255464 252719 255466 252728
rect 255412 252690 255464 252696
rect 255516 252618 255544 253263
rect 255504 252612 255556 252618
rect 255504 252554 255556 252560
rect 254950 252512 255006 252521
rect 254950 252447 255006 252456
rect 254964 251569 254992 252447
rect 255410 251968 255466 251977
rect 255410 251903 255466 251912
rect 255424 251870 255452 251903
rect 255412 251864 255464 251870
rect 255412 251806 255464 251812
rect 254950 251560 255006 251569
rect 254950 251495 255006 251504
rect 255320 251252 255372 251258
rect 255320 251194 255372 251200
rect 254214 249792 254270 249801
rect 254214 249727 254270 249736
rect 254228 249422 254256 249727
rect 254216 249416 254268 249422
rect 254216 249358 254268 249364
rect 255332 248577 255360 251194
rect 255502 251152 255558 251161
rect 255502 251087 255558 251096
rect 255412 250572 255464 250578
rect 255412 250514 255464 250520
rect 255424 250345 255452 250514
rect 255516 250510 255544 251087
rect 255504 250504 255556 250510
rect 255504 250446 255556 250452
rect 255410 250336 255466 250345
rect 255410 250271 255466 250280
rect 255502 249384 255558 249393
rect 255502 249319 255558 249328
rect 255410 248976 255466 248985
rect 255410 248911 255466 248920
rect 255318 248568 255374 248577
rect 255318 248503 255374 248512
rect 255424 248470 255452 248911
rect 255412 248464 255464 248470
rect 255516 248441 255544 249319
rect 255412 248406 255464 248412
rect 255502 248432 255558 248441
rect 255502 248367 255558 248376
rect 255502 248160 255558 248169
rect 255502 248095 255558 248104
rect 255410 247752 255466 247761
rect 255410 247687 255412 247696
rect 255464 247687 255466 247696
rect 255412 247658 255464 247664
rect 255516 247110 255544 248095
rect 255504 247104 255556 247110
rect 255504 247046 255556 247052
rect 255502 246800 255558 246809
rect 255502 246735 255558 246744
rect 254122 246392 254178 246401
rect 254122 246327 254178 246336
rect 255318 246392 255374 246401
rect 255318 246327 255374 246336
rect 254122 243808 254178 243817
rect 254122 243743 254178 243752
rect 254136 239601 254164 243743
rect 254214 242584 254270 242593
rect 254214 242519 254270 242528
rect 254122 239592 254178 239601
rect 254122 239527 254178 239536
rect 254228 237969 254256 242519
rect 255332 238754 255360 246327
rect 255516 245682 255544 246735
rect 255504 245676 255556 245682
rect 255504 245618 255556 245624
rect 255412 245608 255464 245614
rect 255410 245576 255412 245585
rect 255464 245576 255466 245585
rect 255410 245511 255466 245520
rect 255410 245168 255466 245177
rect 255410 245103 255466 245112
rect 255424 244322 255452 245103
rect 255412 244316 255464 244322
rect 255412 244258 255464 244264
rect 255502 244216 255558 244225
rect 255502 244151 255558 244160
rect 255516 243574 255544 244151
rect 255504 243568 255556 243574
rect 255504 243510 255556 243516
rect 255332 238726 255544 238754
rect 254214 237960 254270 237969
rect 254214 237895 254270 237904
rect 255516 235278 255544 238726
rect 255504 235272 255556 235278
rect 255504 235214 255556 235220
rect 255608 222902 255636 298551
rect 255884 297401 255912 298687
rect 256054 297800 256110 297809
rect 256054 297735 256110 297744
rect 255870 297392 255926 297401
rect 255870 297327 255926 297336
rect 256068 296750 256096 297735
rect 256056 296744 256108 296750
rect 256056 296686 256108 296692
rect 255686 295488 255742 295497
rect 255686 295423 255742 295432
rect 255700 231130 255728 295423
rect 256712 295089 256740 326334
rect 256804 325694 256832 364958
rect 257080 353977 257108 533287
rect 258092 507210 258120 568890
rect 258172 567316 258224 567322
rect 258172 567258 258224 567264
rect 258184 538354 258212 567258
rect 259368 561060 259420 561066
rect 259368 561002 259420 561008
rect 259380 552702 259408 561002
rect 259368 552696 259420 552702
rect 259368 552638 259420 552644
rect 258264 545284 258316 545290
rect 258264 545226 258316 545232
rect 258172 538348 258224 538354
rect 258172 538290 258224 538296
rect 258276 525065 258304 545226
rect 258262 525056 258318 525065
rect 258262 524991 258318 525000
rect 258172 521008 258224 521014
rect 258172 520950 258224 520956
rect 258080 507204 258132 507210
rect 258080 507146 258132 507152
rect 258184 480254 258212 520950
rect 258184 480226 258304 480254
rect 258276 476134 258304 480226
rect 258264 476128 258316 476134
rect 258264 476070 258316 476076
rect 258080 455456 258132 455462
rect 258080 455398 258132 455404
rect 257342 454064 257398 454073
rect 257342 453999 257398 454008
rect 257356 442338 257384 453999
rect 257344 442332 257396 442338
rect 257344 442274 257396 442280
rect 257066 353968 257122 353977
rect 257066 353903 257122 353912
rect 258092 338774 258120 455398
rect 258172 449948 258224 449954
rect 258172 449890 258224 449896
rect 258184 390833 258212 449890
rect 258276 443698 258304 476070
rect 258264 443692 258316 443698
rect 258264 443634 258316 443640
rect 258998 398576 259054 398585
rect 258998 398511 259054 398520
rect 258724 396772 258776 396778
rect 258724 396714 258776 396720
rect 258170 390824 258226 390833
rect 258170 390759 258226 390768
rect 258736 386306 258764 396714
rect 259012 395350 259040 398511
rect 259000 395344 259052 395350
rect 259000 395286 259052 395292
rect 259276 391332 259328 391338
rect 259276 391274 259328 391280
rect 258724 386300 258776 386306
rect 258724 386242 258776 386248
rect 259288 384849 259316 391274
rect 259274 384840 259330 384849
rect 259274 384775 259330 384784
rect 259472 351801 259500 601666
rect 262218 599040 262274 599049
rect 262218 598975 262274 598984
rect 261024 589348 261076 589354
rect 261024 589290 261076 589296
rect 259644 561740 259696 561746
rect 259644 561682 259696 561688
rect 259552 550724 259604 550730
rect 259552 550666 259604 550672
rect 259564 469198 259592 550666
rect 259656 533458 259684 561682
rect 260932 560312 260984 560318
rect 260932 560254 260984 560260
rect 260840 553512 260892 553518
rect 260840 553454 260892 553460
rect 259644 533452 259696 533458
rect 259644 533394 259696 533400
rect 259552 469192 259604 469198
rect 259552 469134 259604 469140
rect 259552 460216 259604 460222
rect 259552 460158 259604 460164
rect 259564 429554 259592 460158
rect 259642 458552 259698 458561
rect 259642 458487 259698 458496
rect 259656 442270 259684 458487
rect 260104 454028 260156 454034
rect 260104 453970 260156 453976
rect 260116 452674 260144 453970
rect 260104 452668 260156 452674
rect 260104 452610 260156 452616
rect 259644 442264 259696 442270
rect 259644 442206 259696 442212
rect 259552 429548 259604 429554
rect 259552 429490 259604 429496
rect 259552 401668 259604 401674
rect 259552 401610 259604 401616
rect 259564 383081 259592 401610
rect 259550 383072 259606 383081
rect 259550 383007 259606 383016
rect 259458 351792 259514 351801
rect 259458 351727 259514 351736
rect 259368 347744 259420 347750
rect 259368 347686 259420 347692
rect 258080 338768 258132 338774
rect 258080 338710 258132 338716
rect 256804 325666 256924 325694
rect 256896 311982 256924 325666
rect 258724 324352 258776 324358
rect 258724 324294 258776 324300
rect 256884 311976 256936 311982
rect 256884 311918 256936 311924
rect 256792 301572 256844 301578
rect 256792 301514 256844 301520
rect 256698 295080 256754 295089
rect 256698 295015 256754 295024
rect 256698 294808 256754 294817
rect 256698 294743 256754 294752
rect 256712 293350 256740 294743
rect 256804 293593 256832 301514
rect 256790 293584 256846 293593
rect 256790 293519 256846 293528
rect 256700 293344 256752 293350
rect 256700 293286 256752 293292
rect 256606 292224 256662 292233
rect 256662 292182 256832 292210
rect 256606 292159 256662 292168
rect 256608 291916 256660 291922
rect 256608 291858 256660 291864
rect 256620 291825 256648 291858
rect 256606 291816 256662 291825
rect 256662 291774 256740 291802
rect 256606 291751 256662 291760
rect 256516 291100 256568 291106
rect 256516 291042 256568 291048
rect 256528 291009 256556 291042
rect 256514 291000 256570 291009
rect 256514 290935 256570 290944
rect 256514 290592 256570 290601
rect 256514 290527 256570 290536
rect 256528 289882 256556 290527
rect 256516 289876 256568 289882
rect 256516 289818 256568 289824
rect 256608 289808 256660 289814
rect 256608 289750 256660 289756
rect 256514 289640 256570 289649
rect 256514 289575 256570 289584
rect 256528 289134 256556 289575
rect 256620 289241 256648 289750
rect 256606 289232 256662 289241
rect 256606 289167 256662 289176
rect 256516 289128 256568 289134
rect 256516 289070 256568 289076
rect 255872 288380 255924 288386
rect 255872 288322 255924 288328
rect 255884 288017 255912 288322
rect 255870 288008 255926 288017
rect 255870 287943 255926 287952
rect 255964 287768 256016 287774
rect 255964 287710 256016 287716
rect 255976 287609 256004 287710
rect 255962 287600 256018 287609
rect 255962 287535 256018 287544
rect 255872 287020 255924 287026
rect 255872 286962 255924 286968
rect 255884 286657 255912 286962
rect 255870 286648 255926 286657
rect 255870 286583 255926 286592
rect 256514 286240 256570 286249
rect 256514 286175 256570 286184
rect 256528 285734 256556 286175
rect 256516 285728 256568 285734
rect 256516 285670 256568 285676
rect 256608 285660 256660 285666
rect 256608 285602 256660 285608
rect 256620 285433 256648 285602
rect 256606 285424 256662 285433
rect 256606 285359 256662 285368
rect 256424 284300 256476 284306
rect 256424 284242 256476 284248
rect 255780 283892 255832 283898
rect 255780 283834 255832 283840
rect 255792 283665 255820 283834
rect 255778 283656 255834 283665
rect 255778 283591 255834 283600
rect 256436 283257 256464 284242
rect 256422 283248 256478 283257
rect 256422 283183 256478 283192
rect 255778 271144 255834 271153
rect 255778 271079 255834 271088
rect 255792 268297 255820 271079
rect 255778 268288 255834 268297
rect 255778 268223 255834 268232
rect 255872 244248 255924 244254
rect 255872 244190 255924 244196
rect 255884 243409 255912 244190
rect 255870 243400 255926 243409
rect 255870 243335 255926 243344
rect 255688 231124 255740 231130
rect 255688 231066 255740 231072
rect 255596 222896 255648 222902
rect 255596 222838 255648 222844
rect 256606 220144 256662 220153
rect 256606 220079 256662 220088
rect 256620 219337 256648 220079
rect 256606 219328 256662 219337
rect 256606 219263 256662 219272
rect 256056 216028 256108 216034
rect 256056 215970 256108 215976
rect 255228 198008 255280 198014
rect 255228 197950 255280 197956
rect 254032 168360 254084 168366
rect 254032 168302 254084 168308
rect 252834 154592 252890 154601
rect 252834 154527 252890 154536
rect 252848 145654 252876 154527
rect 252836 145648 252888 145654
rect 252836 145590 252888 145596
rect 252742 114472 252798 114481
rect 252742 114407 252798 114416
rect 253018 114472 253074 114481
rect 253018 114407 253074 114416
rect 253032 113257 253060 114407
rect 253018 113248 253074 113257
rect 253018 113183 253074 113192
rect 253020 112532 253072 112538
rect 253020 112474 253072 112480
rect 253032 111790 253060 112474
rect 252652 111784 252704 111790
rect 252652 111726 252704 111732
rect 253020 111784 253072 111790
rect 253020 111726 253072 111732
rect 252560 109744 252612 109750
rect 252560 109686 252612 109692
rect 251272 17332 251324 17338
rect 251272 17274 251324 17280
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 251284 3482 251312 17274
rect 252664 16574 252692 111726
rect 255240 74594 255268 197950
rect 255964 192500 256016 192506
rect 255964 192442 256016 192448
rect 255320 146804 255372 146810
rect 255320 146746 255372 146752
rect 255332 146334 255360 146746
rect 255320 146328 255372 146334
rect 255320 146270 255372 146276
rect 255228 74588 255280 74594
rect 255228 74530 255280 74536
rect 255332 16574 255360 146270
rect 255976 123486 256004 192442
rect 256068 146810 256096 215970
rect 256146 203552 256202 203561
rect 256146 203487 256202 203496
rect 256160 169017 256188 203487
rect 256620 192506 256648 219263
rect 256712 206310 256740 291774
rect 256804 243273 256832 292182
rect 256896 278089 256924 311918
rect 256974 305824 257030 305833
rect 256974 305759 257030 305768
rect 256988 288425 257016 305759
rect 258080 305720 258132 305726
rect 258080 305662 258132 305668
rect 256974 288416 257030 288425
rect 256974 288351 257030 288360
rect 257986 288416 258042 288425
rect 257986 288351 258042 288360
rect 258000 287745 258028 288351
rect 257986 287736 258042 287745
rect 257986 287671 258042 287680
rect 256882 278080 256938 278089
rect 256882 278015 256938 278024
rect 258092 275670 258120 305662
rect 258172 304292 258224 304298
rect 258172 304234 258224 304240
rect 258184 283898 258212 304234
rect 258736 302297 258764 324294
rect 259274 302424 259330 302433
rect 259274 302359 259330 302368
rect 258722 302288 258778 302297
rect 258722 302223 258778 302232
rect 259288 300218 259316 302359
rect 259276 300212 259328 300218
rect 259276 300154 259328 300160
rect 259276 300076 259328 300082
rect 259276 300018 259328 300024
rect 259288 298081 259316 300018
rect 259274 298072 259330 298081
rect 259274 298007 259330 298016
rect 259380 293282 259408 347686
rect 259736 320204 259788 320210
rect 259736 320146 259788 320152
rect 259552 311160 259604 311166
rect 259552 311102 259604 311108
rect 259460 307828 259512 307834
rect 259460 307770 259512 307776
rect 259472 304298 259500 307770
rect 259460 304292 259512 304298
rect 259460 304234 259512 304240
rect 259458 302288 259514 302297
rect 259458 302223 259514 302232
rect 259472 295662 259500 302223
rect 259460 295656 259512 295662
rect 259460 295598 259512 295604
rect 259368 293276 259420 293282
rect 259368 293218 259420 293224
rect 259460 289128 259512 289134
rect 259460 289070 259512 289076
rect 258172 283892 258224 283898
rect 258172 283834 258224 283840
rect 259276 283620 259328 283626
rect 259276 283562 259328 283568
rect 258722 282296 258778 282305
rect 258722 282231 258778 282240
rect 258356 278656 258408 278662
rect 258356 278598 258408 278604
rect 258368 278050 258396 278598
rect 258356 278044 258408 278050
rect 258356 277986 258408 277992
rect 258080 275664 258132 275670
rect 258080 275606 258132 275612
rect 256882 266928 256938 266937
rect 256882 266863 256938 266872
rect 256790 243264 256846 243273
rect 256790 243199 256846 243208
rect 256790 242312 256846 242321
rect 256790 242247 256846 242256
rect 256804 236609 256832 242247
rect 256896 239426 256924 266863
rect 258078 258224 258134 258233
rect 258078 258159 258134 258168
rect 256976 257372 257028 257378
rect 256976 257314 257028 257320
rect 256884 239420 256936 239426
rect 256884 239362 256936 239368
rect 256790 236600 256846 236609
rect 256790 236535 256846 236544
rect 256988 234598 257016 257314
rect 258092 255785 258120 258159
rect 258078 255776 258134 255785
rect 258078 255711 258134 255720
rect 258264 252748 258316 252754
rect 258264 252690 258316 252696
rect 257988 251320 258040 251326
rect 257988 251262 258040 251268
rect 258000 249422 258028 251262
rect 257988 249416 258040 249422
rect 257988 249358 258040 249364
rect 258170 246256 258226 246265
rect 258170 246191 258226 246200
rect 256976 234592 257028 234598
rect 256976 234534 257028 234540
rect 257344 231124 257396 231130
rect 257344 231066 257396 231072
rect 257356 214606 257384 231066
rect 258184 228449 258212 246191
rect 258276 240825 258304 252690
rect 258262 240816 258318 240825
rect 258262 240751 258318 240760
rect 258170 228440 258226 228449
rect 258170 228375 258226 228384
rect 257344 214600 257396 214606
rect 257344 214542 257396 214548
rect 256700 206304 256752 206310
rect 256700 206246 256752 206252
rect 256608 192500 256660 192506
rect 256608 192442 256660 192448
rect 256146 169008 256202 169017
rect 256146 168943 256202 168952
rect 256056 146804 256108 146810
rect 256056 146746 256108 146752
rect 255964 123480 256016 123486
rect 255964 123422 256016 123428
rect 256712 95849 256740 206246
rect 258368 205698 258396 277986
rect 258080 205692 258132 205698
rect 258080 205634 258132 205640
rect 258356 205692 258408 205698
rect 258356 205634 258408 205640
rect 256698 95840 256754 95849
rect 256698 95775 256754 95784
rect 258092 91050 258120 205634
rect 258736 135250 258764 282231
rect 259288 279478 259316 283562
rect 259366 283520 259422 283529
rect 259366 283455 259422 283464
rect 259380 282849 259408 283455
rect 259366 282840 259422 282849
rect 259366 282775 259422 282784
rect 259472 282305 259500 289070
rect 259564 287774 259592 311102
rect 259642 301472 259698 301481
rect 259642 301407 259698 301416
rect 259552 287768 259604 287774
rect 259552 287710 259604 287716
rect 259458 282296 259514 282305
rect 259458 282231 259514 282240
rect 259656 281081 259684 301407
rect 259748 285734 259776 320146
rect 260116 305658 260144 452610
rect 260196 438796 260248 438802
rect 260196 438738 260248 438744
rect 260208 319433 260236 438738
rect 260380 355360 260432 355366
rect 260380 355302 260432 355308
rect 260286 347032 260342 347041
rect 260286 346967 260342 346976
rect 260194 319424 260250 319433
rect 260194 319359 260250 319368
rect 260300 311409 260328 346967
rect 260392 328438 260420 355302
rect 260852 334694 260880 553454
rect 260944 341465 260972 560254
rect 261036 519586 261064 589290
rect 261024 519580 261076 519586
rect 261024 519522 261076 519528
rect 261116 454096 261168 454102
rect 261116 454038 261168 454044
rect 261024 451308 261076 451314
rect 261024 451250 261076 451256
rect 260930 341456 260986 341465
rect 260930 341391 260986 341400
rect 260840 334688 260892 334694
rect 260840 334630 260892 334636
rect 260380 328432 260432 328438
rect 260380 328374 260432 328380
rect 260840 323808 260892 323814
rect 260840 323750 260892 323756
rect 260852 323066 260880 323750
rect 260840 323060 260892 323066
rect 260840 323002 260892 323008
rect 260286 311400 260342 311409
rect 260286 311335 260342 311344
rect 260104 305652 260156 305658
rect 260104 305594 260156 305600
rect 259826 296712 259882 296721
rect 259826 296647 259882 296656
rect 259840 296614 259868 296647
rect 259828 296608 259880 296614
rect 259828 296550 259880 296556
rect 260748 296608 260800 296614
rect 260748 296550 260800 296556
rect 260760 295390 260788 296550
rect 260748 295384 260800 295390
rect 260748 295326 260800 295332
rect 260852 291106 260880 323002
rect 261036 316034 261064 451250
rect 261128 347750 261156 454038
rect 262232 389065 262260 598975
rect 263600 547936 263652 547942
rect 263600 547878 263652 547884
rect 262312 541000 262364 541006
rect 262312 540942 262364 540948
rect 262324 454034 262352 540942
rect 262404 458924 262456 458930
rect 262404 458866 262456 458872
rect 262312 454028 262364 454034
rect 262312 453970 262364 453976
rect 262310 452840 262366 452849
rect 262310 452775 262366 452784
rect 262218 389056 262274 389065
rect 262218 388991 262274 389000
rect 262220 378072 262272 378078
rect 262220 378014 262272 378020
rect 261116 347744 261168 347750
rect 261116 347686 261168 347692
rect 261208 347132 261260 347138
rect 261208 347074 261260 347080
rect 261220 323814 261248 347074
rect 261208 323808 261260 323814
rect 261208 323750 261260 323756
rect 260944 316006 261064 316034
rect 260944 313342 260972 316006
rect 260932 313336 260984 313342
rect 260932 313278 260984 313284
rect 260840 291100 260892 291106
rect 260840 291042 260892 291048
rect 259736 285728 259788 285734
rect 259736 285670 259788 285676
rect 260102 282160 260158 282169
rect 260102 282095 260158 282104
rect 259642 281072 259698 281081
rect 259642 281007 259698 281016
rect 259458 279848 259514 279857
rect 259458 279783 259514 279792
rect 259276 279472 259328 279478
rect 259276 279414 259328 279420
rect 259368 270836 259420 270842
rect 259368 270778 259420 270784
rect 259380 269822 259408 270778
rect 259368 269816 259420 269822
rect 259368 269758 259420 269764
rect 259368 266416 259420 266422
rect 259368 266358 259420 266364
rect 259380 264178 259408 266358
rect 259368 264172 259420 264178
rect 259368 264114 259420 264120
rect 259368 261384 259420 261390
rect 259368 261326 259420 261332
rect 259380 260166 259408 261326
rect 259368 260160 259420 260166
rect 259368 260102 259420 260108
rect 259472 241466 259500 279783
rect 259642 266520 259698 266529
rect 259642 266455 259698 266464
rect 259552 257372 259604 257378
rect 259552 257314 259604 257320
rect 259564 251326 259592 257314
rect 259552 251320 259604 251326
rect 259552 251262 259604 251268
rect 259552 249416 259604 249422
rect 259552 249358 259604 249364
rect 259460 241460 259512 241466
rect 259460 241402 259512 241408
rect 258816 239420 258868 239426
rect 258816 239362 258868 239368
rect 258828 219434 258856 239362
rect 258816 219428 258868 219434
rect 258816 219370 258868 219376
rect 258724 135244 258776 135250
rect 258724 135186 258776 135192
rect 259472 129742 259500 241402
rect 259564 160750 259592 249358
rect 259656 233238 259684 266455
rect 260116 266218 260144 282095
rect 260944 273970 260972 313278
rect 261022 300656 261078 300665
rect 261022 300591 261078 300600
rect 260932 273964 260984 273970
rect 260932 273906 260984 273912
rect 260104 266212 260156 266218
rect 260104 266154 260156 266160
rect 259736 263764 259788 263770
rect 259736 263706 259788 263712
rect 259748 233918 259776 263706
rect 260748 263628 260800 263634
rect 260748 263570 260800 263576
rect 260760 263537 260788 263570
rect 260746 263528 260802 263537
rect 260746 263463 260802 263472
rect 260746 260536 260802 260545
rect 260746 260471 260748 260480
rect 260800 260471 260802 260480
rect 260748 260442 260800 260448
rect 259736 233912 259788 233918
rect 259736 233854 259788 233860
rect 259644 233232 259696 233238
rect 259644 233174 259696 233180
rect 260196 200864 260248 200870
rect 260196 200806 260248 200812
rect 259552 160744 259604 160750
rect 259552 160686 259604 160692
rect 259460 129736 259512 129742
rect 259460 129678 259512 129684
rect 260104 127696 260156 127702
rect 260104 127638 260156 127644
rect 258722 113248 258778 113257
rect 258722 113183 258778 113192
rect 258080 91044 258132 91050
rect 258080 90986 258132 90992
rect 252664 16546 253520 16574
rect 255332 16546 255912 16574
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253492 480 253520 16546
rect 254676 7608 254728 7614
rect 254676 7550 254728 7556
rect 254688 480 254716 7550
rect 255884 480 255912 16546
rect 256700 15904 256752 15910
rect 256700 15846 256752 15852
rect 256712 490 256740 15846
rect 258264 8968 258316 8974
rect 258264 8910 258316 8916
rect 256896 598 257108 626
rect 256896 490 256924 598
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 462 256924 490
rect 257080 480 257108 598
rect 258276 480 258304 8910
rect 258736 8294 258764 113183
rect 259460 51740 259512 51746
rect 259460 51682 259512 51688
rect 258724 8288 258776 8294
rect 258724 8230 258776 8236
rect 259472 480 259500 51682
rect 260116 17270 260144 127638
rect 260208 111790 260236 200806
rect 260944 191146 260972 273906
rect 261036 242214 261064 300591
rect 262128 300144 262180 300150
rect 262128 300086 262180 300092
rect 262140 299470 262168 300086
rect 262128 299464 262180 299470
rect 262128 299406 262180 299412
rect 261206 291272 261262 291281
rect 261206 291207 261262 291216
rect 261114 254008 261170 254017
rect 261114 253943 261170 253952
rect 261024 242208 261076 242214
rect 261024 242150 261076 242156
rect 261128 239465 261156 253943
rect 261114 239456 261170 239465
rect 261114 239391 261170 239400
rect 260932 191140 260984 191146
rect 260932 191082 260984 191088
rect 261220 159390 261248 291207
rect 261484 290488 261536 290494
rect 261484 290430 261536 290436
rect 261496 273222 261524 290430
rect 262232 285297 262260 378014
rect 262324 347857 262352 452775
rect 262416 407862 262444 458866
rect 262864 434036 262916 434042
rect 262864 433978 262916 433984
rect 262876 432614 262904 433978
rect 262864 432608 262916 432614
rect 262864 432550 262916 432556
rect 262496 431248 262548 431254
rect 262496 431190 262548 431196
rect 262404 407856 262456 407862
rect 262404 407798 262456 407804
rect 262508 398206 262536 431190
rect 262864 403640 262916 403646
rect 262864 403582 262916 403588
rect 262496 398200 262548 398206
rect 262496 398142 262548 398148
rect 262876 378078 262904 403582
rect 262864 378072 262916 378078
rect 262864 378014 262916 378020
rect 263612 366382 263640 547878
rect 263704 480254 263732 601734
rect 265072 590708 265124 590714
rect 265072 590650 265124 590656
rect 264980 576904 265032 576910
rect 264980 576846 265032 576852
rect 263704 480226 263824 480254
rect 263796 461009 263824 480226
rect 263782 461000 263838 461009
rect 263782 460935 263838 460944
rect 263692 442332 263744 442338
rect 263692 442274 263744 442280
rect 263704 383042 263732 442274
rect 263796 438870 263824 460935
rect 263784 438864 263836 438870
rect 263784 438806 263836 438812
rect 263796 437510 263824 438806
rect 263784 437504 263836 437510
rect 263784 437446 263836 437452
rect 264244 435396 264296 435402
rect 264244 435338 264296 435344
rect 263784 431996 263836 432002
rect 263784 431938 263836 431944
rect 263692 383036 263744 383042
rect 263692 382978 263744 382984
rect 263796 373318 263824 431938
rect 264256 389230 264284 435338
rect 264244 389224 264296 389230
rect 264244 389166 264296 389172
rect 263968 375420 264020 375426
rect 263968 375362 264020 375368
rect 263784 373312 263836 373318
rect 263784 373254 263836 373260
rect 263600 366376 263652 366382
rect 263600 366318 263652 366324
rect 263600 362296 263652 362302
rect 263600 362238 263652 362244
rect 262404 354000 262456 354006
rect 262404 353942 262456 353948
rect 262310 347848 262366 347857
rect 262310 347783 262366 347792
rect 262218 285288 262274 285297
rect 262218 285223 262274 285232
rect 262220 284980 262272 284986
rect 262220 284922 262272 284928
rect 262232 283937 262260 284922
rect 262218 283928 262274 283937
rect 262218 283863 262274 283872
rect 262324 277137 262352 347783
rect 262416 278662 262444 353942
rect 262864 315308 262916 315314
rect 262864 315250 262916 315256
rect 262876 306202 262904 315250
rect 262864 306196 262916 306202
rect 262864 306138 262916 306144
rect 262496 303680 262548 303686
rect 262494 303648 262496 303657
rect 262548 303648 262550 303657
rect 262494 303583 262550 303592
rect 262862 299568 262918 299577
rect 262862 299503 262918 299512
rect 262876 291854 262904 299503
rect 263612 291922 263640 362238
rect 263876 311908 263928 311914
rect 263876 311850 263928 311856
rect 263784 296812 263836 296818
rect 263784 296754 263836 296760
rect 263600 291916 263652 291922
rect 263600 291858 263652 291864
rect 262864 291848 262916 291854
rect 262864 291790 262916 291796
rect 263600 285728 263652 285734
rect 263600 285670 263652 285676
rect 263138 285288 263194 285297
rect 263138 285223 263194 285232
rect 263152 284345 263180 285223
rect 263138 284336 263194 284345
rect 263138 284271 263194 284280
rect 262586 281072 262642 281081
rect 262586 281007 262642 281016
rect 262404 278656 262456 278662
rect 262404 278598 262456 278604
rect 262310 277128 262366 277137
rect 262310 277063 262366 277072
rect 261484 273216 261536 273222
rect 261484 273158 261536 273164
rect 262404 271856 262456 271862
rect 262404 271798 262456 271804
rect 262416 270609 262444 271798
rect 262402 270600 262458 270609
rect 262402 270535 262458 270544
rect 262218 270464 262274 270473
rect 262218 270399 262274 270408
rect 262232 270201 262260 270399
rect 262218 270192 262274 270201
rect 262218 270127 262274 270136
rect 261482 262304 261538 262313
rect 261482 262239 261538 262248
rect 261496 258058 261524 262239
rect 261484 258052 261536 258058
rect 261484 257994 261536 258000
rect 262232 215966 262260 270127
rect 262416 227730 262444 270535
rect 262496 251184 262548 251190
rect 262496 251126 262548 251132
rect 262508 250578 262536 251126
rect 262496 250572 262548 250578
rect 262496 250514 262548 250520
rect 262508 228313 262536 250514
rect 262494 228304 262550 228313
rect 262494 228239 262550 228248
rect 262404 227724 262456 227730
rect 262404 227666 262456 227672
rect 262220 215960 262272 215966
rect 262220 215902 262272 215908
rect 261484 195356 261536 195362
rect 261484 195298 261536 195304
rect 261208 159384 261260 159390
rect 261208 159326 261260 159332
rect 260196 111784 260248 111790
rect 260196 111726 260248 111732
rect 261496 84182 261524 195298
rect 262232 88330 262260 215902
rect 262416 116618 262444 227666
rect 262600 164898 262628 281007
rect 262864 278044 262916 278050
rect 262864 277986 262916 277992
rect 262876 251190 262904 277986
rect 262864 251184 262916 251190
rect 262864 251126 262916 251132
rect 263612 166326 263640 285670
rect 263690 284336 263746 284345
rect 263690 284271 263746 284280
rect 263704 207058 263732 284271
rect 263796 240786 263824 296754
rect 263888 285666 263916 311850
rect 263876 285660 263928 285666
rect 263876 285602 263928 285608
rect 263980 280158 264008 375362
rect 264992 318073 265020 576846
rect 265084 359417 265112 590650
rect 266372 561066 266400 697546
rect 267740 596216 267792 596222
rect 267740 596158 267792 596164
rect 266360 561060 266412 561066
rect 266360 561002 266412 561008
rect 266360 557592 266412 557598
rect 266360 557534 266412 557540
rect 265164 525088 265216 525094
rect 265164 525030 265216 525036
rect 265176 387705 265204 525030
rect 265254 480856 265310 480865
rect 265254 480791 265310 480800
rect 265162 387696 265218 387705
rect 265162 387631 265218 387640
rect 265164 374060 265216 374066
rect 265164 374002 265216 374008
rect 265070 359408 265126 359417
rect 265070 359343 265126 359352
rect 264978 318064 265034 318073
rect 264978 317999 265034 318008
rect 264980 316736 265032 316742
rect 264980 316678 265032 316684
rect 264992 282810 265020 316678
rect 265072 306196 265124 306202
rect 265072 306138 265124 306144
rect 265084 290494 265112 306138
rect 265072 290488 265124 290494
rect 265072 290430 265124 290436
rect 264980 282804 265032 282810
rect 264980 282746 265032 282752
rect 263968 280152 264020 280158
rect 263968 280094 264020 280100
rect 264980 280152 265032 280158
rect 264980 280094 265032 280100
rect 263980 279721 264008 280094
rect 263966 279712 264022 279721
rect 263966 279647 264022 279656
rect 263874 262712 263930 262721
rect 263874 262647 263930 262656
rect 263888 262342 263916 262647
rect 263876 262336 263928 262342
rect 263876 262278 263928 262284
rect 263784 240780 263836 240786
rect 263784 240722 263836 240728
rect 263888 216617 263916 262278
rect 263874 216608 263930 216617
rect 263874 216543 263930 216552
rect 264992 212498 265020 280094
rect 265176 259418 265204 374002
rect 265268 370530 265296 480791
rect 265714 387696 265770 387705
rect 265714 387631 265770 387640
rect 265728 387122 265756 387631
rect 265716 387116 265768 387122
rect 265716 387058 265768 387064
rect 265256 370524 265308 370530
rect 265256 370466 265308 370472
rect 266372 327758 266400 557534
rect 266452 543788 266504 543794
rect 266452 543730 266504 543736
rect 266464 336025 266492 543730
rect 266544 527944 266596 527950
rect 266544 527886 266596 527892
rect 266556 386209 266584 527886
rect 266636 437504 266688 437510
rect 266636 437446 266688 437452
rect 266542 386200 266598 386209
rect 266542 386135 266598 386144
rect 266450 336016 266506 336025
rect 266450 335951 266506 335960
rect 266360 327752 266412 327758
rect 266360 327694 266412 327700
rect 266648 318850 266676 437446
rect 267002 386200 267058 386209
rect 267002 386135 267058 386144
rect 267016 385694 267044 386135
rect 267004 385688 267056 385694
rect 267004 385630 267056 385636
rect 267752 369209 267780 596158
rect 269120 564460 269172 564466
rect 269120 564402 269172 564408
rect 267924 480344 267976 480350
rect 267924 480286 267976 480292
rect 267936 436082 267964 480286
rect 268016 449200 268068 449206
rect 268016 449142 268068 449148
rect 267924 436076 267976 436082
rect 267924 436018 267976 436024
rect 267924 432608 267976 432614
rect 267924 432550 267976 432556
rect 267832 407788 267884 407794
rect 267832 407730 267884 407736
rect 267738 369200 267794 369209
rect 267738 369135 267794 369144
rect 267844 368393 267872 407730
rect 267830 368384 267886 368393
rect 267830 368319 267886 368328
rect 267738 334112 267794 334121
rect 267738 334047 267794 334056
rect 266728 328432 266780 328438
rect 266728 328374 266780 328380
rect 266636 318844 266688 318850
rect 266636 318786 266688 318792
rect 266544 317484 266596 317490
rect 266544 317426 266596 317432
rect 265622 298072 265678 298081
rect 265622 298007 265678 298016
rect 265636 297430 265664 298007
rect 265624 297424 265676 297430
rect 265624 297366 265676 297372
rect 265254 260264 265310 260273
rect 265254 260199 265310 260208
rect 265164 259412 265216 259418
rect 265164 259354 265216 259360
rect 265162 259176 265218 259185
rect 265268 259162 265296 260199
rect 265218 259134 265296 259162
rect 265162 259111 265218 259120
rect 265072 255400 265124 255406
rect 265072 255342 265124 255348
rect 265084 252113 265112 255342
rect 265070 252104 265126 252113
rect 265070 252039 265126 252048
rect 265070 247752 265126 247761
rect 265070 247687 265072 247696
rect 265124 247687 265126 247696
rect 265072 247658 265124 247664
rect 265176 238754 265204 259111
rect 265084 238726 265204 238754
rect 265084 225622 265112 238726
rect 265072 225616 265124 225622
rect 265072 225558 265124 225564
rect 264980 212492 265032 212498
rect 264980 212434 265032 212440
rect 263692 207052 263744 207058
rect 263692 206994 263744 207000
rect 263600 166320 263652 166326
rect 263600 166262 263652 166268
rect 262588 164892 262640 164898
rect 262588 164834 262640 164840
rect 263600 155236 263652 155242
rect 263600 155178 263652 155184
rect 263612 154630 263640 155178
rect 263600 154624 263652 154630
rect 263600 154566 263652 154572
rect 262404 116612 262456 116618
rect 262404 116554 262456 116560
rect 262220 88324 262272 88330
rect 262220 88266 262272 88272
rect 261484 84176 261536 84182
rect 261484 84118 261536 84124
rect 262218 79520 262274 79529
rect 262218 79455 262274 79464
rect 260104 17264 260156 17270
rect 260104 17206 260156 17212
rect 262232 16574 262260 79455
rect 262232 16546 262536 16574
rect 261760 8288 261812 8294
rect 261760 8230 261812 8236
rect 260656 3188 260708 3194
rect 260656 3130 260708 3136
rect 260668 480 260696 3130
rect 261772 480 261800 8230
rect 262508 490 262536 16546
rect 263612 3194 263640 154566
rect 263704 94518 263732 206994
rect 264992 98666 265020 212434
rect 265072 206984 265124 206990
rect 265070 206952 265072 206961
rect 265124 206952 265126 206961
rect 265070 206887 265126 206896
rect 265636 153882 265664 297366
rect 266450 295080 266506 295089
rect 266450 295015 266506 295024
rect 266358 284336 266414 284345
rect 266358 284271 266414 284280
rect 265716 247104 265768 247110
rect 265716 247046 265768 247052
rect 265728 206990 265756 247046
rect 266372 220114 266400 284271
rect 266464 236706 266492 295015
rect 266556 284306 266584 317426
rect 266648 285841 266676 318786
rect 266634 285832 266690 285841
rect 266634 285767 266690 285776
rect 266740 284345 266768 328374
rect 267752 322153 267780 334047
rect 267738 322144 267794 322153
rect 267738 322079 267794 322088
rect 267738 307048 267794 307057
rect 267738 306983 267794 306992
rect 267752 289814 267780 306983
rect 267740 289808 267792 289814
rect 267740 289750 267792 289756
rect 267738 287736 267794 287745
rect 267738 287671 267794 287680
rect 266726 284336 266782 284345
rect 266544 284300 266596 284306
rect 266726 284271 266782 284280
rect 266544 284242 266596 284248
rect 266542 269376 266598 269385
rect 266542 269311 266598 269320
rect 266556 238649 266584 269311
rect 266634 252240 266690 252249
rect 266634 252175 266690 252184
rect 266542 238640 266598 238649
rect 266542 238575 266598 238584
rect 266452 236700 266504 236706
rect 266452 236642 266504 236648
rect 266648 233209 266676 252175
rect 267094 235240 267150 235249
rect 267094 235175 267150 235184
rect 266634 233200 266690 233209
rect 266634 233135 266690 233144
rect 267004 232620 267056 232626
rect 267004 232562 267056 232568
rect 266360 220108 266412 220114
rect 266360 220050 266412 220056
rect 265716 206984 265768 206990
rect 265716 206926 265768 206932
rect 265624 153876 265676 153882
rect 265624 153818 265676 153824
rect 266372 102134 266400 220050
rect 267016 141001 267044 232562
rect 267108 204241 267136 235175
rect 267094 204232 267150 204241
rect 267094 204167 267150 204176
rect 267752 158030 267780 287671
rect 267844 271862 267872 368319
rect 267936 345014 267964 432550
rect 268028 392601 268056 449142
rect 269028 433288 269080 433294
rect 269028 433230 269080 433236
rect 269040 432614 269068 433230
rect 269028 432608 269080 432614
rect 269028 432550 269080 432556
rect 268014 392592 268070 392601
rect 268014 392527 268070 392536
rect 267936 344986 268056 345014
rect 268028 341562 268056 344986
rect 268016 341556 268068 341562
rect 268016 341498 268068 341504
rect 268028 341465 268056 341498
rect 268014 341456 268070 341465
rect 268014 341391 268070 341400
rect 267922 323640 267978 323649
rect 267922 323575 267978 323584
rect 267832 271856 267884 271862
rect 267832 271798 267884 271804
rect 267936 267714 267964 323575
rect 269132 314129 269160 564402
rect 269212 552696 269264 552702
rect 269212 552638 269264 552644
rect 269224 472666 269252 552638
rect 269316 550594 269344 702782
rect 271144 702568 271196 702574
rect 271144 702510 271196 702516
rect 270500 587172 270552 587178
rect 270500 587114 270552 587120
rect 269304 550588 269356 550594
rect 269304 550530 269356 550536
rect 269764 476808 269816 476814
rect 269764 476750 269816 476756
rect 269212 472660 269264 472666
rect 269212 472602 269264 472608
rect 269394 466032 269450 466041
rect 269394 465967 269450 465976
rect 269212 446412 269264 446418
rect 269212 446354 269264 446360
rect 269118 314120 269174 314129
rect 269118 314055 269174 314064
rect 268016 302320 268068 302326
rect 268016 302262 268068 302268
rect 267924 267708 267976 267714
rect 267924 267650 267976 267656
rect 267832 262268 267884 262274
rect 267832 262210 267884 262216
rect 267740 158024 267792 158030
rect 267740 157966 267792 157972
rect 267002 140992 267058 141001
rect 267002 140927 267058 140936
rect 266360 102128 266412 102134
rect 266360 102070 266412 102076
rect 264980 98660 265032 98666
rect 264980 98602 265032 98608
rect 263692 94512 263744 94518
rect 263692 94454 263744 94460
rect 264980 58676 265032 58682
rect 264980 58618 265032 58624
rect 263692 29640 263744 29646
rect 263692 29582 263744 29588
rect 263704 16574 263732 29582
rect 263704 16546 264192 16574
rect 263600 3188 263652 3194
rect 263600 3130 263652 3136
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 264992 490 265020 58618
rect 266360 31068 266412 31074
rect 266360 31010 266412 31016
rect 266372 16574 266400 31010
rect 266372 16546 266584 16574
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 16546
rect 267016 4146 267044 140927
rect 267844 109818 267872 262210
rect 267924 250504 267976 250510
rect 267924 250446 267976 250452
rect 267936 250073 267964 250446
rect 267922 250064 267978 250073
rect 267922 249999 267978 250008
rect 268028 216034 268056 302262
rect 269118 285696 269174 285705
rect 269118 285631 269174 285640
rect 269028 268388 269080 268394
rect 269028 268330 269080 268336
rect 269040 267850 269068 268330
rect 268108 267844 268160 267850
rect 268108 267786 268160 267792
rect 269028 267844 269080 267850
rect 269028 267786 269080 267792
rect 268016 216028 268068 216034
rect 268016 215970 268068 215976
rect 268120 149802 268148 267786
rect 268290 262440 268346 262449
rect 268290 262375 268346 262384
rect 268304 262274 268332 262375
rect 268292 262268 268344 262274
rect 268292 262210 268344 262216
rect 269028 251184 269080 251190
rect 269028 251126 269080 251132
rect 269040 250510 269068 251126
rect 269028 250504 269080 250510
rect 269028 250446 269080 250452
rect 268108 149796 268160 149802
rect 268108 149738 268160 149744
rect 268382 142488 268438 142497
rect 268382 142423 268438 142432
rect 268396 127634 268424 142423
rect 269132 133890 269160 285631
rect 269224 247110 269252 446354
rect 269304 443692 269356 443698
rect 269304 443634 269356 443640
rect 269316 322998 269344 443634
rect 269408 389881 269436 465967
rect 269776 445058 269804 476750
rect 269764 445052 269816 445058
rect 269764 444994 269816 445000
rect 270512 403646 270540 587114
rect 270592 575544 270644 575550
rect 270592 575486 270644 575492
rect 270604 461650 270632 575486
rect 271156 536625 271184 702510
rect 271880 600432 271932 600438
rect 271880 600374 271932 600380
rect 271142 536616 271198 536625
rect 271142 536551 271198 536560
rect 270684 522300 270736 522306
rect 270684 522242 270736 522248
rect 270592 461644 270644 461650
rect 270592 461586 270644 461592
rect 270590 451344 270646 451353
rect 270590 451279 270646 451288
rect 270500 403640 270552 403646
rect 270500 403582 270552 403588
rect 269394 389872 269450 389881
rect 269394 389807 269450 389816
rect 270500 385688 270552 385694
rect 270500 385630 270552 385636
rect 269396 380180 269448 380186
rect 269396 380122 269448 380128
rect 269304 322992 269356 322998
rect 269304 322934 269356 322940
rect 269316 289134 269344 322934
rect 269304 289128 269356 289134
rect 269304 289070 269356 289076
rect 269408 272513 269436 380122
rect 269762 311264 269818 311273
rect 269762 311199 269818 311208
rect 269776 283665 269804 311199
rect 269762 283656 269818 283665
rect 269762 283591 269818 283600
rect 270512 274689 270540 385630
rect 270604 282169 270632 451279
rect 270696 380186 270724 522242
rect 271788 409148 271840 409154
rect 271788 409090 271840 409096
rect 271800 408542 271828 409090
rect 270776 408536 270828 408542
rect 270776 408478 270828 408484
rect 271788 408536 271840 408542
rect 271788 408478 271840 408484
rect 270684 380180 270736 380186
rect 270684 380122 270736 380128
rect 270788 362953 270816 408478
rect 270774 362944 270830 362953
rect 270774 362879 270830 362888
rect 270590 282160 270646 282169
rect 270590 282095 270646 282104
rect 270590 281480 270646 281489
rect 270590 281415 270646 281424
rect 270604 280673 270632 281415
rect 270590 280664 270646 280673
rect 270590 280599 270646 280608
rect 270498 274680 270554 274689
rect 270498 274615 270554 274624
rect 269394 272504 269450 272513
rect 269316 272462 269394 272490
rect 269212 247104 269264 247110
rect 269212 247046 269264 247052
rect 269316 223582 269344 272462
rect 269394 272439 269450 272448
rect 269396 267776 269448 267782
rect 269396 267718 269448 267724
rect 269408 235929 269436 267718
rect 270408 244316 270460 244322
rect 270408 244258 270460 244264
rect 270420 244225 270448 244258
rect 270406 244216 270462 244225
rect 270406 244151 270462 244160
rect 269764 241052 269816 241058
rect 269764 240994 269816 241000
rect 269394 235920 269450 235929
rect 269394 235855 269450 235864
rect 269304 223576 269356 223582
rect 269304 223518 269356 223524
rect 269120 133884 269172 133890
rect 269120 133826 269172 133832
rect 267924 127628 267976 127634
rect 267924 127570 267976 127576
rect 268384 127628 268436 127634
rect 268384 127570 268436 127576
rect 267832 109812 267884 109818
rect 267832 109754 267884 109760
rect 267936 16574 267964 127570
rect 269776 72486 269804 240994
rect 270512 211818 270540 274615
rect 270604 226273 270632 280599
rect 270682 273864 270738 273873
rect 270682 273799 270738 273808
rect 270590 226264 270646 226273
rect 270590 226199 270646 226208
rect 270590 222184 270646 222193
rect 270590 222119 270646 222128
rect 270604 221474 270632 222119
rect 270592 221468 270644 221474
rect 270592 221410 270644 221416
rect 270500 211812 270552 211818
rect 270500 211754 270552 211760
rect 270512 97481 270540 211754
rect 270604 108322 270632 221410
rect 270696 162858 270724 273799
rect 270788 271153 270816 362879
rect 271892 358057 271920 600374
rect 273352 597576 273404 597582
rect 273352 597518 273404 597524
rect 273260 558952 273312 558958
rect 273260 558894 273312 558900
rect 271972 546508 272024 546514
rect 271972 546450 272024 546456
rect 271984 389094 272012 546450
rect 272064 451376 272116 451382
rect 272064 451318 272116 451324
rect 271972 389088 272024 389094
rect 271972 389030 272024 389036
rect 271878 358048 271934 358057
rect 271878 357983 271934 357992
rect 272076 346497 272104 451318
rect 272156 394732 272208 394738
rect 272156 394674 272208 394680
rect 272168 364274 272196 394674
rect 273272 372570 273300 558894
rect 273364 465089 273392 597518
rect 274560 583710 274588 703054
rect 280804 702976 280856 702982
rect 280804 702918 280856 702924
rect 274824 604512 274876 604518
rect 274824 604454 274876 604460
rect 274548 583704 274600 583710
rect 274548 583646 274600 583652
rect 274560 583030 274588 583646
rect 274548 583024 274600 583030
rect 274548 582966 274600 582972
rect 273444 574116 273496 574122
rect 273444 574058 273496 574064
rect 273350 465080 273406 465089
rect 273350 465015 273406 465024
rect 273456 463690 273484 574058
rect 273536 533384 273588 533390
rect 273536 533326 273588 533332
rect 273444 463684 273496 463690
rect 273444 463626 273496 463632
rect 273548 425746 273576 533326
rect 273904 464364 273956 464370
rect 273904 464306 273956 464312
rect 273626 449984 273682 449993
rect 273626 449919 273682 449928
rect 273536 425740 273588 425746
rect 273536 425682 273588 425688
rect 273444 395344 273496 395350
rect 273444 395286 273496 395292
rect 273456 379273 273484 395286
rect 273442 379264 273498 379273
rect 273442 379199 273498 379208
rect 273456 379001 273484 379199
rect 273442 378992 273498 379001
rect 273442 378927 273498 378936
rect 273260 372564 273312 372570
rect 273260 372506 273312 372512
rect 272156 364268 272208 364274
rect 272156 364210 272208 364216
rect 272062 346488 272118 346497
rect 272062 346423 272118 346432
rect 271880 324964 271932 324970
rect 271880 324906 271932 324912
rect 271144 298172 271196 298178
rect 271144 298114 271196 298120
rect 271156 287706 271184 298114
rect 271144 287700 271196 287706
rect 271144 287642 271196 287648
rect 271892 282878 271920 324906
rect 271972 302252 272024 302258
rect 271972 302194 272024 302200
rect 271880 282872 271932 282878
rect 271880 282814 271932 282820
rect 271892 282470 271920 282814
rect 271880 282464 271932 282470
rect 271880 282406 271932 282412
rect 271880 276072 271932 276078
rect 271880 276014 271932 276020
rect 270774 271144 270830 271153
rect 270774 271079 270830 271088
rect 270774 248432 270830 248441
rect 270774 248367 270830 248376
rect 270788 239426 270816 248367
rect 270776 239420 270828 239426
rect 270776 239362 270828 239368
rect 270684 162852 270736 162858
rect 270684 162794 270736 162800
rect 271892 153202 271920 276014
rect 271984 200870 272012 302194
rect 272076 273193 272104 346423
rect 272168 295322 272196 364210
rect 272156 295316 272208 295322
rect 272156 295258 272208 295264
rect 272168 294642 272196 295258
rect 272156 294636 272208 294642
rect 272156 294578 272208 294584
rect 273272 281489 273300 372506
rect 273536 333328 273588 333334
rect 273536 333270 273588 333276
rect 273442 303920 273498 303929
rect 273442 303855 273498 303864
rect 273352 282464 273404 282470
rect 273352 282406 273404 282412
rect 273258 281480 273314 281489
rect 273258 281415 273314 281424
rect 272340 276684 272392 276690
rect 272340 276626 272392 276632
rect 272352 276078 272380 276626
rect 272340 276072 272392 276078
rect 272340 276014 272392 276020
rect 273258 276040 273314 276049
rect 273258 275975 273314 275984
rect 272062 273184 272118 273193
rect 272062 273119 272118 273128
rect 272076 272542 272104 273119
rect 272064 272536 272116 272542
rect 272064 272478 272116 272484
rect 272340 254652 272392 254658
rect 272340 254594 272392 254600
rect 272352 253978 272380 254594
rect 272064 253972 272116 253978
rect 272064 253914 272116 253920
rect 272340 253972 272392 253978
rect 272340 253914 272392 253920
rect 272076 224942 272104 253914
rect 272064 224936 272116 224942
rect 272064 224878 272116 224884
rect 271972 200864 272024 200870
rect 271972 200806 272024 200812
rect 271880 153196 271932 153202
rect 271880 153138 271932 153144
rect 273272 131102 273300 275975
rect 273364 212566 273392 282406
rect 273456 241058 273484 303855
rect 273548 283626 273576 333270
rect 273536 283620 273588 283626
rect 273536 283562 273588 283568
rect 273640 269385 273668 449919
rect 273916 391270 273944 464306
rect 274732 463820 274784 463826
rect 274732 463762 274784 463768
rect 273904 391264 273956 391270
rect 273904 391206 273956 391212
rect 274640 337408 274692 337414
rect 274640 337350 274692 337356
rect 273626 269376 273682 269385
rect 273626 269311 273682 269320
rect 273904 259412 273956 259418
rect 273904 259354 273956 259360
rect 273444 241052 273496 241058
rect 273444 240994 273496 241000
rect 273916 238746 273944 259354
rect 273904 238740 273956 238746
rect 273904 238682 273956 238688
rect 274652 238678 274680 337350
rect 274744 259418 274772 463762
rect 274836 435402 274864 604454
rect 278042 601896 278098 601905
rect 278042 601831 278098 601840
rect 276018 599176 276074 599185
rect 276018 599111 276074 599120
rect 274916 565956 274968 565962
rect 274916 565898 274968 565904
rect 274824 435396 274876 435402
rect 274824 435338 274876 435344
rect 274824 424380 274876 424386
rect 274824 424322 274876 424328
rect 274836 351898 274864 424322
rect 274824 351892 274876 351898
rect 274824 351834 274876 351840
rect 274836 279449 274864 351834
rect 274928 331809 274956 565898
rect 276032 468489 276060 599111
rect 277492 584452 277544 584458
rect 277492 584394 277544 584400
rect 277400 563100 277452 563106
rect 277400 563042 277452 563048
rect 276112 550588 276164 550594
rect 276112 550530 276164 550536
rect 276018 468480 276074 468489
rect 276018 468415 276074 468424
rect 276032 433362 276060 468415
rect 276124 455394 276152 550530
rect 276204 482316 276256 482322
rect 276204 482258 276256 482264
rect 276112 455388 276164 455394
rect 276112 455330 276164 455336
rect 276020 433356 276072 433362
rect 276020 433298 276072 433304
rect 276020 398132 276072 398138
rect 276020 398074 276072 398080
rect 276032 376689 276060 398074
rect 276216 396778 276244 482258
rect 276296 458720 276348 458726
rect 276296 458662 276348 458668
rect 277308 458720 277360 458726
rect 277308 458662 277360 458668
rect 276308 458425 276336 458662
rect 276294 458416 276350 458425
rect 276294 458351 276350 458360
rect 276388 455388 276440 455394
rect 276388 455330 276440 455336
rect 276400 454714 276428 455330
rect 276388 454708 276440 454714
rect 276388 454650 276440 454656
rect 276296 436076 276348 436082
rect 276296 436018 276348 436024
rect 276204 396772 276256 396778
rect 276204 396714 276256 396720
rect 276110 382936 276166 382945
rect 276110 382871 276166 382880
rect 276018 376680 276074 376689
rect 276018 376615 276074 376624
rect 274914 331800 274970 331809
rect 274914 331735 274970 331744
rect 274916 309188 274968 309194
rect 274916 309130 274968 309136
rect 274928 283529 274956 309130
rect 276018 309088 276074 309097
rect 276018 309023 276074 309032
rect 276032 307873 276060 309023
rect 276018 307864 276074 307873
rect 276018 307799 276074 307808
rect 274914 283520 274970 283529
rect 274914 283455 274970 283464
rect 274822 279440 274878 279449
rect 274822 279375 274878 279384
rect 276032 276049 276060 307799
rect 276018 276040 276074 276049
rect 276018 275975 276074 275984
rect 276124 271833 276152 382871
rect 276308 309097 276336 436018
rect 276480 398812 276532 398818
rect 276480 398754 276532 398760
rect 276492 398138 276520 398754
rect 276480 398132 276532 398138
rect 276480 398074 276532 398080
rect 277320 389842 277348 458662
rect 277308 389836 277360 389842
rect 277308 389778 277360 389784
rect 277412 342922 277440 563042
rect 277504 398818 277532 584394
rect 277584 553444 277636 553450
rect 277584 553386 277636 553392
rect 277596 499574 277624 553386
rect 278056 542366 278084 601831
rect 280160 599004 280212 599010
rect 280160 598946 280212 598952
rect 278780 580304 278832 580310
rect 278780 580246 278832 580252
rect 278044 542360 278096 542366
rect 278044 542302 278096 542308
rect 277596 499546 277716 499574
rect 277688 496126 277716 499546
rect 277860 497548 277912 497554
rect 277860 497490 277912 497496
rect 277676 496120 277728 496126
rect 277676 496062 277728 496068
rect 277688 457502 277716 496062
rect 277676 457496 277728 457502
rect 277676 457438 277728 457444
rect 277768 422340 277820 422346
rect 277768 422282 277820 422288
rect 277492 398812 277544 398818
rect 277492 398754 277544 398760
rect 277676 380928 277728 380934
rect 277676 380870 277728 380876
rect 277490 369064 277546 369073
rect 277490 368999 277546 369008
rect 277400 342916 277452 342922
rect 277400 342858 277452 342864
rect 277400 322244 277452 322250
rect 277400 322186 277452 322192
rect 276294 309088 276350 309097
rect 276294 309023 276350 309032
rect 276296 305652 276348 305658
rect 276296 305594 276348 305600
rect 276204 296744 276256 296750
rect 276204 296686 276256 296692
rect 276110 271824 276166 271833
rect 276110 271759 276166 271768
rect 274822 265568 274878 265577
rect 274822 265503 274878 265512
rect 274732 259412 274784 259418
rect 274732 259354 274784 259360
rect 274730 257952 274786 257961
rect 274730 257887 274786 257896
rect 274640 238672 274692 238678
rect 274640 238614 274692 238620
rect 273352 212560 273404 212566
rect 273352 212502 273404 212508
rect 273260 131096 273312 131102
rect 273260 131038 273312 131044
rect 270592 108316 270644 108322
rect 270592 108258 270644 108264
rect 270498 97472 270554 97481
rect 270498 97407 270554 97416
rect 273364 89690 273392 212502
rect 274640 204740 274692 204746
rect 274640 204682 274692 204688
rect 274652 204338 274680 204682
rect 274640 204332 274692 204338
rect 274640 204274 274692 204280
rect 274652 120766 274680 204274
rect 274744 177342 274772 257887
rect 274836 204746 274864 265503
rect 276020 264240 276072 264246
rect 276020 264182 276072 264188
rect 276032 261526 276060 264182
rect 276020 261520 276072 261526
rect 276020 261462 276072 261468
rect 274916 255332 274968 255338
rect 274916 255274 274968 255280
rect 274928 232558 274956 255274
rect 274916 232552 274968 232558
rect 274916 232494 274968 232500
rect 274824 204740 274876 204746
rect 274824 204682 274876 204688
rect 274732 177336 274784 177342
rect 274732 177278 274784 177284
rect 276032 149054 276060 261462
rect 276216 195362 276244 296686
rect 276308 232626 276336 305594
rect 277412 288386 277440 322186
rect 277400 288380 277452 288386
rect 277400 288322 277452 288328
rect 277504 243574 277532 368999
rect 277584 304292 277636 304298
rect 277584 304234 277636 304240
rect 277492 243568 277544 243574
rect 277492 243510 277544 243516
rect 277504 238754 277532 243510
rect 277412 238726 277532 238754
rect 276296 232620 276348 232626
rect 276296 232562 276348 232568
rect 276204 195356 276256 195362
rect 276204 195298 276256 195304
rect 276664 160132 276716 160138
rect 276664 160074 276716 160080
rect 276020 149048 276072 149054
rect 276020 148990 276072 148996
rect 276020 131776 276072 131782
rect 276020 131718 276072 131724
rect 274640 120760 274692 120766
rect 274640 120702 274692 120708
rect 273352 89684 273404 89690
rect 273352 89626 273404 89632
rect 270592 84856 270644 84862
rect 270592 84798 270644 84804
rect 269028 72480 269080 72486
rect 269028 72422 269080 72428
rect 269764 72480 269816 72486
rect 269764 72422 269816 72428
rect 267936 16546 268424 16574
rect 267004 4140 267056 4146
rect 267004 4082 267056 4088
rect 267740 4140 267792 4146
rect 267740 4082 267792 4088
rect 267752 480 267780 4082
rect 268396 490 268424 16546
rect 269040 3505 269068 72422
rect 269764 61396 269816 61402
rect 269764 61338 269816 61344
rect 269026 3496 269082 3505
rect 269026 3431 269082 3440
rect 269776 3194 269804 61338
rect 270500 53100 270552 53106
rect 270500 53042 270552 53048
rect 270040 3528 270092 3534
rect 270040 3470 270092 3476
rect 269764 3188 269816 3194
rect 269764 3130 269816 3136
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 3470
rect 270512 626 270540 53042
rect 270604 3534 270632 84798
rect 273258 80744 273314 80753
rect 273258 80679 273314 80688
rect 270592 3528 270644 3534
rect 270592 3470 270644 3476
rect 272432 3188 272484 3194
rect 272432 3130 272484 3136
rect 270512 598 270816 626
rect 270788 490 270816 598
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3130
rect 273272 490 273300 80679
rect 276032 6914 276060 131718
rect 276676 16574 276704 160074
rect 277412 86873 277440 238726
rect 277596 192574 277624 304234
rect 277688 276010 277716 380870
rect 277780 322250 277808 422282
rect 277872 386345 277900 497490
rect 277858 386336 277914 386345
rect 277858 386271 277914 386280
rect 277768 322244 277820 322250
rect 277768 322186 277820 322192
rect 278792 309233 278820 580246
rect 278872 571396 278924 571402
rect 278872 571338 278924 571344
rect 278884 458726 278912 571338
rect 278962 469296 279018 469305
rect 278962 469231 279018 469240
rect 278872 458720 278924 458726
rect 278872 458662 278924 458668
rect 278872 445052 278924 445058
rect 278872 444994 278924 445000
rect 278884 393990 278912 444994
rect 278976 416770 279004 469231
rect 279424 451920 279476 451926
rect 279424 451862 279476 451868
rect 278964 416764 279016 416770
rect 278964 416706 279016 416712
rect 279332 416764 279384 416770
rect 279332 416706 279384 416712
rect 279344 416673 279372 416706
rect 279330 416664 279386 416673
rect 279330 416599 279386 416608
rect 278872 393984 278924 393990
rect 278872 393926 278924 393932
rect 278872 393372 278924 393378
rect 278872 393314 278924 393320
rect 278884 349858 278912 393314
rect 278872 349852 278924 349858
rect 278872 349794 278924 349800
rect 278778 309224 278834 309233
rect 278778 309159 278834 309168
rect 278778 298752 278834 298761
rect 278778 298687 278834 298696
rect 277676 276004 277728 276010
rect 277676 275946 277728 275952
rect 277674 271824 277730 271833
rect 277674 271759 277730 271768
rect 277688 209681 277716 271759
rect 278044 248464 278096 248470
rect 278044 248406 278096 248412
rect 278056 233238 278084 248406
rect 278044 233232 278096 233238
rect 278044 233174 278096 233180
rect 277674 209672 277730 209681
rect 277674 209607 277730 209616
rect 277584 192568 277636 192574
rect 277584 192510 277636 192516
rect 278044 104848 278096 104854
rect 278044 104790 278096 104796
rect 277398 86864 277454 86873
rect 277398 86799 277454 86808
rect 277400 28280 277452 28286
rect 277400 28222 277452 28228
rect 277412 16574 277440 28222
rect 276676 16546 276796 16574
rect 277412 16546 277992 16574
rect 276032 6886 276704 6914
rect 276020 4412 276072 4418
rect 276020 4354 276072 4360
rect 274822 3496 274878 3505
rect 274822 3431 274878 3440
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 3431
rect 276032 480 276060 4354
rect 276676 490 276704 6886
rect 276768 3466 276796 16546
rect 277964 3482 277992 16546
rect 278056 4418 278084 104790
rect 278686 86864 278742 86873
rect 278686 86799 278742 86808
rect 278700 85649 278728 86799
rect 278686 85640 278742 85649
rect 278686 85575 278742 85584
rect 278792 77217 278820 298687
rect 278884 277370 278912 349794
rect 278962 309224 279018 309233
rect 278962 309159 279018 309168
rect 278872 277364 278924 277370
rect 278872 277306 278924 277312
rect 278976 262177 279004 309159
rect 278962 262168 279018 262177
rect 278962 262103 279018 262112
rect 278964 260160 279016 260166
rect 278964 260102 279016 260108
rect 278872 251864 278924 251870
rect 278872 251806 278924 251812
rect 278884 186998 278912 251806
rect 278976 231130 279004 260102
rect 279332 252816 279384 252822
rect 279332 252758 279384 252764
rect 279344 251870 279372 252758
rect 279332 251864 279384 251870
rect 279332 251806 279384 251812
rect 279436 246265 279464 451862
rect 280172 409154 280200 598946
rect 280252 555484 280304 555490
rect 280252 555426 280304 555432
rect 280264 464370 280292 555426
rect 280816 536489 280844 702918
rect 283852 700330 283880 703520
rect 285588 702840 285640 702846
rect 285588 702782 285640 702788
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 281540 603152 281592 603158
rect 281540 603094 281592 603100
rect 280802 536480 280858 536489
rect 280802 536415 280858 536424
rect 280252 464364 280304 464370
rect 280252 464306 280304 464312
rect 280252 454708 280304 454714
rect 280252 454650 280304 454656
rect 280160 409148 280212 409154
rect 280160 409090 280212 409096
rect 280160 383716 280212 383722
rect 280160 383658 280212 383664
rect 280172 278730 280200 383658
rect 280264 317422 280292 454650
rect 280436 419552 280488 419558
rect 280436 419494 280488 419500
rect 280344 400240 280396 400246
rect 280344 400182 280396 400188
rect 280356 352578 280384 400182
rect 280448 380769 280476 419494
rect 281552 419490 281580 603094
rect 284300 592680 284352 592686
rect 284300 592622 284352 592628
rect 283564 572756 283616 572762
rect 283564 572698 283616 572704
rect 281632 567860 281684 567866
rect 281632 567802 281684 567808
rect 281540 419484 281592 419490
rect 281540 419426 281592 419432
rect 281552 418810 281580 419426
rect 281540 418804 281592 418810
rect 281540 418746 281592 418752
rect 281540 389836 281592 389842
rect 281540 389778 281592 389784
rect 280434 380760 280490 380769
rect 280434 380695 280490 380704
rect 280344 352572 280396 352578
rect 280344 352514 280396 352520
rect 280252 317416 280304 317422
rect 280252 317358 280304 317364
rect 280252 291848 280304 291854
rect 280252 291790 280304 291796
rect 280160 278724 280212 278730
rect 280160 278666 280212 278672
rect 280158 271144 280214 271153
rect 280158 271079 280214 271088
rect 279422 246256 279478 246265
rect 279422 246191 279478 246200
rect 278964 231124 279016 231130
rect 278964 231066 279016 231072
rect 280172 227633 280200 271079
rect 280158 227624 280214 227633
rect 280158 227559 280214 227568
rect 278872 186992 278924 186998
rect 278872 186934 278924 186940
rect 280172 115258 280200 227559
rect 280264 198014 280292 291790
rect 280356 270502 280384 352514
rect 280436 317416 280488 317422
rect 280436 317358 280488 317364
rect 280448 316062 280476 317358
rect 280436 316056 280488 316062
rect 280436 315998 280488 316004
rect 280344 270496 280396 270502
rect 280344 270438 280396 270444
rect 280344 269816 280396 269822
rect 280344 269758 280396 269764
rect 280356 229090 280384 269758
rect 280448 268394 280476 315998
rect 281552 314702 281580 389778
rect 281644 389162 281672 567802
rect 282920 538280 282972 538286
rect 282920 538222 282972 538228
rect 281724 534744 281776 534750
rect 281724 534686 281776 534692
rect 281632 389156 281684 389162
rect 281632 389098 281684 389104
rect 281632 382968 281684 382974
rect 281632 382910 281684 382916
rect 281540 314696 281592 314702
rect 281540 314638 281592 314644
rect 281540 300212 281592 300218
rect 281540 300154 281592 300160
rect 280436 268388 280488 268394
rect 280436 268330 280488 268336
rect 281448 246356 281500 246362
rect 281448 246298 281500 246304
rect 281460 245682 281488 246298
rect 280804 245676 280856 245682
rect 280804 245618 280856 245624
rect 281448 245676 281500 245682
rect 281448 245618 281500 245624
rect 280344 229084 280396 229090
rect 280344 229026 280396 229032
rect 280252 198008 280304 198014
rect 280252 197950 280304 197956
rect 280816 124166 280844 245618
rect 280896 140888 280948 140894
rect 280896 140830 280948 140836
rect 280804 124160 280856 124166
rect 280804 124102 280856 124108
rect 280160 115252 280212 115258
rect 280160 115194 280212 115200
rect 280804 103556 280856 103562
rect 280908 103514 280936 140830
rect 280856 103504 280936 103514
rect 280804 103498 280936 103504
rect 280816 103486 280936 103498
rect 278778 77208 278834 77217
rect 278778 77143 278834 77152
rect 280066 77208 280122 77217
rect 280066 77143 280122 77152
rect 280080 76566 280108 77143
rect 280068 76560 280120 76566
rect 280068 76502 280120 76508
rect 278780 32428 278832 32434
rect 278780 32370 278832 32376
rect 278792 16574 278820 32370
rect 278792 16546 279096 16574
rect 278044 4412 278096 4418
rect 278044 4354 278096 4360
rect 276756 3460 276808 3466
rect 277964 3454 278360 3482
rect 276756 3402 276808 3408
rect 276952 598 277164 626
rect 276952 490 276980 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 462 276980 490
rect 277136 480 277164 598
rect 278332 480 278360 3454
rect 279068 490 279096 16546
rect 280712 11756 280764 11762
rect 280712 11698 280764 11704
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 11698
rect 280816 7614 280844 103486
rect 281552 102814 281580 300154
rect 281644 274650 281672 382910
rect 281736 380866 281764 534686
rect 281816 532024 281868 532030
rect 281816 531966 281868 531972
rect 281828 456929 281856 531966
rect 281814 456920 281870 456929
rect 281814 456855 281870 456864
rect 281828 412622 281856 456855
rect 281816 412616 281868 412622
rect 281816 412558 281868 412564
rect 281816 405748 281868 405754
rect 281816 405690 281868 405696
rect 281724 380860 281776 380866
rect 281724 380802 281776 380808
rect 281828 368490 281856 405690
rect 281816 368484 281868 368490
rect 281816 368426 281868 368432
rect 281828 354674 281856 368426
rect 281736 354646 281856 354674
rect 281736 281450 281764 354646
rect 281816 314696 281868 314702
rect 281816 314638 281868 314644
rect 281724 281444 281776 281450
rect 281724 281386 281776 281392
rect 281828 276690 281856 314638
rect 282932 311137 282960 538222
rect 283102 450120 283158 450129
rect 283102 450055 283158 450064
rect 283010 385656 283066 385665
rect 283010 385591 283066 385600
rect 282918 311128 282974 311137
rect 282918 311063 282974 311072
rect 282920 307760 282972 307766
rect 282920 307702 282972 307708
rect 282932 306406 282960 307702
rect 282920 306400 282972 306406
rect 282920 306342 282972 306348
rect 281816 276684 281868 276690
rect 281816 276626 281868 276632
rect 281632 274644 281684 274650
rect 281632 274586 281684 274592
rect 282932 273873 282960 306342
rect 282918 273864 282974 273873
rect 282918 273799 282974 273808
rect 281632 272536 281684 272542
rect 281632 272478 281684 272484
rect 281644 151201 281672 272478
rect 282920 267164 282972 267170
rect 282920 267106 282972 267112
rect 282932 266422 282960 267106
rect 282920 266416 282972 266422
rect 282920 266358 282972 266364
rect 281722 262848 281778 262857
rect 281722 262783 281778 262792
rect 281736 224262 281764 262783
rect 281816 233232 281868 233238
rect 281816 233174 281868 233180
rect 281828 231878 281856 233174
rect 281816 231872 281868 231878
rect 281816 231814 281868 231820
rect 281724 224256 281776 224262
rect 281724 224198 281776 224204
rect 281828 215286 281856 231814
rect 281816 215280 281868 215286
rect 281816 215222 281868 215228
rect 282932 154562 282960 266358
rect 283024 240106 283052 385591
rect 283116 307766 283144 450055
rect 283196 416832 283248 416838
rect 283196 416774 283248 416780
rect 283208 378146 283236 416774
rect 283576 391270 283604 572698
rect 283656 417444 283708 417450
rect 283656 417386 283708 417392
rect 283668 416838 283696 417386
rect 283656 416832 283708 416838
rect 283656 416774 283708 416780
rect 283564 391264 283616 391270
rect 283564 391206 283616 391212
rect 284312 387802 284340 592622
rect 284392 583024 284444 583030
rect 284392 582966 284444 582972
rect 284404 460934 284432 582966
rect 285600 536858 285628 702782
rect 288714 604752 288770 604761
rect 288714 604687 288770 604696
rect 289726 604752 289782 604761
rect 289726 604687 289782 604696
rect 287060 597644 287112 597650
rect 287060 597586 287112 597592
rect 285680 594108 285732 594114
rect 285680 594050 285732 594056
rect 285692 593434 285720 594050
rect 285680 593428 285732 593434
rect 285680 593370 285732 593376
rect 285588 536852 285640 536858
rect 285588 536794 285640 536800
rect 285692 466585 285720 593370
rect 285864 542360 285916 542366
rect 285864 542302 285916 542308
rect 285678 466576 285734 466585
rect 285678 466511 285734 466520
rect 285678 462904 285734 462913
rect 285678 462839 285734 462848
rect 284404 460906 284524 460934
rect 284496 456113 284524 460906
rect 284482 456104 284538 456113
rect 284482 456039 284538 456048
rect 284392 427100 284444 427106
rect 284392 427042 284444 427048
rect 284404 426494 284432 427042
rect 284392 426488 284444 426494
rect 284392 426430 284444 426436
rect 284300 387796 284352 387802
rect 284300 387738 284352 387744
rect 283196 378140 283248 378146
rect 283196 378082 283248 378088
rect 283104 307760 283156 307766
rect 283104 307702 283156 307708
rect 283208 254658 283236 378082
rect 284298 373280 284354 373289
rect 284298 373215 284354 373224
rect 283196 254652 283248 254658
rect 283196 254594 283248 254600
rect 283102 253872 283158 253881
rect 283102 253807 283158 253816
rect 283116 252618 283144 253807
rect 283104 252612 283156 252618
rect 283104 252554 283156 252560
rect 283012 240100 283064 240106
rect 283012 240042 283064 240048
rect 283116 195294 283144 252554
rect 284312 242185 284340 373215
rect 284404 252822 284432 426430
rect 284496 320249 284524 456039
rect 284482 320240 284538 320249
rect 284482 320175 284538 320184
rect 284496 267170 284524 320175
rect 284944 287700 284996 287706
rect 284944 287642 284996 287648
rect 284484 267164 284536 267170
rect 284484 267106 284536 267112
rect 284482 262304 284538 262313
rect 284482 262239 284538 262248
rect 284392 252816 284444 252822
rect 284392 252758 284444 252764
rect 284298 242176 284354 242185
rect 284298 242111 284354 242120
rect 283104 195288 283156 195294
rect 283104 195230 283156 195236
rect 282920 154556 282972 154562
rect 282920 154498 282972 154504
rect 281630 151192 281686 151201
rect 281630 151127 281686 151136
rect 282184 137284 282236 137290
rect 282184 137226 282236 137232
rect 281540 102808 281592 102814
rect 281540 102750 281592 102756
rect 281540 71052 281592 71058
rect 281540 70994 281592 71000
rect 280804 7608 280856 7614
rect 280804 7550 280856 7556
rect 281552 490 281580 70994
rect 282196 2990 282224 137226
rect 284312 89622 284340 242111
rect 284496 213217 284524 262239
rect 284482 213208 284538 213217
rect 284482 213143 284538 213152
rect 284956 144226 284984 287642
rect 285126 263528 285182 263537
rect 285126 263463 285182 263472
rect 285140 262313 285168 263463
rect 285126 262304 285182 262313
rect 285126 262239 285182 262248
rect 285692 244254 285720 462839
rect 285772 442264 285824 442270
rect 285772 442206 285824 442212
rect 285784 264246 285812 442206
rect 285876 419558 285904 542302
rect 287072 472666 287100 597586
rect 287152 587920 287204 587926
rect 287152 587862 287204 587868
rect 287060 472660 287112 472666
rect 287060 472602 287112 472608
rect 287060 471300 287112 471306
rect 287060 471242 287112 471248
rect 285864 419552 285916 419558
rect 285864 419494 285916 419500
rect 285864 418804 285916 418810
rect 285864 418746 285916 418752
rect 285876 358766 285904 418746
rect 285864 358760 285916 358766
rect 285864 358702 285916 358708
rect 285772 264240 285824 264246
rect 285772 264182 285824 264188
rect 285772 259480 285824 259486
rect 285772 259422 285824 259428
rect 285784 254590 285812 259422
rect 285876 257281 285904 358702
rect 287072 300150 287100 471242
rect 287164 451926 287192 587862
rect 288624 565888 288676 565894
rect 288624 565830 288676 565836
rect 288440 556232 288492 556238
rect 288440 556174 288492 556180
rect 287612 472660 287664 472666
rect 287612 472602 287664 472608
rect 287624 472161 287652 472602
rect 287610 472152 287666 472161
rect 287610 472087 287666 472096
rect 288348 456068 288400 456074
rect 288348 456010 288400 456016
rect 288360 455569 288388 456010
rect 287334 455560 287390 455569
rect 287334 455495 287390 455504
rect 288346 455560 288402 455569
rect 288346 455495 288402 455504
rect 287242 454744 287298 454753
rect 287242 454679 287298 454688
rect 287152 451920 287204 451926
rect 287152 451862 287204 451868
rect 287150 301064 287206 301073
rect 287150 300999 287206 301008
rect 287060 300144 287112 300150
rect 287060 300086 287112 300092
rect 285956 294636 286008 294642
rect 285956 294578 286008 294584
rect 285862 257272 285918 257281
rect 285862 257207 285918 257216
rect 285772 254584 285824 254590
rect 285772 254526 285824 254532
rect 285680 244248 285732 244254
rect 285680 244190 285732 244196
rect 285680 218816 285732 218822
rect 285680 218758 285732 218764
rect 285128 217320 285180 217326
rect 285128 217262 285180 217268
rect 285140 216753 285168 217262
rect 285126 216744 285182 216753
rect 285126 216679 285182 216688
rect 285140 200114 285168 216679
rect 285048 200086 285168 200114
rect 284944 144220 284996 144226
rect 284944 144162 284996 144168
rect 284944 119400 284996 119406
rect 284944 119342 284996 119348
rect 284392 107636 284444 107642
rect 284392 107578 284444 107584
rect 284404 106962 284432 107578
rect 284392 106956 284444 106962
rect 284392 106898 284444 106904
rect 284300 89616 284352 89622
rect 284300 89558 284352 89564
rect 284312 89010 284340 89558
rect 284300 89004 284352 89010
rect 284300 88946 284352 88952
rect 284956 74497 284984 119342
rect 285048 107642 285076 200086
rect 285036 107636 285088 107642
rect 285036 107578 285088 107584
rect 285692 104854 285720 218758
rect 285784 144129 285812 254526
rect 285968 219366 285996 294578
rect 285956 219360 286008 219366
rect 285956 219302 286008 219308
rect 285968 218822 285996 219302
rect 285956 218816 286008 218822
rect 285956 218758 286008 218764
rect 285770 144120 285826 144129
rect 285770 144055 285826 144064
rect 285680 104848 285732 104854
rect 285680 104790 285732 104796
rect 287164 78577 287192 300999
rect 287256 263634 287284 454679
rect 287244 263628 287296 263634
rect 287244 263570 287296 263576
rect 287256 145586 287284 263570
rect 287348 259486 287376 455495
rect 288452 367810 288480 556174
rect 288530 463720 288586 463729
rect 288530 463655 288586 463664
rect 288440 367804 288492 367810
rect 288440 367746 288492 367752
rect 288440 295384 288492 295390
rect 288440 295326 288492 295332
rect 287336 259480 287388 259486
rect 287336 259422 287388 259428
rect 287244 145580 287296 145586
rect 287244 145522 287296 145528
rect 287704 140820 287756 140826
rect 287704 140762 287756 140768
rect 287150 78568 287206 78577
rect 287150 78503 287206 78512
rect 284942 74488 284998 74497
rect 284942 74423 284998 74432
rect 284956 73273 284984 74423
rect 284298 73264 284354 73273
rect 284298 73199 284354 73208
rect 284942 73264 284998 73273
rect 284942 73199 284998 73208
rect 282184 2984 282236 2990
rect 282184 2926 282236 2932
rect 283104 2984 283156 2990
rect 283104 2926 283156 2932
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 2926
rect 284312 480 284340 73199
rect 287060 68332 287112 68338
rect 287060 68274 287112 68280
rect 286324 50380 286376 50386
rect 286324 50322 286376 50328
rect 284392 18624 284444 18630
rect 284392 18566 284444 18572
rect 284404 16574 284432 18566
rect 284404 16546 284984 16574
rect 284956 490 284984 16546
rect 286336 6186 286364 50322
rect 287072 16574 287100 68274
rect 287072 16546 287376 16574
rect 286324 6180 286376 6186
rect 286324 6122 286376 6128
rect 286600 3460 286652 3466
rect 286600 3402 286652 3408
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 3402
rect 287348 490 287376 16546
rect 287716 3058 287744 140762
rect 288452 79393 288480 295326
rect 288544 264217 288572 463655
rect 288636 378049 288664 565830
rect 288728 439550 288756 604687
rect 289740 604518 289768 604687
rect 289728 604512 289780 604518
rect 289728 604454 289780 604460
rect 299480 600364 299532 600370
rect 299480 600306 299532 600312
rect 293960 596828 294012 596834
rect 293960 596770 294012 596776
rect 292580 589960 292632 589966
rect 292580 589902 292632 589908
rect 289912 568608 289964 568614
rect 289912 568550 289964 568556
rect 289728 566500 289780 566506
rect 289728 566442 289780 566448
rect 289740 565894 289768 566442
rect 289728 565888 289780 565894
rect 289728 565830 289780 565836
rect 289818 459640 289874 459649
rect 289818 459575 289874 459584
rect 288716 439544 288768 439550
rect 288716 439486 288768 439492
rect 288622 378040 288678 378049
rect 288622 377975 288678 377984
rect 288624 300892 288676 300898
rect 288624 300834 288676 300840
rect 288530 264208 288586 264217
rect 288530 264143 288586 264152
rect 288544 181490 288572 264143
rect 288532 181484 288584 181490
rect 288532 181426 288584 181432
rect 288636 140894 288664 300834
rect 288728 263537 288756 439486
rect 288714 263528 288770 263537
rect 288714 263463 288770 263472
rect 289832 245614 289860 459575
rect 289924 390561 289952 568550
rect 291200 536852 291252 536858
rect 291200 536794 291252 536800
rect 290004 465112 290056 465118
rect 290004 465054 290056 465060
rect 289910 390552 289966 390561
rect 289910 390487 289966 390496
rect 289924 389201 289952 390487
rect 289910 389192 289966 389201
rect 289910 389127 289966 389136
rect 290016 304298 290044 465054
rect 291212 384985 291240 536794
rect 291292 529236 291344 529242
rect 291292 529178 291344 529184
rect 291198 384976 291254 384985
rect 291198 384911 291254 384920
rect 291304 379506 291332 529178
rect 291382 472016 291438 472025
rect 291382 471951 291438 471960
rect 291396 427106 291424 471951
rect 291384 427100 291436 427106
rect 291384 427042 291436 427048
rect 291384 403028 291436 403034
rect 291384 402970 291436 402976
rect 291396 382265 291424 402970
rect 291476 391264 291528 391270
rect 291476 391206 291528 391212
rect 291382 382256 291438 382265
rect 291382 382191 291438 382200
rect 291292 379500 291344 379506
rect 291292 379442 291344 379448
rect 291198 311944 291254 311953
rect 291198 311879 291254 311888
rect 290004 304292 290056 304298
rect 290004 304234 290056 304240
rect 289912 293344 289964 293350
rect 289912 293286 289964 293292
rect 289820 245608 289872 245614
rect 289820 245550 289872 245556
rect 289832 244322 289860 245550
rect 289820 244316 289872 244322
rect 289820 244258 289872 244264
rect 288624 140888 288676 140894
rect 288624 140830 288676 140836
rect 289084 140072 289136 140078
rect 289084 140014 289136 140020
rect 288438 79384 288494 79393
rect 288438 79319 288494 79328
rect 288346 78568 288402 78577
rect 288346 78503 288402 78512
rect 288360 77994 288388 78503
rect 288348 77988 288400 77994
rect 288348 77930 288400 77936
rect 288440 19984 288492 19990
rect 288440 19926 288492 19932
rect 288452 16574 288480 19926
rect 288452 16546 289032 16574
rect 287704 3052 287756 3058
rect 287704 2994 287756 3000
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 16546
rect 289096 3534 289124 140014
rect 289924 119406 289952 293286
rect 291108 251864 291160 251870
rect 291108 251806 291160 251812
rect 291120 251258 291148 251806
rect 291108 251252 291160 251258
rect 291108 251194 291160 251200
rect 291120 233714 291148 251194
rect 290464 233708 290516 233714
rect 290464 233650 290516 233656
rect 291108 233708 291160 233714
rect 291108 233650 291160 233656
rect 290476 208350 290504 233650
rect 291120 233306 291148 233650
rect 291108 233300 291160 233306
rect 291108 233242 291160 233248
rect 290464 208344 290516 208350
rect 290464 208286 290516 208292
rect 289912 119400 289964 119406
rect 289912 119342 289964 119348
rect 291212 111110 291240 311879
rect 291290 308000 291346 308009
rect 291290 307935 291346 307944
rect 291304 117201 291332 307935
rect 291396 278050 291424 382191
rect 291488 376553 291516 391206
rect 291474 376544 291530 376553
rect 291474 376479 291530 376488
rect 292592 356726 292620 589902
rect 292672 460964 292724 460970
rect 292672 460906 292724 460912
rect 292580 356720 292632 356726
rect 292580 356662 292632 356668
rect 291476 339516 291528 339522
rect 291476 339458 291528 339464
rect 291488 284986 291516 339458
rect 292580 320884 292632 320890
rect 292580 320826 292632 320832
rect 291476 284980 291528 284986
rect 291476 284922 291528 284928
rect 292592 281518 292620 320826
rect 292684 319462 292712 460906
rect 293972 338745 294000 596770
rect 298100 591320 298152 591326
rect 298100 591262 298152 591268
rect 296810 453248 296866 453257
rect 296810 453183 296866 453192
rect 295338 437608 295394 437617
rect 295338 437543 295394 437552
rect 294052 342304 294104 342310
rect 294052 342246 294104 342252
rect 293958 338736 294014 338745
rect 293958 338671 294014 338680
rect 292672 319456 292724 319462
rect 292672 319398 292724 319404
rect 294064 287026 294092 342246
rect 294052 287020 294104 287026
rect 294052 286962 294104 286968
rect 292670 282160 292726 282169
rect 292670 282095 292726 282104
rect 292580 281512 292632 281518
rect 292580 281454 292632 281460
rect 291384 278044 291436 278050
rect 291384 277986 291436 277992
rect 291382 268560 291438 268569
rect 291382 268495 291438 268504
rect 291396 200122 291424 268495
rect 292684 220794 292712 282095
rect 295352 260137 295380 437543
rect 295522 309360 295578 309369
rect 295522 309295 295578 309304
rect 295432 264988 295484 264994
rect 295432 264930 295484 264936
rect 295338 260128 295394 260137
rect 295338 260063 295394 260072
rect 293960 244316 294012 244322
rect 293960 244258 294012 244264
rect 292672 220788 292724 220794
rect 292672 220730 292724 220736
rect 291384 200116 291436 200122
rect 291384 200058 291436 200064
rect 293972 164218 294000 244258
rect 293960 164212 294012 164218
rect 293960 164154 294012 164160
rect 294420 164212 294472 164218
rect 294420 164154 294472 164160
rect 294432 163538 294460 164154
rect 294420 163532 294472 163538
rect 294420 163474 294472 163480
rect 295340 127628 295392 127634
rect 295340 127570 295392 127576
rect 295352 126954 295380 127570
rect 295340 126948 295392 126954
rect 295340 126890 295392 126896
rect 291290 117192 291346 117201
rect 291290 117127 291346 117136
rect 291658 117192 291714 117201
rect 291658 117127 291714 117136
rect 291672 116618 291700 117127
rect 291660 116612 291712 116618
rect 291660 116554 291712 116560
rect 291200 111104 291252 111110
rect 291200 111046 291252 111052
rect 291212 110498 291240 111046
rect 291200 110492 291252 110498
rect 291200 110434 291252 110440
rect 291844 110492 291896 110498
rect 291844 110434 291896 110440
rect 291856 45626 291884 110434
rect 292672 76560 292724 76566
rect 292672 76502 292724 76508
rect 291936 46232 291988 46238
rect 291936 46174 291988 46180
rect 291844 45620 291896 45626
rect 291844 45562 291896 45568
rect 291200 25560 291252 25566
rect 291200 25502 291252 25508
rect 291212 16574 291240 25502
rect 291212 16546 291424 16574
rect 289084 3528 289136 3534
rect 289084 3470 289136 3476
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 290200 480 290228 3470
rect 291396 480 291424 16546
rect 291948 3534 291976 46174
rect 292684 16574 292712 76502
rect 295352 16574 295380 126890
rect 295444 124914 295472 264930
rect 295536 217326 295564 309295
rect 296718 306504 296774 306513
rect 296718 306439 296774 306448
rect 295524 217320 295576 217326
rect 295524 217262 295576 217268
rect 295432 124908 295484 124914
rect 295432 124850 295484 124856
rect 296732 37262 296760 306439
rect 296824 297430 296852 453183
rect 298112 371890 298140 591262
rect 298192 577516 298244 577522
rect 298192 577458 298244 577464
rect 298204 391338 298232 577458
rect 298284 420980 298336 420986
rect 298284 420922 298336 420928
rect 298192 391332 298244 391338
rect 298192 391274 298244 391280
rect 298100 371884 298152 371890
rect 298100 371826 298152 371832
rect 296812 297424 296864 297430
rect 296812 297366 296864 297372
rect 298100 294024 298152 294030
rect 298100 293966 298152 293972
rect 298112 188358 298140 293966
rect 298296 246362 298324 420922
rect 299492 329089 299520 600306
rect 299584 592686 299612 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 348804 703186 348832 703520
rect 348792 703180 348844 703186
rect 348792 703122 348844 703128
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 364996 702914 365024 703520
rect 364984 702908 365036 702914
rect 364984 702850 365036 702856
rect 397472 702794 397500 703520
rect 413664 703118 413692 703520
rect 413652 703112 413704 703118
rect 413652 703054 413704 703060
rect 429856 702982 429884 703520
rect 429844 702976 429896 702982
rect 429844 702918 429896 702924
rect 462332 702846 462360 703520
rect 397380 702766 397500 702794
rect 462320 702840 462372 702846
rect 462320 702782 462372 702788
rect 397380 702710 397408 702766
rect 397368 702704 397420 702710
rect 397368 702646 397420 702652
rect 478524 702642 478552 703520
rect 494808 702778 494836 703520
rect 494796 702772 494848 702778
rect 494796 702714 494848 702720
rect 478512 702636 478564 702642
rect 478512 702578 478564 702584
rect 527192 702574 527220 703520
rect 527180 702568 527232 702574
rect 527180 702510 527232 702516
rect 543476 702506 543504 703520
rect 543464 702500 543516 702506
rect 543464 702442 543516 702448
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 582840 700324 582892 700330
rect 582840 700266 582892 700272
rect 582470 697232 582526 697241
rect 582470 697167 582526 697176
rect 582378 617536 582434 617545
rect 582378 617471 582434 617480
rect 582392 606490 582420 617471
rect 582380 606484 582432 606490
rect 582380 606426 582432 606432
rect 299572 592680 299624 592686
rect 299572 592622 299624 592628
rect 582378 591016 582434 591025
rect 582378 590951 582434 590960
rect 582392 584458 582420 590951
rect 582380 584452 582432 584458
rect 582380 584394 582432 584400
rect 582378 577688 582434 577697
rect 582378 577623 582434 577632
rect 582392 537538 582420 577623
rect 582484 566506 582512 697167
rect 582562 683904 582618 683913
rect 582562 683839 582618 683848
rect 582576 570654 582604 683839
rect 582654 644056 582710 644065
rect 582654 643991 582710 644000
rect 582668 603673 582696 643991
rect 582746 630864 582802 630873
rect 582746 630799 582802 630808
rect 582760 607889 582788 630799
rect 582852 609249 582880 700266
rect 582930 670712 582986 670721
rect 582930 670647 582986 670656
rect 582838 609240 582894 609249
rect 582838 609175 582894 609184
rect 582746 607880 582802 607889
rect 582746 607815 582802 607824
rect 582840 604512 582892 604518
rect 582840 604454 582892 604460
rect 582654 603664 582710 603673
rect 582654 603599 582710 603608
rect 582746 601760 582802 601769
rect 582746 601695 582802 601704
rect 582656 593428 582708 593434
rect 582656 593370 582708 593376
rect 582564 570648 582616 570654
rect 582564 570590 582616 570596
rect 582472 566500 582524 566506
rect 582472 566442 582524 566448
rect 582470 537840 582526 537849
rect 582470 537775 582526 537784
rect 582380 537532 582432 537538
rect 582380 537474 582432 537480
rect 582484 528554 582512 537775
rect 582392 528526 582512 528554
rect 579802 484664 579858 484673
rect 579802 484599 579858 484608
rect 579816 484362 579844 484599
rect 579804 484356 579856 484362
rect 579804 484298 579856 484304
rect 302240 474836 302292 474842
rect 302240 474778 302292 474784
rect 299572 466472 299624 466478
rect 299572 466414 299624 466420
rect 299478 329080 299534 329089
rect 299478 329015 299534 329024
rect 299480 293276 299532 293282
rect 299480 293218 299532 293224
rect 298284 246356 298336 246362
rect 298284 246298 298336 246304
rect 298100 188352 298152 188358
rect 298100 188294 298152 188300
rect 299492 155242 299520 293218
rect 299584 251870 299612 466414
rect 302252 287706 302280 474778
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456074 580212 458079
rect 580172 456068 580224 456074
rect 580172 456010 580224 456016
rect 582392 418810 582420 528526
rect 582668 511329 582696 593370
rect 582760 524521 582788 601695
rect 582852 564369 582880 604454
rect 582838 564360 582894 564369
rect 582838 564295 582894 564304
rect 582944 538257 582972 670647
rect 582930 538248 582986 538257
rect 582930 538183 582986 538192
rect 582746 524512 582802 524521
rect 582746 524447 582802 524456
rect 582654 511320 582710 511329
rect 582654 511255 582710 511264
rect 582472 472660 582524 472666
rect 582472 472602 582524 472608
rect 582380 418804 582432 418810
rect 582380 418746 582432 418752
rect 582378 418296 582434 418305
rect 582378 418231 582434 418240
rect 582392 391270 582420 418231
rect 582484 404977 582512 472602
rect 582654 471472 582710 471481
rect 582654 471407 582710 471416
rect 582564 427100 582616 427106
rect 582564 427042 582616 427048
rect 582470 404968 582526 404977
rect 582470 404903 582526 404912
rect 582380 391264 582432 391270
rect 582380 391206 582432 391212
rect 582380 387116 582432 387122
rect 582380 387058 582432 387064
rect 582392 378457 582420 387058
rect 582378 378448 582434 378457
rect 582378 378383 582434 378392
rect 582470 365120 582526 365129
rect 582470 365055 582526 365064
rect 302330 305008 302386 305017
rect 302330 304943 302386 304952
rect 302240 287700 302292 287706
rect 302240 287642 302292 287648
rect 299572 251864 299624 251870
rect 299572 251806 299624 251812
rect 299480 155236 299532 155242
rect 299480 155178 299532 155184
rect 298744 144220 298796 144226
rect 298744 144162 298796 144168
rect 298100 47592 298152 47598
rect 298100 47534 298152 47540
rect 296812 45620 296864 45626
rect 296812 45562 296864 45568
rect 296720 37256 296772 37262
rect 296720 37198 296772 37204
rect 296824 16574 296852 45562
rect 298008 37256 298060 37262
rect 298008 37198 298060 37204
rect 298020 36582 298048 37198
rect 298008 36576 298060 36582
rect 298008 36518 298060 36524
rect 292684 16546 293264 16574
rect 295352 16546 295656 16574
rect 296824 16546 297312 16574
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 292580 3052 292632 3058
rect 292580 2994 292632 3000
rect 292592 480 292620 2994
rect 293236 490 293264 16546
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 293512 598 293724 626
rect 293512 490 293540 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 462 293540 490
rect 293696 480 293724 598
rect 294892 480 294920 3470
rect 295628 490 295656 16546
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 16546
rect 298112 490 298140 47534
rect 298756 3534 298784 144162
rect 299480 129056 299532 129062
rect 299480 128998 299532 129004
rect 298744 3528 298796 3534
rect 298744 3470 298796 3476
rect 299492 2650 299520 128998
rect 302344 126954 302372 304943
rect 582378 302832 582434 302841
rect 582378 302767 582434 302776
rect 303620 300144 303672 300150
rect 303620 300086 303672 300092
rect 303632 172514 303660 300086
rect 580172 278044 580224 278050
rect 580172 277986 580224 277992
rect 580184 272241 580212 277986
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 580920 257378 580948 258839
rect 580908 257372 580960 257378
rect 580908 257314 580960 257320
rect 580264 233300 580316 233306
rect 580264 233242 580316 233248
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 580276 219065 580304 233242
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580170 192536 580226 192545
rect 580170 192471 580172 192480
rect 580224 192471 580226 192480
rect 580172 192442 580224 192448
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178702 580212 179143
rect 580172 178696 580224 178702
rect 580172 178638 580224 178644
rect 341524 173188 341576 173194
rect 341524 173130 341576 173136
rect 303620 172508 303672 172514
rect 303620 172450 303672 172456
rect 304080 172508 304132 172514
rect 304080 172450 304132 172456
rect 304092 171834 304120 172450
rect 304080 171828 304132 171834
rect 304080 171770 304132 171776
rect 320180 171828 320232 171834
rect 320180 171770 320232 171776
rect 316038 159352 316094 159361
rect 316038 159287 316094 159296
rect 303618 157448 303674 157457
rect 303618 157383 303674 157392
rect 302884 133952 302936 133958
rect 302884 133894 302936 133900
rect 302332 126948 302384 126954
rect 302332 126890 302384 126896
rect 299570 39264 299626 39273
rect 299570 39199 299626 39208
rect 299584 16574 299612 39199
rect 300858 26888 300914 26897
rect 300858 26823 300914 26832
rect 300872 16574 300900 26823
rect 299584 16546 299704 16574
rect 300872 16546 301544 16574
rect 299480 2644 299532 2650
rect 299480 2586 299532 2592
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 16546
rect 300768 2644 300820 2650
rect 300768 2586 300820 2592
rect 300780 480 300808 2586
rect 301516 490 301544 16546
rect 302896 15910 302924 133894
rect 302974 21312 303030 21321
rect 302974 21247 303030 21256
rect 302884 15904 302936 15910
rect 302884 15846 302936 15852
rect 302884 14544 302936 14550
rect 302884 14486 302936 14492
rect 302896 3482 302924 14486
rect 302988 4010 303016 21247
rect 303632 16574 303660 157383
rect 305644 149728 305696 149734
rect 305644 149670 305696 149676
rect 304264 116612 304316 116618
rect 304264 116554 304316 116560
rect 303632 16546 303936 16574
rect 302976 4004 303028 4010
rect 302976 3946 303028 3952
rect 302896 3454 303200 3482
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 3454
rect 303908 490 303936 16546
rect 304276 4049 304304 116554
rect 305656 5574 305684 149670
rect 313280 122120 313332 122126
rect 313280 122062 313332 122068
rect 309784 102808 309836 102814
rect 309784 102750 309836 102756
rect 307024 84924 307076 84930
rect 307024 84866 307076 84872
rect 305644 5568 305696 5574
rect 305644 5510 305696 5516
rect 304262 4040 304318 4049
rect 304262 3975 304318 3984
rect 306748 4004 306800 4010
rect 306748 3946 306800 3952
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3470
rect 306760 480 306788 3946
rect 307036 3534 307064 84866
rect 309140 44872 309192 44878
rect 309140 44814 309192 44820
rect 309152 16574 309180 44814
rect 309796 18018 309824 102750
rect 311900 35216 311952 35222
rect 311900 35158 311952 35164
rect 309784 18012 309836 18018
rect 309784 17954 309836 17960
rect 311912 16574 311940 35158
rect 313292 16574 313320 122062
rect 309152 16546 309824 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 309048 5568 309100 5574
rect 309048 5510 309100 5516
rect 307942 4040 307998 4049
rect 307942 3975 307998 3984
rect 307024 3528 307076 3534
rect 307024 3470 307076 3476
rect 307956 480 307984 3975
rect 309060 480 309088 5510
rect 309796 490 309824 16546
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 3470
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 314660 15904 314712 15910
rect 314660 15846 314712 15852
rect 314672 490 314700 15846
rect 316052 3482 316080 159287
rect 317420 148368 317472 148374
rect 317420 148310 317472 148316
rect 316132 18012 316184 18018
rect 316132 17954 316184 17960
rect 316144 3602 316172 17954
rect 317432 6914 317460 148310
rect 318064 74588 318116 74594
rect 318064 74530 318116 74536
rect 318076 16574 318104 74530
rect 318076 16546 318196 16574
rect 317432 6886 318104 6914
rect 316132 3596 316184 3602
rect 316132 3538 316184 3544
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 316052 3454 316264 3482
rect 314856 598 315068 626
rect 314856 490 314884 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 462 314884 490
rect 315040 480 315068 598
rect 316236 480 316264 3454
rect 317340 480 317368 3538
rect 318076 490 318104 6886
rect 318168 3262 318196 16546
rect 320192 3534 320220 171770
rect 323584 150476 323636 150482
rect 323584 150418 323636 150424
rect 322204 99408 322256 99414
rect 322204 99350 322256 99356
rect 320272 54528 320324 54534
rect 320272 54470 320324 54476
rect 320284 16574 320312 54470
rect 322216 18630 322244 99350
rect 322296 63572 322348 63578
rect 322296 63514 322348 63520
rect 322204 18624 322256 18630
rect 322204 18566 322256 18572
rect 320284 16546 320496 16574
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 320180 3528 320232 3534
rect 320180 3470 320232 3476
rect 318156 3256 318208 3262
rect 318156 3198 318208 3204
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3470
rect 320468 490 320496 16546
rect 322112 3256 322164 3262
rect 322112 3198 322164 3204
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 3198
rect 322308 3194 322336 63514
rect 322940 43444 322992 43450
rect 322940 43386 322992 43392
rect 322296 3188 322348 3194
rect 322296 3130 322348 3136
rect 322952 490 322980 43386
rect 323596 4010 323624 150418
rect 327080 145648 327132 145654
rect 327080 145590 327132 145596
rect 324412 112464 324464 112470
rect 324412 112406 324464 112412
rect 324424 11762 324452 112406
rect 327092 16574 327120 145590
rect 333980 135924 334032 135930
rect 333980 135866 334032 135872
rect 331220 93152 331272 93158
rect 331220 93094 331272 93100
rect 327092 16546 328040 16574
rect 324412 11756 324464 11762
rect 324412 11698 324464 11704
rect 325608 11756 325660 11762
rect 325608 11698 325660 11704
rect 323584 4004 323636 4010
rect 323584 3946 323636 3952
rect 324412 3188 324464 3194
rect 324412 3130 324464 3136
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 3130
rect 325620 480 325648 11698
rect 326804 4004 326856 4010
rect 326804 3946 326856 3952
rect 326816 480 326844 3946
rect 328012 480 328040 16546
rect 330392 7608 330444 7614
rect 330392 7550 330444 7556
rect 329196 6180 329248 6186
rect 329196 6122 329248 6128
rect 329208 480 329236 6122
rect 330404 480 330432 7550
rect 331232 490 331260 93094
rect 332600 18624 332652 18630
rect 332600 18566 332652 18572
rect 332612 16574 332640 18566
rect 332612 16546 332732 16574
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 16546
rect 333992 3074 334020 135866
rect 338118 87544 338174 87553
rect 338118 87479 338174 87488
rect 335358 65512 335414 65521
rect 335358 65447 335414 65456
rect 334072 40724 334124 40730
rect 334072 40666 334124 40672
rect 334084 16574 334112 40666
rect 335372 16574 335400 65447
rect 336740 17264 336792 17270
rect 336740 17206 336792 17212
rect 336752 16574 336780 17206
rect 338132 16574 338160 87479
rect 339500 82884 339552 82890
rect 339500 82826 339552 82832
rect 334084 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 333900 3046 334020 3074
rect 333900 480 333928 3046
rect 334636 490 334664 16546
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 16546
rect 337028 490 337056 16546
rect 337304 598 337516 626
rect 337304 490 337332 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 462 337332 490
rect 337488 480 337516 598
rect 338684 480 338712 16546
rect 339512 490 339540 82826
rect 340972 13116 341024 13122
rect 340972 13058 341024 13064
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 13058
rect 341536 3369 341564 173130
rect 342260 153876 342312 153882
rect 342260 153818 342312 153824
rect 341522 3360 341578 3369
rect 341522 3295 341578 3304
rect 342272 3074 342300 153818
rect 351920 126268 351972 126274
rect 351920 126210 351972 126216
rect 345664 109744 345716 109750
rect 345664 109686 345716 109692
rect 345020 77988 345072 77994
rect 345020 77930 345072 77936
rect 343640 36576 343692 36582
rect 343640 36518 343692 36524
rect 343652 16574 343680 36518
rect 345032 16574 345060 77930
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 342904 10328 342956 10334
rect 342904 10270 342956 10276
rect 342180 3046 342300 3074
rect 342180 480 342208 3046
rect 342916 490 342944 10270
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 16546
rect 345308 490 345336 16546
rect 345676 3194 345704 109686
rect 349160 106956 349212 106962
rect 349160 106898 349212 106904
rect 349172 5574 349200 106898
rect 346952 5568 347004 5574
rect 346952 5510 347004 5516
rect 349160 5568 349212 5574
rect 349160 5510 349212 5516
rect 345664 3188 345716 3194
rect 345664 3130 345716 3136
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 5510
rect 351644 3528 351696 3534
rect 351644 3470 351696 3476
rect 350446 3360 350502 3369
rect 350446 3295 350502 3304
rect 348056 3256 348108 3262
rect 348056 3198 348108 3204
rect 348068 480 348096 3198
rect 349252 3188 349304 3194
rect 349252 3130 349304 3136
rect 349264 480 349292 3130
rect 350460 480 350488 3295
rect 351656 480 351684 3470
rect 351932 3262 351960 126210
rect 580264 89752 580316 89758
rect 580264 89694 580316 89700
rect 353298 82104 353354 82113
rect 353298 82039 353354 82048
rect 353312 3534 353340 82039
rect 580276 73001 580304 89694
rect 580262 72992 580318 73001
rect 580262 72927 580318 72936
rect 580172 49020 580224 49026
rect 580172 48962 580224 48968
rect 580184 46345 580212 48962
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 353300 3528 353352 3534
rect 582392 3482 582420 302767
rect 582484 251841 582512 365055
rect 582576 351937 582604 427042
rect 582668 417450 582696 471407
rect 582746 431624 582802 431633
rect 582746 431559 582802 431568
rect 582656 417444 582708 417450
rect 582656 417386 582708 417392
rect 582760 390561 582788 431559
rect 582746 390552 582802 390561
rect 582746 390487 582802 390496
rect 582562 351928 582618 351937
rect 582562 351863 582618 351872
rect 582654 312080 582710 312089
rect 582654 312015 582710 312024
rect 582564 289876 582616 289882
rect 582564 289818 582616 289824
rect 582470 251832 582526 251841
rect 582470 251767 582526 251776
rect 582470 248432 582526 248441
rect 582470 248367 582526 248376
rect 582484 245585 582512 248367
rect 582470 245576 582526 245585
rect 582470 245511 582526 245520
rect 582472 200796 582524 200802
rect 582472 200738 582524 200744
rect 353300 3470 353352 3476
rect 582208 3454 582420 3482
rect 581000 3324 581052 3330
rect 581000 3266 581052 3272
rect 351920 3256 351972 3262
rect 351920 3198 351972 3204
rect 581012 480 581040 3266
rect 582208 480 582236 3454
rect 582484 3210 582512 200738
rect 582576 3330 582604 289818
rect 582668 251190 582696 312015
rect 582656 251184 582708 251190
rect 582656 251126 582708 251132
rect 582656 235272 582708 235278
rect 582656 235214 582708 235220
rect 582668 152697 582696 235214
rect 583024 175296 583076 175302
rect 583024 175238 583076 175244
rect 582748 169788 582800 169794
rect 582748 169730 582800 169736
rect 582654 152688 582710 152697
rect 582654 152623 582710 152632
rect 582654 138680 582710 138689
rect 582654 138615 582710 138624
rect 582668 19825 582696 138615
rect 582760 59673 582788 169730
rect 582838 165880 582894 165889
rect 582838 165815 582894 165824
rect 582852 124166 582880 165815
rect 582932 163532 582984 163538
rect 582932 163474 582984 163480
rect 582944 126041 582972 163474
rect 583036 139369 583064 175238
rect 583114 146432 583170 146441
rect 583114 146367 583170 146376
rect 583022 139360 583078 139369
rect 583022 139295 583078 139304
rect 582930 126032 582986 126041
rect 582930 125967 582986 125976
rect 582840 124160 582892 124166
rect 582840 124102 582892 124108
rect 583128 112849 583156 146367
rect 583114 112840 583170 112849
rect 583114 112775 583170 112784
rect 583022 99512 583078 99521
rect 583022 99447 583078 99456
rect 582840 89004 582892 89010
rect 582840 88946 582892 88952
rect 582746 59664 582802 59673
rect 582746 59599 582802 59608
rect 582654 19816 582710 19825
rect 582654 19751 582710 19760
rect 582852 6633 582880 88946
rect 582932 80708 582984 80714
rect 582932 80650 582984 80656
rect 582944 33153 582972 80650
rect 583036 73166 583064 99447
rect 583024 73160 583076 73166
rect 583024 73102 583076 73108
rect 582930 33144 582986 33153
rect 582930 33079 582986 33088
rect 582838 6624 582894 6633
rect 582838 6559 582894 6568
rect 582564 3324 582616 3330
rect 582564 3266 582616 3272
rect 582484 3182 583432 3210
rect 583404 480 583432 3182
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 3330 579944 3386 580000
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 566888 3478 566944
rect 2778 553852 2834 553888
rect 2778 553832 2780 553852
rect 2780 553832 2832 553852
rect 2832 553832 2834 553852
rect 55034 582528 55090 582584
rect 15842 541048 15898 541104
rect 3146 527856 3202 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3422 501744 3478 501800
rect 3330 475632 3386 475688
rect 3422 462576 3478 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3514 410488 3570 410544
rect 3422 397432 3478 397488
rect 3422 377304 3478 377360
rect 3514 371320 3570 371376
rect 7562 391856 7618 391912
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 3146 345344 3202 345400
rect 19338 342896 19394 342952
rect 8298 335960 8354 336016
rect 4066 319232 4122 319288
rect 3422 306176 3478 306232
rect 3422 293120 3478 293176
rect 3422 290400 3478 290456
rect 5538 300056 5594 300112
rect 4158 294480 4214 294536
rect 3422 267144 3478 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 2778 215872 2834 215928
rect 3514 214940 3570 214976
rect 3514 214920 3516 214940
rect 3516 214920 3568 214940
rect 3568 214920 3570 214940
rect 3514 201864 3570 201920
rect 3422 188808 3478 188864
rect 3422 162832 3478 162888
rect 2870 136720 2926 136776
rect 2870 110608 2926 110664
rect 3054 97552 3110 97608
rect 3330 84632 3386 84688
rect 3514 71576 3570 71632
rect 3422 58520 3478 58576
rect 3514 45464 3570 45520
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 4250 149776 4306 149832
rect 3422 6432 3478 6488
rect 12438 334600 12494 334656
rect 11058 298696 11114 298752
rect 11150 25472 11206 25528
rect 16578 330384 16634 330440
rect 15198 320728 15254 320784
rect 13818 236000 13874 236056
rect 17958 302232 18014 302288
rect 20718 331744 20774 331800
rect 22098 327120 22154 327176
rect 26238 323584 26294 323640
rect 24858 291760 24914 291816
rect 22742 235184 22798 235240
rect 28998 301416 29054 301472
rect 27618 297336 27674 297392
rect 27710 152360 27766 152416
rect 34518 328480 34574 328536
rect 39946 389136 40002 389192
rect 42706 437552 42762 437608
rect 41326 337320 41382 337376
rect 38658 233824 38714 233880
rect 35990 202136 36046 202192
rect 41418 325760 41474 325816
rect 52366 456864 52422 456920
rect 43994 149096 44050 149152
rect 43994 120672 44050 120728
rect 46846 285776 46902 285832
rect 50802 387640 50858 387696
rect 49606 268368 49662 268424
rect 50802 264968 50858 265024
rect 50986 387640 51042 387696
rect 50894 239400 50950 239456
rect 49606 237904 49662 237960
rect 53470 434696 53526 434752
rect 52366 214512 52422 214568
rect 56322 254088 56378 254144
rect 57610 425584 57666 425640
rect 57702 310392 57758 310448
rect 57702 283056 57758 283112
rect 56506 254088 56562 254144
rect 56414 218592 56470 218648
rect 55034 146920 55090 146976
rect 59082 391448 59138 391504
rect 60554 519424 60610 519480
rect 57794 274760 57850 274816
rect 57242 135904 57298 135960
rect 52550 77832 52606 77888
rect 56598 40568 56654 40624
rect 58346 266464 58402 266520
rect 57886 264968 57942 265024
rect 59082 271904 59138 271960
rect 60646 442992 60702 443048
rect 59174 266464 59230 266520
rect 59082 160656 59138 160712
rect 66166 603064 66222 603120
rect 61750 284824 61806 284880
rect 61106 273300 61108 273320
rect 61108 273300 61160 273320
rect 61160 273300 61162 273320
rect 61106 273264 61162 273300
rect 61934 273264 61990 273320
rect 61842 270680 61898 270736
rect 60554 261024 60610 261080
rect 61750 261024 61806 261080
rect 60462 245520 60518 245576
rect 59266 139440 59322 139496
rect 59174 94424 59230 94480
rect 61750 235864 61806 235920
rect 61842 144880 61898 144936
rect 62118 252728 62174 252784
rect 62026 221448 62082 221504
rect 61934 138080 61990 138136
rect 65798 548256 65854 548312
rect 65890 546760 65946 546816
rect 66626 579944 66682 580000
rect 66442 578584 66498 578640
rect 67178 577360 67234 577416
rect 66626 573144 66682 573200
rect 66626 571784 66682 571840
rect 66626 570152 66682 570208
rect 66810 564712 66866 564768
rect 66718 563352 66774 563408
rect 66166 561584 66222 561640
rect 66810 559272 66866 559328
rect 66166 558048 66222 558104
rect 66074 546352 66130 546408
rect 65890 534656 65946 534712
rect 65982 525000 66038 525056
rect 66718 553560 66774 553616
rect 66810 544040 66866 544096
rect 66534 543088 66590 543144
rect 66626 539960 66682 540016
rect 66074 434560 66130 434616
rect 67362 575320 67418 575376
rect 67546 576408 67602 576464
rect 67454 569880 67510 569936
rect 67454 567568 67510 567624
rect 67362 555192 67418 555248
rect 67270 552200 67326 552256
rect 79322 599392 79378 599448
rect 74262 581168 74318 581224
rect 75366 581032 75422 581088
rect 88982 601840 89038 601896
rect 79966 581168 80022 581224
rect 82726 582664 82782 582720
rect 83002 582528 83058 582584
rect 71502 580760 71558 580816
rect 80886 580760 80942 580816
rect 84198 580760 84254 580816
rect 89258 580760 89314 580816
rect 67638 566616 67694 566672
rect 67730 561992 67786 562048
rect 67638 556552 67694 556608
rect 95238 563624 95294 563680
rect 94686 558592 94742 558648
rect 67822 527720 67878 527776
rect 68926 525000 68982 525056
rect 67730 469784 67786 469840
rect 69662 448432 69718 448488
rect 66810 433356 66866 433392
rect 66810 433336 66812 433356
rect 66812 433336 66864 433356
rect 66864 433336 66866 433356
rect 66166 432540 66222 432576
rect 66166 432520 66168 432540
rect 66168 432520 66220 432540
rect 66220 432520 66222 432540
rect 64602 375264 64658 375320
rect 63314 289720 63370 289776
rect 64602 287680 64658 287736
rect 64786 287680 64842 287736
rect 64786 283328 64842 283384
rect 63406 255312 63462 255368
rect 63406 252728 63462 252784
rect 64510 135224 64566 135280
rect 66810 430344 66866 430400
rect 67362 431432 67418 431488
rect 67362 429392 67418 429448
rect 67270 429256 67326 429312
rect 67362 426264 67418 426320
rect 67362 425584 67418 425640
rect 66994 425176 67050 425232
rect 66718 424088 66774 424144
rect 66810 423272 66866 423328
rect 66810 421096 66866 421152
rect 65890 279656 65946 279712
rect 65890 268504 65946 268560
rect 66442 418920 66498 418976
rect 66442 418124 66498 418160
rect 66442 418104 66444 418124
rect 66444 418104 66496 418124
rect 66496 418104 66498 418124
rect 66902 420008 66958 420064
rect 66810 417016 66866 417072
rect 66902 415928 66958 415984
rect 66810 414840 66866 414896
rect 67362 414024 67418 414080
rect 66626 412936 66682 412992
rect 66902 411848 66958 411904
rect 66810 410760 66866 410816
rect 66442 408856 66498 408912
rect 66810 407788 66866 407824
rect 66810 407768 66812 407788
rect 66812 407768 66864 407788
rect 66864 407768 66866 407788
rect 66442 406680 66498 406736
rect 66902 404504 66958 404560
rect 66442 403688 66498 403744
rect 66442 401512 66498 401568
rect 67270 400424 67326 400480
rect 66810 399608 66866 399664
rect 67086 398520 67142 398576
rect 66810 397468 66812 397488
rect 66812 397468 66864 397488
rect 66864 397468 66866 397488
rect 66810 397432 66866 397468
rect 66258 396344 66314 396400
rect 66626 392264 66682 392320
rect 67546 428168 67602 428224
rect 67546 427372 67602 427408
rect 67546 427352 67548 427372
rect 67548 427352 67600 427372
rect 67600 427352 67602 427372
rect 67546 422184 67602 422240
rect 67546 418104 67602 418160
rect 67454 405592 67510 405648
rect 67454 398520 67510 398576
rect 67454 365608 67510 365664
rect 68926 438096 68982 438152
rect 67638 409672 67694 409728
rect 67638 402600 67694 402656
rect 67730 393372 67786 393408
rect 67730 393352 67732 393372
rect 67732 393352 67784 393372
rect 67784 393352 67786 393372
rect 67638 376488 67694 376544
rect 68558 391176 68614 391232
rect 69202 434288 69258 434344
rect 70490 436212 70546 436248
rect 70490 436192 70492 436212
rect 70492 436192 70544 436212
rect 70544 436192 70546 436212
rect 70858 436192 70914 436248
rect 69846 434696 69902 434752
rect 94318 539824 94374 539880
rect 89718 539688 89774 539744
rect 74446 452648 74502 452704
rect 72606 434832 72662 434888
rect 70674 433644 70676 433664
rect 70676 433644 70728 433664
rect 70728 433644 70730 433664
rect 70674 433608 70730 433644
rect 74078 433608 74134 433664
rect 80150 538328 80206 538384
rect 76562 442992 76618 443048
rect 75182 436192 75238 436248
rect 74814 433608 74870 433664
rect 75458 433744 75514 433800
rect 76194 433608 76250 433664
rect 77390 437552 77446 437608
rect 81346 525816 81402 525872
rect 80058 458768 80114 458824
rect 81346 457408 81402 457464
rect 84014 538056 84070 538112
rect 84290 533296 84346 533352
rect 79322 437552 79378 437608
rect 80242 436328 80298 436384
rect 80058 436192 80114 436248
rect 82082 436056 82138 436112
rect 80978 434288 81034 434344
rect 87694 536696 87750 536752
rect 88338 530712 88394 530768
rect 88982 484336 89038 484392
rect 88982 482976 89038 483032
rect 83738 434424 83794 434480
rect 84566 434288 84622 434344
rect 90362 469240 90418 469296
rect 91006 469240 91062 469296
rect 94594 538872 94650 538928
rect 94778 555464 94834 555520
rect 90362 438096 90418 438152
rect 89350 436736 89406 436792
rect 85854 434288 85910 434344
rect 91098 436056 91154 436112
rect 94778 523640 94834 523696
rect 95422 565800 95478 565856
rect 95330 558864 95386 558920
rect 95330 545672 95386 545728
rect 95238 520920 95294 520976
rect 94594 482160 94650 482216
rect 115294 604424 115350 604480
rect 98550 581168 98606 581224
rect 96802 578856 96858 578912
rect 97906 577496 97962 577552
rect 97906 576680 97962 576736
rect 96802 574776 96858 574832
rect 96894 573416 96950 573472
rect 97906 572636 97908 572656
rect 97908 572636 97960 572656
rect 97960 572636 97962 572656
rect 97906 572600 97962 572636
rect 97722 571396 97778 571432
rect 97722 571376 97724 571396
rect 97724 571376 97776 571396
rect 97776 571376 97778 571396
rect 97906 570016 97962 570072
rect 96710 569064 96766 569120
rect 97446 569064 97502 569120
rect 96802 567840 96858 567896
rect 96894 561040 96950 561096
rect 96710 556824 96766 556880
rect 96618 552064 96674 552120
rect 96434 533296 96490 533352
rect 96986 559544 97042 559600
rect 97906 556844 97962 556880
rect 97906 556824 97908 556844
rect 97908 556824 97960 556844
rect 97960 556824 97962 556844
rect 96986 554104 97042 554160
rect 96894 541728 96950 541784
rect 95330 444896 95386 444952
rect 97906 552744 97962 552800
rect 97906 552064 97962 552120
rect 97538 544312 97594 544368
rect 97538 542952 97594 543008
rect 97906 541728 97962 541784
rect 98090 562264 98146 562320
rect 101402 551928 101458 551984
rect 105542 581032 105598 581088
rect 95698 434288 95754 434344
rect 96894 436056 96950 436112
rect 98734 462304 98790 462360
rect 98642 451832 98698 451888
rect 98642 436736 98698 436792
rect 100206 434288 100262 434344
rect 107658 436192 107714 436248
rect 108946 436192 109002 436248
rect 112994 454008 113050 454064
rect 92662 434152 92718 434208
rect 90638 433880 90694 433936
rect 101218 433744 101274 433800
rect 78126 433608 78182 433664
rect 85854 433608 85910 433664
rect 87326 433608 87382 433664
rect 87970 433608 88026 433664
rect 89626 433608 89682 433664
rect 90086 433608 90142 433664
rect 91558 433608 91614 433664
rect 92938 433608 92994 433664
rect 98458 433608 98514 433664
rect 99838 433608 99894 433664
rect 100942 433608 100998 433664
rect 105174 433608 105230 433664
rect 106738 433608 106794 433664
rect 109498 433608 109554 433664
rect 111706 433608 111762 433664
rect 113270 428168 113326 428224
rect 113178 420824 113234 420880
rect 113086 407108 113142 407144
rect 113086 407088 113088 407108
rect 113088 407088 113140 407108
rect 113140 407088 113142 407108
rect 82174 390904 82230 390960
rect 85486 390904 85542 390960
rect 83186 390632 83242 390688
rect 67362 324944 67418 325000
rect 67270 282104 67326 282160
rect 67270 281288 67326 281344
rect 66810 278840 66866 278896
rect 66902 276392 66958 276448
rect 66074 272312 66130 272368
rect 65982 266600 66038 266656
rect 65890 240760 65946 240816
rect 66442 274760 66498 274816
rect 66810 273128 66866 273184
rect 66626 272312 66682 272368
rect 66810 271904 66866 271960
rect 66534 270680 66590 270736
rect 66810 269864 66866 269920
rect 66810 268232 66866 268288
rect 66810 264988 66866 265024
rect 66810 264968 66812 264988
rect 66812 264968 66864 264988
rect 66864 264968 66866 264988
rect 66626 264152 66682 264208
rect 67086 263336 67142 263392
rect 66902 262520 66958 262576
rect 66258 260888 66314 260944
rect 66810 258440 66866 258496
rect 66258 257624 66314 257680
rect 67546 281288 67602 281344
rect 67546 278024 67602 278080
rect 67454 263336 67510 263392
rect 67362 256808 67418 256864
rect 66810 255176 66866 255232
rect 66994 253544 67050 253600
rect 66810 251912 66866 251968
rect 66810 250280 66866 250336
rect 66442 248648 66498 248704
rect 66810 247832 66866 247888
rect 66718 243752 66774 243808
rect 66810 242120 66866 242176
rect 66166 162696 66222 162752
rect 64786 136992 64842 137048
rect 64694 136856 64750 136912
rect 66074 153176 66130 153232
rect 65982 121352 66038 121408
rect 66810 133592 66866 133648
rect 66810 131960 66866 132016
rect 66258 131144 66314 131200
rect 67178 129784 67234 129840
rect 66810 128152 66866 128208
rect 66166 125976 66222 126032
rect 66902 124344 66958 124400
rect 66810 123800 66866 123856
rect 66258 122984 66314 123040
rect 66350 122168 66406 122224
rect 66902 120672 66958 120728
rect 66810 120536 66866 120592
rect 66810 120028 66812 120048
rect 66812 120028 66864 120048
rect 66864 120028 66866 120048
rect 66810 119992 66866 120028
rect 66902 119176 66958 119232
rect 66810 118360 66866 118416
rect 66902 117544 66958 117600
rect 66074 117000 66130 117056
rect 66810 116184 66866 116240
rect 66810 115368 66866 115424
rect 66810 114552 66866 114608
rect 66810 113736 66866 113792
rect 65982 113192 66038 113248
rect 66810 112376 66866 112432
rect 66902 111560 66958 111616
rect 66810 110744 66866 110800
rect 66902 110200 66958 110256
rect 66810 109384 66866 109440
rect 66442 108568 66498 108624
rect 66718 107752 66774 107808
rect 66994 106956 67050 106992
rect 66994 106936 66996 106956
rect 66996 106936 67048 106956
rect 67048 106936 67050 106956
rect 66534 105596 66590 105632
rect 66534 105576 66536 105596
rect 66536 105576 66588 105596
rect 66588 105576 66590 105596
rect 66350 104796 66352 104816
rect 66352 104796 66404 104816
rect 66404 104796 66406 104816
rect 66350 104760 66406 104796
rect 67454 246200 67510 246256
rect 67454 233144 67510 233200
rect 67362 150592 67418 150648
rect 67362 106936 67418 106992
rect 67270 103944 67326 104000
rect 66534 103128 66590 103184
rect 66626 102584 66682 102640
rect 64786 83680 64842 83736
rect 63406 82728 63462 82784
rect 66810 101768 66866 101824
rect 67270 100136 67326 100192
rect 66810 99628 66812 99648
rect 66812 99628 66864 99648
rect 66864 99628 66866 99648
rect 66810 99592 66866 99628
rect 66810 98776 66866 98832
rect 66810 94968 66866 95024
rect 72422 390360 72478 390416
rect 72422 389272 72478 389328
rect 71686 383560 71742 383616
rect 70490 383424 70546 383480
rect 70398 362208 70454 362264
rect 70306 307808 70362 307864
rect 69662 291080 69718 291136
rect 69018 288496 69074 288552
rect 69846 287136 69902 287192
rect 67822 283192 67878 283248
rect 73066 386960 73122 387016
rect 73802 382880 73858 382936
rect 73158 371184 73214 371240
rect 71870 283600 71926 283656
rect 72422 283600 72478 283656
rect 70858 282920 70914 282976
rect 71594 283464 71650 283520
rect 71962 283464 72018 283520
rect 77206 390360 77262 390416
rect 77206 388728 77262 388784
rect 77482 388456 77538 388512
rect 77206 369144 77262 369200
rect 74630 288632 74686 288688
rect 73802 285776 73858 285832
rect 73250 283464 73306 283520
rect 73894 284144 73950 284200
rect 75826 283464 75882 283520
rect 78586 385056 78642 385112
rect 76654 309032 76710 309088
rect 76562 284144 76618 284200
rect 77298 306448 77354 306504
rect 78770 386824 78826 386880
rect 80058 390088 80114 390144
rect 79414 384920 79470 384976
rect 78678 284144 78734 284200
rect 79966 293120 80022 293176
rect 81300 390088 81356 390144
rect 80886 385736 80942 385792
rect 80702 378664 80758 378720
rect 80058 291080 80114 291136
rect 82726 387504 82782 387560
rect 81990 376352 82046 376408
rect 80794 311072 80850 311128
rect 82634 304136 82690 304192
rect 82082 291080 82138 291136
rect 79046 283464 79102 283520
rect 82910 346432 82966 346488
rect 92018 390768 92074 390824
rect 89718 390632 89774 390688
rect 86866 382880 86922 382936
rect 85578 382200 85634 382256
rect 84106 312432 84162 312488
rect 84014 308352 84070 308408
rect 71870 283192 71926 283248
rect 81990 283056 82046 283112
rect 83094 285776 83150 285832
rect 83462 305768 83518 305824
rect 84014 285776 84070 285832
rect 86774 313928 86830 313984
rect 84106 285640 84162 285696
rect 87970 389136 88026 389192
rect 89626 385872 89682 385928
rect 88338 373224 88394 373280
rect 86958 307672 87014 307728
rect 86866 285640 86922 285696
rect 87326 291080 87382 291136
rect 88246 306992 88302 307048
rect 89442 316648 89498 316704
rect 88430 294616 88486 294672
rect 88246 291080 88302 291136
rect 87602 290400 87658 290456
rect 87326 289856 87382 289912
rect 88614 287816 88670 287872
rect 88430 283056 88486 283112
rect 89166 285912 89222 285968
rect 81990 282920 82046 282976
rect 82634 282920 82690 282976
rect 83462 282920 83518 282976
rect 86314 282920 86370 282976
rect 89074 282920 89130 282976
rect 90454 388864 90510 388920
rect 91098 384240 91154 384296
rect 99470 390904 99526 390960
rect 106002 390904 106058 390960
rect 96802 390768 96858 390824
rect 93398 387504 93454 387560
rect 91006 311072 91062 311128
rect 90362 305632 90418 305688
rect 89718 289584 89774 289640
rect 90270 286048 90326 286104
rect 89810 283464 89866 283520
rect 95146 382336 95202 382392
rect 93766 315288 93822 315344
rect 91098 301552 91154 301608
rect 91006 286048 91062 286104
rect 92294 284144 92350 284200
rect 92386 283600 92442 283656
rect 94502 309712 94558 309768
rect 93950 284280 94006 284336
rect 94042 283464 94098 283520
rect 97078 390768 97134 390824
rect 96894 389000 96950 389056
rect 97630 389000 97686 389056
rect 97262 377440 97318 377496
rect 98918 389136 98974 389192
rect 99470 387912 99526 387968
rect 95330 312432 95386 312488
rect 95238 289992 95294 290048
rect 94686 283328 94742 283384
rect 99286 370504 99342 370560
rect 96894 283328 96950 283384
rect 90730 282920 90786 282976
rect 67822 277208 67878 277264
rect 67730 260072 67786 260128
rect 68190 258712 68246 258768
rect 67730 251096 67786 251152
rect 67822 249464 67878 249520
rect 100666 390360 100722 390416
rect 99470 316648 99526 316704
rect 100114 289856 100170 289912
rect 98918 282920 98974 282976
rect 99470 271224 99526 271280
rect 99378 258984 99434 259040
rect 98366 258712 98422 258768
rect 98090 247016 98146 247072
rect 71134 241712 71190 241768
rect 74906 241712 74962 241768
rect 76654 241712 76710 241768
rect 69294 241440 69350 241496
rect 69570 241440 69626 241496
rect 71318 241440 71374 241496
rect 71778 240080 71834 240136
rect 67730 132776 67786 132832
rect 67730 128968 67786 129024
rect 67546 97960 67602 98016
rect 67454 97144 67510 97200
rect 67546 86672 67602 86728
rect 60738 46144 60794 46200
rect 67914 143792 67970 143848
rect 67822 127608 67878 127664
rect 70398 155896 70454 155952
rect 70398 154808 70454 154864
rect 69110 143384 69166 143440
rect 69018 142976 69074 143032
rect 70214 139576 70270 139632
rect 70306 135088 70362 135144
rect 70306 134988 70308 135008
rect 70308 134988 70360 135008
rect 70360 134988 70362 135008
rect 70306 134952 70362 134988
rect 72790 239808 72846 239864
rect 73526 239944 73582 240000
rect 72882 239400 72938 239456
rect 74446 240080 74502 240136
rect 71778 233996 71780 234016
rect 71780 233996 71832 234016
rect 71832 233996 71834 234016
rect 71778 233960 71834 233996
rect 75458 240080 75514 240136
rect 76562 238856 76618 238912
rect 72422 157392 72478 157448
rect 71042 155896 71098 155952
rect 71318 138216 71374 138272
rect 73618 139304 73674 139360
rect 77666 241712 77722 241768
rect 78402 241712 78458 241768
rect 79874 241712 79930 241768
rect 77298 238584 77354 238640
rect 74722 149640 74778 149696
rect 74446 134816 74502 134872
rect 75918 176160 75974 176216
rect 75642 134680 75698 134736
rect 77666 240080 77722 240136
rect 78402 240080 78458 240136
rect 77574 236544 77630 236600
rect 80150 238448 80206 238504
rect 80150 237904 80206 237960
rect 81990 241712 82046 241768
rect 83738 241712 83794 241768
rect 85946 241712 86002 241768
rect 86590 241712 86646 241768
rect 91558 241712 91614 241768
rect 77942 164328 77998 164384
rect 79966 141344 80022 141400
rect 79598 137284 79654 137320
rect 79598 137264 79600 137284
rect 79600 137264 79652 137284
rect 79652 137264 79654 137284
rect 78770 136584 78826 136640
rect 82910 238312 82966 238368
rect 82174 176704 82230 176760
rect 84290 238584 84346 238640
rect 83554 220088 83610 220144
rect 85578 211792 85634 211848
rect 88430 240080 88486 240136
rect 83554 177248 83610 177304
rect 82082 140800 82138 140856
rect 83002 156032 83058 156088
rect 86314 172352 86370 172408
rect 86314 171128 86370 171184
rect 86130 143520 86186 143576
rect 84842 142024 84898 142080
rect 84750 139984 84806 140040
rect 86958 164464 87014 164520
rect 86866 144744 86922 144800
rect 90270 241576 90326 241632
rect 89626 239944 89682 240000
rect 90822 241576 90878 241632
rect 88246 151000 88302 151056
rect 89718 167048 89774 167104
rect 88982 149640 89038 149696
rect 89166 147736 89222 147792
rect 88430 142024 88486 142080
rect 89074 137264 89130 137320
rect 91098 240080 91154 240136
rect 91098 236000 91154 236056
rect 91926 239436 91928 239456
rect 91928 239436 91980 239456
rect 91980 239436 91982 239456
rect 91926 239400 91982 239436
rect 92386 236408 92442 236464
rect 90822 144744 90878 144800
rect 90822 140800 90878 140856
rect 91006 136856 91062 136912
rect 91098 135904 91154 135960
rect 91282 135904 91338 135960
rect 94778 237224 94834 237280
rect 94134 234096 94190 234152
rect 92478 145560 92534 145616
rect 94870 138080 94926 138136
rect 67914 125160 67970 125216
rect 67822 100952 67878 101008
rect 68558 95784 68614 95840
rect 69018 94424 69074 94480
rect 68006 93336 68062 93392
rect 67822 91976 67878 92032
rect 68374 89528 68430 89584
rect 69846 91024 69902 91080
rect 69846 85312 69902 85368
rect 69018 82048 69074 82104
rect 68006 60560 68062 60616
rect 71778 92384 71834 92440
rect 70858 86536 70914 86592
rect 70398 76472 70454 76528
rect 71778 87896 71834 87952
rect 74308 92656 74364 92712
rect 74860 92656 74916 92712
rect 73342 92384 73398 92440
rect 74446 71712 74502 71768
rect 75366 92520 75422 92576
rect 76884 92656 76940 92712
rect 76286 92248 76342 92304
rect 78954 91024 79010 91080
rect 78402 89664 78458 89720
rect 78034 89392 78090 89448
rect 77298 80008 77354 80064
rect 81438 92384 81494 92440
rect 82082 88032 82138 88088
rect 83554 92384 83610 92440
rect 83002 86808 83058 86864
rect 89626 92676 89682 92712
rect 89626 92656 89628 92676
rect 89628 92656 89680 92676
rect 89680 92656 89682 92676
rect 85670 83952 85726 84008
rect 90362 84768 90418 84824
rect 89902 75792 89958 75848
rect 95974 164464 96030 164520
rect 95974 164192 96030 164248
rect 95330 120264 95386 120320
rect 92754 92248 92810 92304
rect 94502 90364 94558 90400
rect 94502 90344 94504 90364
rect 94504 90344 94556 90364
rect 94556 90344 94558 90364
rect 91466 83816 91522 83872
rect 91098 81368 91154 81424
rect 96710 133048 96766 133104
rect 96710 132232 96766 132288
rect 96802 130872 96858 130928
rect 96710 130056 96766 130112
rect 96618 125432 96674 125488
rect 96526 103556 96582 103592
rect 96526 103536 96528 103556
rect 96528 103536 96580 103556
rect 96580 103536 96582 103556
rect 95422 89528 95478 89584
rect 96710 114008 96766 114064
rect 97354 144744 97410 144800
rect 97354 131416 97410 131472
rect 97446 127608 97502 127664
rect 97630 127064 97686 127120
rect 97262 126248 97318 126304
rect 97538 124616 97594 124672
rect 97906 124108 97908 124128
rect 97908 124108 97960 124128
rect 97960 124108 97962 124128
rect 97906 124072 97962 124108
rect 97170 123256 97226 123312
rect 97538 122440 97594 122496
rect 97722 120808 97778 120864
rect 97538 120264 97594 120320
rect 97722 119448 97778 119504
rect 97906 118652 97962 118688
rect 97906 118632 97908 118652
rect 97908 118632 97960 118652
rect 97960 118632 97962 118652
rect 97354 117000 97410 117056
rect 97906 116456 97962 116512
rect 97906 115640 97962 115696
rect 97814 114824 97870 114880
rect 97538 113464 97594 113520
rect 97906 112648 97962 112704
rect 96894 111868 96896 111888
rect 96896 111868 96948 111888
rect 96948 111868 96950 111888
rect 96894 111832 96950 111868
rect 97354 111016 97410 111072
rect 97814 109656 97870 109712
rect 96986 107208 97042 107264
rect 97906 108024 97962 108080
rect 97538 105848 97594 105904
rect 96894 105032 96950 105088
rect 97722 104216 97778 104272
rect 97906 102856 97962 102912
rect 97906 102060 97962 102096
rect 97906 102040 97908 102060
rect 97908 102040 97960 102060
rect 97960 102040 97962 102060
rect 97906 101224 97962 101280
rect 100206 283328 100262 283384
rect 100850 282648 100906 282704
rect 100758 281832 100814 281888
rect 100850 281016 100906 281072
rect 100758 279384 100814 279440
rect 100758 277752 100814 277808
rect 100022 262248 100078 262304
rect 99562 249192 99618 249248
rect 98734 223488 98790 223544
rect 98734 222264 98790 222320
rect 98090 110200 98146 110256
rect 98734 104080 98790 104136
rect 97538 100408 97594 100464
rect 97906 99592 97962 99648
rect 98642 99456 98698 99512
rect 96894 99048 96950 99104
rect 97354 98232 97410 98288
rect 97906 97416 97962 97472
rect 96894 96600 96950 96656
rect 97262 95240 97318 95296
rect 96986 94460 96988 94480
rect 96988 94460 97040 94480
rect 97040 94460 97042 94480
rect 96986 94424 97042 94460
rect 96802 84768 96858 84824
rect 97906 93608 97962 93664
rect 100666 245928 100722 245984
rect 101034 276936 101090 276992
rect 100850 276120 100906 276176
rect 100942 275304 100998 275360
rect 101034 275168 101090 275224
rect 100850 274488 100906 274544
rect 103334 382880 103390 382936
rect 101402 273672 101458 273728
rect 100850 272856 100906 272912
rect 101494 271224 101550 271280
rect 100850 270444 100852 270464
rect 100852 270444 100904 270464
rect 100904 270444 100906 270464
rect 100850 270408 100906 270444
rect 100850 267960 100906 268016
rect 101034 266328 101090 266384
rect 100850 265512 100906 265568
rect 100942 264696 100998 264752
rect 100850 263064 100906 263120
rect 101126 262248 101182 262304
rect 100850 261468 100852 261488
rect 100852 261468 100904 261488
rect 100904 261468 100906 261488
rect 100850 261432 100906 261468
rect 101034 261432 101090 261488
rect 100850 260616 100906 260672
rect 101954 259800 102010 259856
rect 101402 257352 101458 257408
rect 100942 256536 100998 256592
rect 100850 255720 100906 255776
rect 100850 254904 100906 254960
rect 100850 253272 100906 253328
rect 100850 250824 100906 250880
rect 100942 250008 100998 250064
rect 100850 248376 100906 248432
rect 100850 245112 100906 245168
rect 100850 243480 100906 243536
rect 100850 242664 100906 242720
rect 101034 244296 101090 244352
rect 100758 230424 100814 230480
rect 101494 216688 101550 216744
rect 100758 151000 100814 151056
rect 100022 93064 100078 93120
rect 100114 86536 100170 86592
rect 98642 82728 98698 82784
rect 98918 82728 98974 82784
rect 104254 390360 104310 390416
rect 103334 281424 103390 281480
rect 103334 280200 103390 280256
rect 105266 390360 105322 390416
rect 105174 388592 105230 388648
rect 106002 379344 106058 379400
rect 103518 239400 103574 239456
rect 103518 236680 103574 236736
rect 104714 272448 104770 272504
rect 104254 246744 104310 246800
rect 104162 233144 104218 233200
rect 104162 220088 104218 220144
rect 102782 151000 102838 151056
rect 102966 150456 103022 150512
rect 102782 117816 102838 117872
rect 104254 150592 104310 150648
rect 104162 90344 104218 90400
rect 103518 30912 103574 30968
rect 101034 3440 101090 3496
rect 104530 90344 104586 90400
rect 104530 89392 104586 89448
rect 107382 390904 107438 390960
rect 111982 390496 112038 390552
rect 106094 267008 106150 267064
rect 106094 266328 106150 266384
rect 108302 389816 108358 389872
rect 107750 380840 107806 380896
rect 106922 317464 106978 317520
rect 106186 238312 106242 238368
rect 106186 237360 106242 237416
rect 105082 91024 105138 91080
rect 105634 89800 105690 89856
rect 104990 83816 105046 83872
rect 105634 80008 105690 80064
rect 109682 371864 109738 371920
rect 109038 371320 109094 371376
rect 109682 371320 109738 371376
rect 108302 269184 108358 269240
rect 108302 266328 108358 266384
rect 107014 238448 107070 238504
rect 107658 234096 107714 234152
rect 110510 385736 110566 385792
rect 109774 263608 109830 263664
rect 109038 237360 109094 237416
rect 107658 92248 107714 92304
rect 108486 144880 108542 144936
rect 109038 88032 109094 88088
rect 112534 283192 112590 283248
rect 110510 236544 110566 236600
rect 111246 135904 111302 135960
rect 111154 89664 111210 89720
rect 113362 418920 113418 418976
rect 114926 429256 114982 429312
rect 115110 424940 115112 424960
rect 115112 424940 115164 424960
rect 115164 424940 115166 424960
rect 115110 424904 115166 424940
rect 114558 423000 114614 423056
rect 114650 420008 114706 420064
rect 114558 417832 114614 417888
rect 114466 406408 114522 406464
rect 113454 402328 113510 402384
rect 113270 304136 113326 304192
rect 112626 253952 112682 254008
rect 112718 232464 112774 232520
rect 114926 414840 114982 414896
rect 114834 400424 114890 400480
rect 116214 553968 116270 554024
rect 115294 516704 115350 516760
rect 115294 468424 115350 468480
rect 115754 433336 115810 433392
rect 115846 432248 115902 432304
rect 115846 428168 115902 428224
rect 115846 427080 115902 427136
rect 115754 425992 115810 426048
rect 115846 424088 115902 424144
rect 115846 423000 115902 423056
rect 115294 421912 115350 421968
rect 115846 418920 115902 418976
rect 115846 416780 115848 416800
rect 115848 416780 115900 416800
rect 115900 416780 115902 416800
rect 115846 416744 115902 416780
rect 115846 415676 115902 415712
rect 115846 415656 115848 415676
rect 115848 415656 115900 415676
rect 115900 415656 115902 415676
rect 115202 413752 115258 413808
rect 115846 412684 115902 412720
rect 115846 412664 115848 412684
rect 115848 412664 115900 412684
rect 115900 412664 115902 412684
rect 115754 411576 115810 411632
rect 115846 410488 115902 410544
rect 115846 409708 115848 409728
rect 115848 409708 115900 409728
rect 115900 409708 115902 409728
rect 115846 409672 115902 409708
rect 115846 408584 115902 408640
rect 115202 406408 115258 406464
rect 115846 405592 115902 405648
rect 115846 404504 115902 404560
rect 115846 403416 115902 403472
rect 115386 401240 115442 401296
rect 115846 399336 115902 399392
rect 115846 398284 115848 398304
rect 115848 398284 115900 398304
rect 115900 398284 115902 398304
rect 115846 398248 115902 398284
rect 115846 397160 115902 397216
rect 115754 396344 115810 396400
rect 115846 395256 115902 395312
rect 115846 394168 115902 394224
rect 115846 393080 115902 393136
rect 115846 392012 115902 392048
rect 115846 391992 115848 392012
rect 115848 391992 115900 392012
rect 115900 391992 115902 392012
rect 118698 584976 118754 585032
rect 119342 584976 119398 585032
rect 117318 460944 117374 461000
rect 118698 436192 118754 436248
rect 117410 389816 117466 389872
rect 116214 385736 116270 385792
rect 115938 300192 115994 300248
rect 114006 161472 114062 161528
rect 111890 109520 111946 109576
rect 115294 281424 115350 281480
rect 115294 267824 115350 267880
rect 115202 226888 115258 226944
rect 114742 104080 114798 104136
rect 116674 285776 116730 285832
rect 122102 582664 122158 582720
rect 122746 451832 122802 451888
rect 122746 451288 122802 451344
rect 119342 383424 119398 383480
rect 119986 377304 120042 377360
rect 117502 275168 117558 275224
rect 116858 142704 116914 142760
rect 116858 137264 116914 137320
rect 116030 83952 116086 84008
rect 120722 307808 120778 307864
rect 118790 234096 118846 234152
rect 120078 204992 120134 205048
rect 120170 140664 120226 140720
rect 120170 139984 120226 140040
rect 121550 236680 121606 236736
rect 122930 451288 122986 451344
rect 122838 387504 122894 387560
rect 123482 387504 123538 387560
rect 122930 378664 122986 378720
rect 123482 323720 123538 323776
rect 122102 306992 122158 307048
rect 122838 301552 122894 301608
rect 122102 165688 122158 165744
rect 121550 62736 121606 62792
rect 123482 233960 123538 234016
rect 124954 376624 125010 376680
rect 124862 332560 124918 332616
rect 124218 233960 124274 234016
rect 125138 235728 125194 235784
rect 129002 438912 129058 438968
rect 129002 391856 129058 391912
rect 127806 298016 127862 298072
rect 128266 298016 128322 298072
rect 127806 297336 127862 297392
rect 127714 236544 127770 236600
rect 126610 124072 126666 124128
rect 127714 120672 127770 120728
rect 129738 384920 129794 384976
rect 129002 241440 129058 241496
rect 129002 192480 129058 192536
rect 129094 127608 129150 127664
rect 130474 334736 130530 334792
rect 131854 328616 131910 328672
rect 133142 473184 133198 473240
rect 133694 473184 133750 473240
rect 133142 471960 133198 472016
rect 132498 434696 132554 434752
rect 133142 331200 133198 331256
rect 135166 458768 135222 458824
rect 134706 297336 134762 297392
rect 135902 327392 135958 327448
rect 134706 133864 134762 133920
rect 135994 324944 136050 325000
rect 137374 373224 137430 373280
rect 137282 369008 137338 369064
rect 137282 316648 137338 316704
rect 136086 149232 136142 149288
rect 139306 382200 139362 382256
rect 139306 381656 139362 381712
rect 137466 333240 137522 333296
rect 137558 284280 137614 284336
rect 137374 238584 137430 238640
rect 137374 237904 137430 237960
rect 138018 211012 138020 211032
rect 138020 211012 138072 211032
rect 138072 211012 138074 211032
rect 138018 210976 138074 211012
rect 137466 134408 137522 134464
rect 140042 311888 140098 311944
rect 138846 272448 138902 272504
rect 141422 375128 141478 375184
rect 140686 331064 140742 331120
rect 138754 160112 138810 160168
rect 138754 121624 138810 121680
rect 143446 610000 143502 610056
rect 142894 475224 142950 475280
rect 142066 306992 142122 307048
rect 141698 295296 141754 295352
rect 142066 295296 142122 295352
rect 141514 127608 141570 127664
rect 143354 475224 143410 475280
rect 143354 474816 143410 474872
rect 144734 605920 144790 605976
rect 144642 449112 144698 449168
rect 144274 377984 144330 378040
rect 144274 373224 144330 373280
rect 144182 361528 144238 361584
rect 142986 286320 143042 286376
rect 144090 331064 144146 331120
rect 143538 329840 143594 329896
rect 144090 329840 144146 329896
rect 142986 162832 143042 162888
rect 144734 377984 144790 378040
rect 144734 310392 144790 310448
rect 144734 309712 144790 309768
rect 144182 272448 144238 272504
rect 145562 311072 145618 311128
rect 144826 257896 144882 257952
rect 145654 283464 145710 283520
rect 147494 516704 147550 516760
rect 147494 390496 147550 390552
rect 147494 389272 147550 389328
rect 146942 373224 146998 373280
rect 146206 333240 146262 333296
rect 146942 309304 146998 309360
rect 145654 151816 145710 151872
rect 147126 317464 147182 317520
rect 148874 523640 148930 523696
rect 148322 381520 148378 381576
rect 148414 284960 148470 285016
rect 150162 455504 150218 455560
rect 149058 397976 149114 398032
rect 149702 376352 149758 376408
rect 149702 333376 149758 333432
rect 148874 316004 148876 316024
rect 148876 316004 148928 316024
rect 148928 316004 148930 316024
rect 148874 315968 148930 316004
rect 148690 313248 148746 313304
rect 148598 285912 148654 285968
rect 148598 243480 148654 243536
rect 148506 228248 148562 228304
rect 148598 153720 148654 153776
rect 150346 397976 150402 398032
rect 151082 535336 151138 535392
rect 151634 450064 151690 450120
rect 151266 347792 151322 347848
rect 150438 113736 150494 113792
rect 152462 533296 152518 533352
rect 151174 241576 151230 241632
rect 151174 220088 151230 220144
rect 151174 144880 151230 144936
rect 151174 98232 151230 98288
rect 151174 86672 151230 86728
rect 152738 321544 152794 321600
rect 152554 318144 152610 318200
rect 152554 317464 152610 317520
rect 152646 301144 152702 301200
rect 173806 611360 173862 611416
rect 160742 608640 160798 608696
rect 155866 607280 155922 607336
rect 153934 570560 153990 570616
rect 153934 458088 153990 458144
rect 153842 456048 153898 456104
rect 153106 420824 153162 420880
rect 152922 318144 152978 318200
rect 153198 335416 153254 335472
rect 153290 326304 153346 326360
rect 153106 289720 153162 289776
rect 153106 289040 153162 289096
rect 154302 384376 154358 384432
rect 154394 368328 154450 368384
rect 155222 398928 155278 398984
rect 155682 387640 155738 387696
rect 155682 386960 155738 387016
rect 154486 343576 154542 343632
rect 154486 342896 154542 342952
rect 154026 338680 154082 338736
rect 154486 330520 154542 330576
rect 154118 319368 154174 319424
rect 155222 314744 155278 314800
rect 154486 162696 154542 162752
rect 154486 158752 154542 158808
rect 153934 154672 153990 154728
rect 153934 145560 153990 145616
rect 155406 261432 155462 261488
rect 156602 366968 156658 367024
rect 157246 366968 157302 367024
rect 156602 306992 156658 307048
rect 155866 136448 155922 136504
rect 155866 135224 155922 135280
rect 156694 240760 156750 240816
rect 156694 136448 156750 136504
rect 158626 564984 158682 565040
rect 158442 331744 158498 331800
rect 158810 451868 158812 451888
rect 158812 451868 158864 451888
rect 158864 451868 158866 451888
rect 158810 451832 158866 451868
rect 165526 600480 165582 600536
rect 159914 451832 159970 451888
rect 159914 442992 159970 443048
rect 159914 316648 159970 316704
rect 159362 312024 159418 312080
rect 158626 266328 158682 266384
rect 158718 235864 158774 235920
rect 158718 234640 158774 234696
rect 158074 160656 158130 160712
rect 161294 471144 161350 471200
rect 161202 391176 161258 391232
rect 160374 390360 160430 390416
rect 160374 389136 160430 389192
rect 160190 306856 160246 306912
rect 158718 143384 158774 143440
rect 159362 143384 159418 143440
rect 158718 142704 158774 142760
rect 159638 234640 159694 234696
rect 159638 204176 159694 204232
rect 159546 153176 159602 153232
rect 159362 139440 159418 139496
rect 161386 389136 161442 389192
rect 163594 442992 163650 443048
rect 161570 390360 161626 390416
rect 161478 376488 161534 376544
rect 162122 376488 162178 376544
rect 160742 143248 160798 143304
rect 159638 139440 159694 139496
rect 159362 111832 159418 111888
rect 161294 326304 161350 326360
rect 163870 384920 163926 384976
rect 163870 384240 163926 384296
rect 162122 327256 162178 327312
rect 162122 323720 162178 323776
rect 162122 317464 162178 317520
rect 162122 253816 162178 253872
rect 160926 146920 160982 146976
rect 162674 244296 162730 244352
rect 164146 457408 164202 457464
rect 163962 290400 164018 290456
rect 162858 266328 162914 266384
rect 163502 218592 163558 218648
rect 164882 384920 164938 384976
rect 165526 336096 165582 336152
rect 166446 460128 166502 460184
rect 166446 453192 166502 453248
rect 166354 414568 166410 414624
rect 165618 284824 165674 284880
rect 165618 284280 165674 284336
rect 166262 330520 166318 330576
rect 166262 302776 166318 302832
rect 168194 529080 168250 529136
rect 167642 483656 167698 483712
rect 166538 428440 166594 428496
rect 166998 369824 167054 369880
rect 165066 238584 165122 238640
rect 166446 284280 166502 284336
rect 166906 231784 166962 231840
rect 167734 386280 167790 386336
rect 167734 371184 167790 371240
rect 167734 369824 167790 369880
rect 168194 369688 168250 369744
rect 167642 318008 167698 318064
rect 167090 285640 167146 285696
rect 169114 579672 169170 579728
rect 169206 513324 169262 513360
rect 169206 513304 169208 513324
rect 169208 513304 169260 513324
rect 169260 513304 169262 513324
rect 169114 489096 169170 489152
rect 169022 365608 169078 365664
rect 167642 260480 167698 260536
rect 166446 136992 166502 137048
rect 168286 235864 168342 235920
rect 167734 234640 167790 234696
rect 168286 234640 168342 234696
rect 172334 589872 172390 589928
rect 170402 502968 170458 503024
rect 170494 471144 170550 471200
rect 169666 465704 169722 465760
rect 169114 311344 169170 311400
rect 170862 471144 170918 471200
rect 170770 439456 170826 439512
rect 170954 465704 171010 465760
rect 170954 390768 171010 390824
rect 170494 386144 170550 386200
rect 170494 366832 170550 366888
rect 169298 260480 169354 260536
rect 171782 462848 171838 462904
rect 171046 383560 171102 383616
rect 171874 386144 171930 386200
rect 171782 369688 171838 369744
rect 173162 581032 173218 581088
rect 172334 457544 172390 457600
rect 173162 553968 173218 554024
rect 173622 440816 173678 440872
rect 173162 397976 173218 398032
rect 172426 393896 172482 393952
rect 172242 386144 172298 386200
rect 173622 387640 173678 387696
rect 173622 381656 173678 381712
rect 173162 379208 173218 379264
rect 170402 250416 170458 250472
rect 169758 237224 169814 237280
rect 169114 235728 169170 235784
rect 169666 235728 169722 235784
rect 169666 136584 169722 136640
rect 171138 257896 171194 257952
rect 171782 341400 171838 341456
rect 172242 330384 172298 330440
rect 171230 239808 171286 239864
rect 171782 224848 171838 224904
rect 172334 210976 172390 211032
rect 173714 322904 173770 322960
rect 173254 270408 173310 270464
rect 173162 244296 173218 244352
rect 172518 239808 172574 239864
rect 172518 239400 172574 239456
rect 172426 176568 172482 176624
rect 172334 92792 172390 92848
rect 175094 482160 175150 482216
rect 175002 450200 175058 450256
rect 173806 311208 173862 311264
rect 173898 288360 173954 288416
rect 173898 287680 173954 287736
rect 173714 244568 173770 244624
rect 173714 244296 173770 244352
rect 175554 343576 175610 343632
rect 178774 547032 178830 547088
rect 177302 390904 177358 390960
rect 175186 316104 175242 316160
rect 174634 288360 174690 288416
rect 175186 302504 175242 302560
rect 177670 382336 177726 382392
rect 177302 322904 177358 322960
rect 175186 256012 175242 256048
rect 175186 255992 175188 256012
rect 175188 255992 175240 256012
rect 175240 255992 175242 256012
rect 174542 138624 174598 138680
rect 174542 138080 174598 138136
rect 176658 312024 176714 312080
rect 176658 311344 176714 311400
rect 176658 309712 176714 309768
rect 176106 306720 176162 306776
rect 176106 298016 176162 298072
rect 177762 342896 177818 342952
rect 177670 312024 177726 312080
rect 177486 310528 177542 310584
rect 176658 260072 176714 260128
rect 176198 249056 176254 249112
rect 175922 156168 175978 156224
rect 176014 146240 176070 146296
rect 176566 146240 176622 146296
rect 176014 145016 176070 145072
rect 176014 141344 176070 141400
rect 176014 138080 176070 138136
rect 178038 398792 178094 398848
rect 180614 539688 180670 539744
rect 179510 538328 179566 538384
rect 178038 390904 178094 390960
rect 178682 269728 178738 269784
rect 178682 257216 178738 257272
rect 177762 253952 177818 254008
rect 177394 92112 177450 92168
rect 176658 76472 176714 76528
rect 176566 65456 176622 65512
rect 179142 387504 179198 387560
rect 179418 391992 179474 392048
rect 180614 485832 180670 485888
rect 180522 435920 180578 435976
rect 180522 417424 180578 417480
rect 178774 239944 178830 240000
rect 179234 237904 179290 237960
rect 178866 96600 178922 96656
rect 179234 96600 179290 96656
rect 178866 92384 178922 92440
rect 180154 384240 180210 384296
rect 181442 464480 181498 464536
rect 180706 394032 180762 394088
rect 180798 393352 180854 393408
rect 180706 391992 180762 392048
rect 180246 380704 180302 380760
rect 182178 448432 182234 448488
rect 183006 485016 183062 485072
rect 182914 469240 182970 469296
rect 183006 467744 183062 467800
rect 182914 454824 182970 454880
rect 182822 435920 182878 435976
rect 182822 389272 182878 389328
rect 180246 289040 180302 289096
rect 180154 253952 180210 254008
rect 181442 254088 181498 254144
rect 180246 229744 180302 229800
rect 180062 86808 180118 86864
rect 181994 320864 182050 320920
rect 183282 390632 183338 390688
rect 184202 597760 184258 597816
rect 184202 468560 184258 468616
rect 184662 458768 184718 458824
rect 183374 351056 183430 351112
rect 182822 306584 182878 306640
rect 182914 291896 182970 291952
rect 182914 283464 182970 283520
rect 182086 247424 182142 247480
rect 181534 241032 181590 241088
rect 181534 231104 181590 231160
rect 181534 204856 181590 204912
rect 181442 77832 181498 77888
rect 182546 236000 182602 236056
rect 185582 601976 185638 602032
rect 186962 600616 187018 600672
rect 186226 578312 186282 578368
rect 184846 449132 184902 449168
rect 184846 449112 184848 449132
rect 184848 449112 184900 449132
rect 184900 449112 184902 449132
rect 187330 555192 187386 555248
rect 185674 480800 185730 480856
rect 186226 475360 186282 475416
rect 186134 449384 186190 449440
rect 184938 390632 184994 390688
rect 184938 389816 184994 389872
rect 184294 373904 184350 373960
rect 184846 345616 184902 345672
rect 182914 237904 182970 237960
rect 182914 143656 182970 143712
rect 185674 309440 185730 309496
rect 186042 290400 186098 290456
rect 184846 240760 184902 240816
rect 183558 60560 183614 60616
rect 147126 3440 147182 3496
rect 184386 143520 184442 143576
rect 184754 120692 184810 120728
rect 184754 120672 184756 120692
rect 184756 120672 184808 120692
rect 184808 120672 184810 120692
rect 184846 92656 184902 92712
rect 185582 257236 185638 257272
rect 185582 257216 185584 257236
rect 185584 257216 185636 257236
rect 185636 257216 185638 257236
rect 187606 599528 187662 599584
rect 187146 468560 187202 468616
rect 188342 584976 188398 585032
rect 188434 537920 188490 537976
rect 188342 536016 188398 536072
rect 188342 511264 188398 511320
rect 187606 458496 187662 458552
rect 187790 458224 187846 458280
rect 188342 460264 188398 460320
rect 187606 446392 187662 446448
rect 186318 390904 186374 390960
rect 189722 612720 189778 612776
rect 187054 386960 187110 387016
rect 186962 383016 187018 383072
rect 187606 390496 187662 390552
rect 187698 386144 187754 386200
rect 188526 394032 188582 394088
rect 204350 611360 204406 611416
rect 202878 610000 202934 610056
rect 198738 608640 198794 608696
rect 191654 607824 191710 607880
rect 191194 603608 191250 603664
rect 191102 598984 191158 599040
rect 190642 596264 190698 596320
rect 190642 595176 190698 595232
rect 191010 591232 191066 591288
rect 190458 586508 190460 586528
rect 190460 586508 190512 586528
rect 190512 586508 190514 586528
rect 190458 586472 190514 586508
rect 196714 604696 196770 604752
rect 191746 598848 191802 598904
rect 191654 596808 191710 596864
rect 191746 594632 191802 594688
rect 191654 593408 191710 593464
rect 191286 589328 191342 589384
rect 191194 586200 191250 586256
rect 191102 578312 191158 578368
rect 191562 578312 191618 578368
rect 191010 576136 191066 576192
rect 191194 575592 191250 575648
rect 191286 574504 191342 574560
rect 191010 573280 191066 573336
rect 191562 572756 191618 572792
rect 191562 572736 191564 572756
rect 191564 572736 191616 572756
rect 191616 572736 191618 572756
rect 191286 572192 191342 572248
rect 191562 570832 191618 570888
rect 190918 570560 190974 570616
rect 190366 568656 190422 568712
rect 190458 567568 190514 567624
rect 190458 564984 190514 565040
rect 191102 564848 191158 564904
rect 190826 564712 190882 564768
rect 191010 563660 191012 563680
rect 191012 563660 191064 563680
rect 191064 563660 191066 563680
rect 191010 563624 191066 563660
rect 191194 560904 191250 560960
rect 191102 560632 191158 560688
rect 190918 558184 190974 558240
rect 191746 592320 191802 592376
rect 194690 600344 194746 600400
rect 192758 599256 192814 599312
rect 198554 600480 198610 600536
rect 197358 600344 197414 600400
rect 193310 597760 193366 597816
rect 197174 598984 197230 599040
rect 199842 604560 199898 604616
rect 201682 600344 201738 600400
rect 208674 603200 208730 603256
rect 211618 601976 211674 602032
rect 211618 601704 211674 601760
rect 209962 600480 210018 600536
rect 212538 599256 212594 599312
rect 213366 599120 213422 599176
rect 215298 600344 215354 600400
rect 216402 600344 216458 600400
rect 218242 609184 218298 609240
rect 219530 600752 219586 600808
rect 218242 599528 218298 599584
rect 221370 600752 221426 600808
rect 222198 612720 222254 612776
rect 222842 612720 222898 612776
rect 222290 600616 222346 600672
rect 222658 600616 222714 600672
rect 202602 598984 202658 599040
rect 207110 598984 207166 599040
rect 210422 598984 210478 599040
rect 214010 598984 214066 599040
rect 216678 598984 216734 599040
rect 218702 598984 218758 599040
rect 220910 598984 220966 599040
rect 224222 599120 224278 599176
rect 229650 601840 229706 601896
rect 228638 599120 228694 599176
rect 231490 600344 231546 600400
rect 234066 607280 234122 607336
rect 239218 606056 239274 606112
rect 238482 604424 238538 604480
rect 237562 600480 237618 600536
rect 236642 600344 236698 600400
rect 245474 605920 245530 605976
rect 243634 600616 243690 600672
rect 244186 600480 244242 600536
rect 248786 600480 248842 600536
rect 248418 599392 248474 599448
rect 250074 600344 250130 600400
rect 249338 599256 249394 599312
rect 253386 600480 253442 600536
rect 224038 598984 224094 599040
rect 226062 598984 226118 599040
rect 226798 598984 226854 599040
rect 230018 598984 230074 599040
rect 232410 598984 232466 599040
rect 233238 598984 233294 599040
rect 234710 598984 234766 599040
rect 236826 598984 236882 599040
rect 240690 598984 240746 599040
rect 247774 598984 247830 599040
rect 250902 598984 250958 599040
rect 252834 598984 252890 599040
rect 193494 598440 193550 598496
rect 253478 600344 253534 600400
rect 193402 592728 193458 592784
rect 253386 592048 253442 592104
rect 253570 599256 253626 599312
rect 253570 598984 253626 599040
rect 253938 587356 253994 587412
rect 191746 585148 191748 585168
rect 191748 585148 191800 585168
rect 191800 585148 191802 585168
rect 191746 585112 191802 585148
rect 191746 583888 191802 583944
rect 191746 582664 191802 582720
rect 191746 581576 191802 581632
rect 191746 578856 191802 578912
rect 191746 578040 191802 578096
rect 191746 567196 191748 567216
rect 191748 567196 191800 567216
rect 191800 567196 191802 567216
rect 191746 567160 191802 567196
rect 191746 561992 191802 562048
rect 191746 557776 191802 557832
rect 190826 554804 190882 554840
rect 190826 554784 190828 554804
rect 190828 554784 190880 554804
rect 190880 554784 190882 554804
rect 190918 553832 190974 553888
rect 191378 550704 191434 550760
rect 191746 556416 191802 556472
rect 191746 552084 191802 552120
rect 191746 552064 191748 552084
rect 191748 552064 191800 552084
rect 191800 552064 191802 552084
rect 191562 549752 191618 549808
rect 191746 549344 191802 549400
rect 191562 547984 191618 548040
rect 191286 547032 191342 547088
rect 191562 546524 191564 546544
rect 191564 546524 191616 546544
rect 191616 546524 191618 546544
rect 191562 546488 191618 546524
rect 191194 545400 191250 545456
rect 191102 544176 191158 544232
rect 190642 544040 190698 544096
rect 191562 542544 191618 542600
rect 190826 541456 190882 541512
rect 191470 540232 191526 540288
rect 191562 540096 191618 540152
rect 189722 469240 189778 469296
rect 191654 458768 191710 458824
rect 190366 456864 190422 456920
rect 188986 385600 189042 385656
rect 188986 378120 189042 378176
rect 190182 387368 190238 387424
rect 188342 375264 188398 375320
rect 187054 307944 187110 308000
rect 186410 305088 186466 305144
rect 186226 302504 186282 302560
rect 186410 297336 186466 297392
rect 186318 250416 186374 250472
rect 187514 304988 187516 305008
rect 187516 304988 187568 305008
rect 187568 304988 187570 305008
rect 187514 304952 187570 304988
rect 188434 373224 188490 373280
rect 188434 362888 188490 362944
rect 190274 384376 190330 384432
rect 189722 376488 189778 376544
rect 190182 376488 190238 376544
rect 187698 309168 187754 309224
rect 188066 305632 188122 305688
rect 187790 305224 187846 305280
rect 187054 286320 187110 286376
rect 186226 242392 186282 242448
rect 186318 242120 186374 242176
rect 185582 221448 185638 221504
rect 187054 241440 187110 241496
rect 187698 245792 187754 245848
rect 187146 234504 187202 234560
rect 189078 270408 189134 270464
rect 189078 269184 189134 269240
rect 189078 253816 189134 253872
rect 189814 351192 189870 351248
rect 191470 456048 191526 456104
rect 191562 449132 191618 449168
rect 191562 449112 191564 449132
rect 191564 449112 191616 449132
rect 191616 449112 191618 449132
rect 191562 447788 191564 447808
rect 191564 447788 191616 447808
rect 191616 447788 191618 447808
rect 191562 447752 191618 447788
rect 191010 446392 191066 446448
rect 191010 445032 191066 445088
rect 191562 442040 191618 442096
rect 191562 440680 191618 440736
rect 191654 437960 191710 438016
rect 191654 436600 191710 436656
rect 191654 435240 191710 435296
rect 191654 433608 191710 433664
rect 191654 432248 191710 432304
rect 191746 430888 191802 430944
rect 191010 429528 191066 429584
rect 190826 428168 190882 428224
rect 191746 426808 191802 426864
rect 191746 425448 191802 425504
rect 191010 423816 191066 423872
rect 191746 422456 191802 422512
rect 191746 417016 191802 417072
rect 191654 415384 191710 415440
rect 191194 414044 191250 414080
rect 191194 414024 191196 414044
rect 191196 414024 191248 414044
rect 191248 414024 191250 414044
rect 191102 412664 191158 412720
rect 191010 406952 191066 407008
rect 191010 402872 191066 402928
rect 191010 400152 191066 400208
rect 190826 398520 190882 398576
rect 191746 411304 191802 411360
rect 191746 409944 191802 410000
rect 191746 405628 191748 405648
rect 191748 405628 191800 405648
rect 191800 405628 191802 405648
rect 191746 405592 191802 405628
rect 191746 404268 191748 404288
rect 191748 404268 191800 404288
rect 191800 404268 191802 404288
rect 191746 404232 191802 404268
rect 191746 401548 191748 401568
rect 191748 401548 191800 401568
rect 191800 401548 191802 401568
rect 191746 401512 191802 401548
rect 191194 397160 191250 397216
rect 191102 387368 191158 387424
rect 191746 395800 191802 395856
rect 190458 370504 190514 370560
rect 190550 338680 190606 338736
rect 191746 338716 191748 338736
rect 191748 338716 191800 338736
rect 191800 338716 191802 338736
rect 191746 338680 191802 338716
rect 191746 335960 191802 336016
rect 190458 334736 190514 334792
rect 191562 330384 191618 330440
rect 189078 252592 189134 252648
rect 188986 245792 189042 245848
rect 189078 245656 189134 245712
rect 188894 234368 188950 234424
rect 188434 233960 188490 234016
rect 187514 154536 187570 154592
rect 186962 146512 187018 146568
rect 186962 135904 187018 135960
rect 187054 106664 187110 106720
rect 185122 93064 185178 93120
rect 185582 78648 185638 78704
rect 186226 78648 186282 78704
rect 187054 84088 187110 84144
rect 184294 60560 184350 60616
rect 188434 154808 188490 154864
rect 188342 144744 188398 144800
rect 188526 146376 188582 146432
rect 188342 143792 188398 143848
rect 189722 242936 189778 242992
rect 189998 299512 190054 299568
rect 189906 295432 189962 295488
rect 191470 300872 191526 300928
rect 191470 298696 191526 298752
rect 191470 297608 191526 297664
rect 191470 294344 191526 294400
rect 191470 293256 191526 293312
rect 191470 292168 191526 292224
rect 191470 291080 191526 291136
rect 190826 290012 190882 290048
rect 190826 289992 190828 290012
rect 190828 289992 190880 290012
rect 190880 289992 190882 290012
rect 191470 288904 191526 288960
rect 191470 287816 191526 287872
rect 191378 286728 191434 286784
rect 191470 285640 191526 285696
rect 191470 284552 191526 284608
rect 191470 282376 191526 282432
rect 191470 281288 191526 281344
rect 191470 280236 191472 280256
rect 191472 280236 191524 280256
rect 191524 280236 191526 280256
rect 191470 280200 191526 280236
rect 191470 279112 191526 279168
rect 191470 278024 191526 278080
rect 190642 276936 190698 276992
rect 191654 322088 191710 322144
rect 191562 275848 191618 275904
rect 190826 273672 190882 273728
rect 191562 272584 191618 272640
rect 191562 271496 191618 271552
rect 191470 270408 191526 270464
rect 191562 269356 191564 269376
rect 191564 269356 191616 269376
rect 191616 269356 191618 269376
rect 191562 269320 191618 269356
rect 191470 269184 191526 269240
rect 191562 268232 191618 268288
rect 190642 264968 190698 265024
rect 191378 260616 191434 260672
rect 190458 258032 190514 258088
rect 190642 257352 190698 257408
rect 191010 255212 191012 255232
rect 191012 255212 191064 255232
rect 191064 255212 191066 255232
rect 191010 255176 191066 255212
rect 191010 251932 191066 251968
rect 191010 251912 191012 251932
rect 191012 251912 191064 251932
rect 191064 251912 191066 251932
rect 191010 249736 191066 249792
rect 189906 239808 189962 239864
rect 189814 215872 189870 215928
rect 191654 266056 191710 266112
rect 191654 262792 191710 262848
rect 191654 261704 191710 261760
rect 191654 259528 191710 259584
rect 191654 256264 191710 256320
rect 191654 250824 191710 250880
rect 191562 248512 191618 248568
rect 193126 553084 193182 553140
rect 194138 535472 194194 535528
rect 195426 536016 195482 536072
rect 194690 531936 194746 531992
rect 192666 450336 192722 450392
rect 192758 448568 192814 448624
rect 192666 447344 192722 447400
rect 193126 461624 193182 461680
rect 193034 443672 193090 443728
rect 192390 419736 192446 419792
rect 193402 454824 193458 454880
rect 193310 452512 193366 452568
rect 193218 449384 193274 449440
rect 197450 535472 197506 535528
rect 195426 498752 195482 498808
rect 195334 491816 195390 491872
rect 195242 478080 195298 478136
rect 195334 476720 195390 476776
rect 199382 536560 199438 536616
rect 199382 535336 199438 535392
rect 198738 529080 198794 529136
rect 196622 468560 196678 468616
rect 197450 452512 197506 452568
rect 198002 490592 198058 490648
rect 197910 454008 197966 454064
rect 197542 450336 197598 450392
rect 202970 538056 203026 538112
rect 202970 536832 203026 536888
rect 203522 536832 203578 536888
rect 204442 530576 204498 530632
rect 205086 530576 205142 530632
rect 203522 512624 203578 512680
rect 202142 509768 202198 509824
rect 201498 462304 201554 462360
rect 201406 458904 201462 458960
rect 200210 456184 200266 456240
rect 198830 453192 198886 453248
rect 200854 452648 200910 452704
rect 201406 452648 201462 452704
rect 203614 489232 203670 489288
rect 202878 483656 202934 483712
rect 202786 465840 202842 465896
rect 202786 462304 202842 462360
rect 202142 454688 202198 454744
rect 203614 467200 203670 467256
rect 204902 461488 204958 461544
rect 202970 457544 203026 457600
rect 202970 454008 203026 454064
rect 202878 450472 202934 450528
rect 204074 450472 204130 450528
rect 207386 538192 207442 538248
rect 208122 535472 208178 535528
rect 206374 471144 206430 471200
rect 206466 457408 206522 457464
rect 212446 536424 212502 536480
rect 209042 489096 209098 489152
rect 209042 482976 209098 483032
rect 210238 492768 210294 492824
rect 209042 471144 209098 471200
rect 209778 470600 209834 470656
rect 209870 464616 209926 464672
rect 208398 460264 208454 460320
rect 207294 450200 207350 450256
rect 207570 450200 207626 450256
rect 212630 533296 212686 533352
rect 213274 533296 213330 533352
rect 213274 523640 213330 523696
rect 215390 536696 215446 536752
rect 214562 464480 214618 464536
rect 213918 464344 213974 464400
rect 213918 463664 213974 463720
rect 212630 454688 212686 454744
rect 218978 533296 219034 533352
rect 219530 530576 219586 530632
rect 220082 533296 220138 533352
rect 215390 461624 215446 461680
rect 215390 460264 215446 460320
rect 215390 455504 215446 455560
rect 218702 485016 218758 485072
rect 218702 482160 218758 482216
rect 223578 538192 223634 538248
rect 222842 535472 222898 535528
rect 219438 456864 219494 456920
rect 219806 456864 219862 456920
rect 222934 533976 222990 534032
rect 224682 538192 224738 538248
rect 223946 533296 224002 533352
rect 226522 535472 226578 535528
rect 223486 456864 223542 456920
rect 222198 454688 222254 454744
rect 222106 454008 222162 454064
rect 222106 453192 222162 453248
rect 223670 457408 223726 457464
rect 223670 456864 223726 456920
rect 227718 490456 227774 490512
rect 229650 533976 229706 534032
rect 228454 493448 228510 493504
rect 231122 522280 231178 522336
rect 228362 469784 228418 469840
rect 227810 464616 227866 464672
rect 205638 450064 205694 450120
rect 231214 491136 231270 491192
rect 232502 533296 232558 533352
rect 231950 480800 232006 480856
rect 231858 479440 231914 479496
rect 231306 474816 231362 474872
rect 231214 467064 231270 467120
rect 231122 459584 231178 459640
rect 230570 455912 230626 455968
rect 232134 458360 232190 458416
rect 231306 455912 231362 455968
rect 231306 455504 231362 455560
rect 235354 533296 235410 533352
rect 234618 500112 234674 500168
rect 235906 496032 235962 496088
rect 232502 453872 232558 453928
rect 233514 453872 233570 453928
rect 233514 451424 233570 451480
rect 235998 462848 236054 462904
rect 234894 454008 234950 454064
rect 235906 454008 235962 454064
rect 240782 481480 240838 481536
rect 240782 460264 240838 460320
rect 239402 453872 239458 453928
rect 239218 451832 239274 451888
rect 239218 451288 239274 451344
rect 243542 538736 243598 538792
rect 243634 535472 243690 535528
rect 244278 518064 244334 518120
rect 241426 456864 241482 456920
rect 242162 452784 242218 452840
rect 244278 462848 244334 462904
rect 247130 485016 247186 485072
rect 244922 460128 244978 460184
rect 244922 452648 244978 452704
rect 245934 450200 245990 450256
rect 228822 450064 228878 450120
rect 204166 449928 204222 449984
rect 250074 533296 250130 533352
rect 249798 527040 249854 527096
rect 250442 485832 250498 485888
rect 249062 456048 249118 456104
rect 253202 536016 253258 536072
rect 251362 492632 251418 492688
rect 251086 466520 251142 466576
rect 251086 465840 251142 465896
rect 250442 452104 250498 452160
rect 253386 556144 253442 556200
rect 255318 603064 255374 603120
rect 255962 598848 256018 598904
rect 255410 597644 255466 597680
rect 255410 597624 255412 597644
rect 255412 597624 255464 597644
rect 255464 597624 255466 597644
rect 255410 596536 255466 596592
rect 255318 594224 255374 594280
rect 255410 590960 255466 591016
rect 255410 589872 255466 589928
rect 255410 588104 255466 588160
rect 255410 585112 255466 585168
rect 255318 584160 255374 584216
rect 254030 582256 254086 582312
rect 254030 577496 254086 577552
rect 253938 538736 253994 538792
rect 254122 547848 254178 547904
rect 254214 542408 254270 542464
rect 253938 507864 253994 507920
rect 253386 481480 253442 481536
rect 251914 451424 251970 451480
rect 246118 449656 246174 449712
rect 247130 449656 247186 449712
rect 253938 472096 253994 472152
rect 253938 471144 253994 471200
rect 253570 448024 253626 448080
rect 193126 419736 193182 419792
rect 253570 413616 253626 413672
rect 192574 413208 192630 413264
rect 192482 408584 192538 408640
rect 192666 391040 192722 391096
rect 193126 390904 193182 390960
rect 193126 389408 193182 389464
rect 193402 391040 193458 391096
rect 194138 389816 194194 389872
rect 198186 387640 198242 387696
rect 201130 386280 201186 386336
rect 200210 386008 200266 386064
rect 198830 384376 198886 384432
rect 198738 383560 198794 383616
rect 198738 382880 198794 382936
rect 195978 362208 196034 362264
rect 195242 357992 195298 358048
rect 193310 320864 193366 320920
rect 192022 295976 192078 296032
rect 192022 295296 192078 295352
rect 196622 341400 196678 341456
rect 195978 316648 196034 316704
rect 195426 316104 195482 316160
rect 195334 315288 195390 315344
rect 192942 301824 192998 301880
rect 193770 301688 193826 301744
rect 193494 300736 193550 300792
rect 193494 300056 193550 300112
rect 193678 300056 193734 300112
rect 193126 298832 193182 298888
rect 192942 296928 192998 296984
rect 193678 295160 193734 295216
rect 195978 309304 196034 309360
rect 195334 301824 195390 301880
rect 195058 301688 195114 301744
rect 195978 300872 196034 300928
rect 197358 320728 197414 320784
rect 204810 389136 204866 389192
rect 204810 388728 204866 388784
rect 200762 338680 200818 338736
rect 201682 336232 201738 336288
rect 201498 331744 201554 331800
rect 200210 313248 200266 313304
rect 200762 313248 200818 313304
rect 198738 305632 198794 305688
rect 198738 304272 198794 304328
rect 201682 329160 201738 329216
rect 202050 323584 202106 323640
rect 204258 326304 204314 326360
rect 203062 318824 203118 318880
rect 208398 373224 208454 373280
rect 206374 356632 206430 356688
rect 204718 319368 204774 319424
rect 204902 319368 204958 319424
rect 206282 349696 206338 349752
rect 205638 328344 205694 328400
rect 205638 327392 205694 327448
rect 204994 315288 205050 315344
rect 205822 305088 205878 305144
rect 207294 333376 207350 333432
rect 207110 329840 207166 329896
rect 206374 328344 206430 328400
rect 206282 305088 206338 305144
rect 208398 331200 208454 331256
rect 208214 302504 208270 302560
rect 212538 389408 212594 389464
rect 213182 385600 213238 385656
rect 209778 369008 209834 369064
rect 212630 378664 212686 378720
rect 211802 359352 211858 359408
rect 209042 323584 209098 323640
rect 212538 333240 212594 333296
rect 208490 321544 208546 321600
rect 209134 321544 209190 321600
rect 208582 318144 208638 318200
rect 208582 313928 208638 313984
rect 211342 312024 211398 312080
rect 211250 311072 211306 311128
rect 213458 384240 213514 384296
rect 214562 353912 214618 353968
rect 214378 345752 214434 345808
rect 214378 341536 214434 341592
rect 213918 334736 213974 334792
rect 213090 314744 213146 314800
rect 213182 313384 213238 313440
rect 213826 306720 213882 306776
rect 221554 388864 221610 388920
rect 220082 386144 220138 386200
rect 218794 384240 218850 384296
rect 218334 381656 218390 381712
rect 217414 355272 217470 355328
rect 217322 344256 217378 344312
rect 214010 318688 214066 318744
rect 214562 318688 214618 318744
rect 214010 317464 214066 317520
rect 216678 329704 216734 329760
rect 216678 328616 216734 328672
rect 217138 305224 217194 305280
rect 217414 329704 217470 329760
rect 219438 334600 219494 334656
rect 219346 329024 219402 329080
rect 217322 305224 217378 305280
rect 219530 329160 219586 329216
rect 220726 377848 220782 377904
rect 224958 386280 225014 386336
rect 225786 386280 225842 386336
rect 222934 364928 222990 364984
rect 224222 343032 224278 343088
rect 222106 334600 222162 334656
rect 221002 327120 221058 327176
rect 222106 327120 222162 327176
rect 220082 315288 220138 315344
rect 220818 302232 220874 302288
rect 222290 328480 222346 328536
rect 223578 326984 223634 327040
rect 224222 326984 224278 327040
rect 223578 325760 223634 325816
rect 223854 304272 223910 304328
rect 223762 301144 223818 301200
rect 224958 385600 225014 385656
rect 225602 363568 225658 363624
rect 226982 351736 227038 351792
rect 225602 342896 225658 342952
rect 226982 339496 227038 339552
rect 224958 337320 225014 337376
rect 225142 337320 225198 337376
rect 225142 335416 225198 335472
rect 225878 311208 225934 311264
rect 226430 309440 226486 309496
rect 226890 306584 226946 306640
rect 229650 389272 229706 389328
rect 227810 381520 227866 381576
rect 228454 377304 228510 377360
rect 229742 369144 229798 369200
rect 228546 362208 228602 362264
rect 228270 311888 228326 311944
rect 227626 304136 227682 304192
rect 226982 303592 227038 303648
rect 227994 303592 228050 303648
rect 226890 301688 226946 301744
rect 229282 332560 229338 332616
rect 230386 333240 230442 333296
rect 230386 332560 230442 332616
rect 232594 387504 232650 387560
rect 230570 316784 230626 316840
rect 229742 308080 229798 308136
rect 235354 384376 235410 384432
rect 233146 312024 233202 312080
rect 233422 309032 233478 309088
rect 233422 307944 233478 308000
rect 234526 325080 234582 325136
rect 233974 318008 234030 318064
rect 233974 309032 234030 309088
rect 238022 356768 238078 356824
rect 237286 314064 237342 314120
rect 235998 313928 236054 313984
rect 236734 300872 236790 300928
rect 240782 389816 240838 389872
rect 239034 384240 239090 384296
rect 240046 359080 240102 359136
rect 238114 330520 238170 330576
rect 238666 313928 238722 313984
rect 238022 304272 238078 304328
rect 238206 302368 238262 302424
rect 239126 302776 239182 302832
rect 240782 305768 240838 305824
rect 242898 388592 242954 388648
rect 242898 386144 242954 386200
rect 244738 389000 244794 389056
rect 244370 384376 244426 384432
rect 244278 383016 244334 383072
rect 243082 379344 243138 379400
rect 242254 362208 242310 362264
rect 242162 305632 242218 305688
rect 242990 303728 243046 303784
rect 248878 390904 248934 390960
rect 250718 390768 250774 390824
rect 247774 389000 247830 389056
rect 248602 389000 248658 389056
rect 249246 389000 249302 389056
rect 249522 389000 249578 389056
rect 247682 384920 247738 384976
rect 247682 380840 247738 380896
rect 245658 373904 245714 373960
rect 245658 372680 245714 372736
rect 246302 372680 246358 372736
rect 244370 366832 244426 366888
rect 244830 311888 244886 311944
rect 243542 303728 243598 303784
rect 246394 362208 246450 362264
rect 246302 346976 246358 347032
rect 246394 343032 246450 343088
rect 245014 311888 245070 311944
rect 244922 303592 244978 303648
rect 246394 307128 246450 307184
rect 246946 304952 247002 305008
rect 247130 325760 247186 325816
rect 247682 307944 247738 308000
rect 252558 390904 252614 390960
rect 249246 371864 249302 371920
rect 249614 371864 249670 371920
rect 249614 364928 249670 364984
rect 249614 311208 249670 311264
rect 249062 304136 249118 304192
rect 251822 361528 251878 361584
rect 248970 302368 249026 302424
rect 249706 302368 249762 302424
rect 251914 330656 251970 330712
rect 251822 309304 251878 309360
rect 251362 306448 251418 306504
rect 250810 303728 250866 303784
rect 251914 306992 251970 307048
rect 252282 306856 252338 306912
rect 252282 302232 252338 302288
rect 249706 300872 249762 300928
rect 254214 431996 254270 432032
rect 254214 431976 254216 431996
rect 254216 431976 254268 431996
rect 254268 431976 254270 431996
rect 254214 427896 254270 427952
rect 254122 415112 254178 415168
rect 254030 392808 254086 392864
rect 254030 391992 254086 392048
rect 255410 583208 255466 583264
rect 256330 592728 256386 592784
rect 255410 579672 255466 579728
rect 255410 576952 255466 577008
rect 255410 575864 255466 575920
rect 255410 574640 255466 574696
rect 255594 574096 255650 574152
rect 255502 572872 255558 572928
rect 255410 572600 255466 572656
rect 255410 571512 255466 571568
rect 255410 570596 255412 570616
rect 255412 570596 255464 570616
rect 255464 570596 255466 570616
rect 255410 570560 255466 570596
rect 255410 569336 255466 569392
rect 255410 568656 255466 568712
rect 255778 567568 255834 567624
rect 255686 566344 255742 566400
rect 255594 565836 255596 565856
rect 255596 565836 255648 565856
rect 255648 565836 255650 565856
rect 255594 565800 255650 565836
rect 255594 564712 255650 564768
rect 255594 563100 255650 563136
rect 255594 563080 255596 563100
rect 255596 563080 255648 563100
rect 255648 563080 255650 563100
rect 255594 561856 255650 561912
rect 255594 560768 255650 560824
rect 255594 559544 255650 559600
rect 255594 557912 255650 557968
rect 255594 556824 255650 556880
rect 256606 554920 256662 554976
rect 255686 554104 255742 554160
rect 255594 553560 255650 553616
rect 255594 552744 255650 552800
rect 255594 550840 255650 550896
rect 255594 550160 255650 550216
rect 255594 548392 255650 548448
rect 255594 546760 255650 546816
rect 255594 545808 255650 545864
rect 255686 545128 255742 545184
rect 255594 544040 255650 544096
rect 255594 541184 255650 541240
rect 255594 538872 255650 538928
rect 255502 537920 255558 537976
rect 256790 551112 256846 551168
rect 257066 533296 257122 533352
rect 256790 531256 256846 531312
rect 255502 466656 255558 466712
rect 255502 465704 255558 465760
rect 255594 460264 255650 460320
rect 255594 448840 255650 448896
rect 255594 447752 255650 447808
rect 255594 447480 255650 447536
rect 255962 446120 256018 446176
rect 255502 444760 255558 444816
rect 255502 443400 255558 443456
rect 255502 442040 255558 442096
rect 255502 439048 255558 439104
rect 255502 437688 255558 437744
rect 255870 437552 255926 437608
rect 255870 436328 255926 436384
rect 255502 434968 255558 435024
rect 255502 433608 255558 433664
rect 255410 430616 255466 430672
rect 255410 429256 255466 429312
rect 255410 426536 255466 426592
rect 256606 425176 256662 425232
rect 255502 423544 255558 423600
rect 255502 422184 255558 422240
rect 255502 420824 255558 420880
rect 255410 419484 255466 419520
rect 255410 419464 255412 419484
rect 255412 419464 255464 419484
rect 255464 419464 255466 419484
rect 255502 418104 255558 418160
rect 255410 416764 255466 416800
rect 255410 416744 255412 416764
rect 255412 416744 255464 416764
rect 255464 416744 255466 416764
rect 255318 415112 255374 415168
rect 255502 412392 255558 412448
rect 255502 411032 255558 411088
rect 255410 409672 255466 409728
rect 255410 408312 255466 408368
rect 255502 406952 255558 407008
rect 254214 388456 254270 388512
rect 254214 388048 254270 388104
rect 253938 375264 253994 375320
rect 253202 334600 253258 334656
rect 255410 403960 255466 404016
rect 255410 402600 255466 402656
rect 255410 401240 255466 401296
rect 255410 399880 255466 399936
rect 255410 395528 255466 395584
rect 255410 394168 255466 394224
rect 254122 375264 254178 375320
rect 253294 329160 253350 329216
rect 252466 311208 252522 311264
rect 192482 291760 192538 291816
rect 193126 283464 193182 283520
rect 192022 263880 192078 263936
rect 191746 247560 191802 247616
rect 191286 244296 191342 244352
rect 191654 244296 191710 244352
rect 191838 242800 191894 242856
rect 191746 242120 191802 242176
rect 191286 235184 191342 235240
rect 189078 152360 189134 152416
rect 188434 92248 188490 92304
rect 188526 91160 188582 91216
rect 190366 138624 190422 138680
rect 190274 138488 190330 138544
rect 189998 136720 190054 136776
rect 189906 133864 189962 133920
rect 190274 129784 190330 129840
rect 193678 244160 193734 244216
rect 193586 242392 193642 242448
rect 194506 241984 194562 242040
rect 193678 241304 193734 241360
rect 192482 157936 192538 157992
rect 190458 134680 190514 134736
rect 192482 149096 192538 149152
rect 191746 136312 191802 136368
rect 191746 135496 191802 135552
rect 192942 139848 192998 139904
rect 191746 134408 191802 134464
rect 192482 134408 192538 134464
rect 190458 125704 190514 125760
rect 190274 110744 190330 110800
rect 189722 95240 189778 95296
rect 189814 89528 189870 89584
rect 189078 83680 189134 83736
rect 189078 82864 189134 82920
rect 189722 82864 189778 82920
rect 190458 121624 190514 121680
rect 191654 131144 191710 131200
rect 193034 131960 193090 132016
rect 191654 129240 191710 129296
rect 191746 128424 191802 128480
rect 192298 127608 192354 127664
rect 192390 126520 192446 126576
rect 191746 122984 191802 123040
rect 191194 121388 191196 121408
rect 191196 121388 191248 121408
rect 191248 121388 191250 121408
rect 191194 121352 191250 121388
rect 191746 120264 191802 120320
rect 191746 119448 191802 119504
rect 191746 118632 191802 118688
rect 191102 117544 191158 117600
rect 191286 116728 191342 116784
rect 191746 115912 191802 115968
rect 191010 115096 191066 115152
rect 191746 114008 191802 114064
rect 191194 113228 191196 113248
rect 191196 113228 191248 113248
rect 191248 113228 191250 113248
rect 191194 113192 191250 113228
rect 191378 110472 191434 110528
rect 191562 109656 191618 109712
rect 191194 108876 191196 108896
rect 191196 108876 191248 108896
rect 191248 108876 191250 108896
rect 191194 108840 191250 108876
rect 191194 107772 191250 107808
rect 191194 107752 191196 107772
rect 191196 107752 191248 107772
rect 191248 107752 191250 107772
rect 191746 106936 191802 106992
rect 191746 106120 191802 106176
rect 191746 105032 191802 105088
rect 191746 104216 191802 104272
rect 191654 103400 191710 103456
rect 191102 102584 191158 102640
rect 190642 99864 190698 99920
rect 190642 97144 190698 97200
rect 191654 101496 191710 101552
rect 191562 100680 191618 100736
rect 191562 99456 191618 99512
rect 191102 93880 191158 93936
rect 191102 85312 191158 85368
rect 191654 97960 191710 98016
rect 191654 94424 191710 94480
rect 191562 83408 191618 83464
rect 191746 93608 191802 93664
rect 191102 77152 191158 77208
rect 191654 77152 191710 77208
rect 193034 126520 193090 126576
rect 192942 124888 192998 124944
rect 191102 62056 191158 62112
rect 193218 157392 193274 157448
rect 196622 241032 196678 241088
rect 194506 238040 194562 238096
rect 197358 237904 197414 237960
rect 196714 236000 196770 236056
rect 196622 234504 196678 234560
rect 197358 233144 197414 233200
rect 198646 233144 198702 233200
rect 195978 214512 196034 214568
rect 196622 214512 196678 214568
rect 193770 182824 193826 182880
rect 193862 157392 193918 157448
rect 196070 157392 196126 157448
rect 196622 157392 196678 157448
rect 193310 142840 193366 142896
rect 194690 142704 194746 142760
rect 194690 142160 194746 142216
rect 197266 163376 197322 163432
rect 196622 142296 196678 142352
rect 200762 236544 200818 236600
rect 198646 158072 198702 158128
rect 203614 232464 203670 232520
rect 203614 227568 203670 227624
rect 204902 216552 204958 216608
rect 204902 215328 204958 215384
rect 205546 215328 205602 215384
rect 200762 153720 200818 153776
rect 201590 148280 201646 148336
rect 196806 140392 196862 140448
rect 207018 177248 207074 177304
rect 205822 176704 205878 176760
rect 207018 176704 207074 176760
rect 207662 176704 207718 176760
rect 205546 155896 205602 155952
rect 204442 149640 204498 149696
rect 204258 141072 204314 141128
rect 205454 140936 205510 140992
rect 207110 145016 207166 145072
rect 207018 143248 207074 143304
rect 211802 239944 211858 240000
rect 211802 224168 211858 224224
rect 210422 222128 210478 222184
rect 211066 222128 211122 222184
rect 210422 171128 210478 171184
rect 208490 151136 208546 151192
rect 208122 143248 208178 143304
rect 202878 140392 202934 140448
rect 203522 140392 203578 140448
rect 209502 140528 209558 140584
rect 210514 144064 210570 144120
rect 213274 222264 213330 222320
rect 211802 189624 211858 189680
rect 211158 156032 211214 156088
rect 211066 151000 211122 151056
rect 211802 149640 211858 149696
rect 214654 192480 214710 192536
rect 213274 159296 213330 159352
rect 212814 142432 212870 142488
rect 216678 238040 216734 238096
rect 215390 237904 215446 237960
rect 216678 237224 216734 237280
rect 217966 237224 218022 237280
rect 215942 164328 215998 164384
rect 215298 153856 215354 153912
rect 211894 140664 211950 140720
rect 208214 140392 208270 140448
rect 220082 210840 220138 210896
rect 222198 230424 222254 230480
rect 220082 167048 220138 167104
rect 219438 149504 219494 149560
rect 218334 147736 218390 147792
rect 218242 143384 218298 143440
rect 220174 149504 220230 149560
rect 218794 146376 218850 146432
rect 220082 146376 220138 146432
rect 220174 141072 220230 141128
rect 222198 154672 222254 154728
rect 221922 142296 221978 142352
rect 219990 140800 220046 140856
rect 223762 141344 223818 141400
rect 225050 136584 225106 136640
rect 193218 124072 193274 124128
rect 225234 123800 225290 123856
rect 226338 139032 226394 139088
rect 226338 136312 226394 136368
rect 226338 133320 226394 133376
rect 226338 131960 226394 132016
rect 226338 126520 226394 126576
rect 226522 124616 226578 124672
rect 226338 122984 226394 123040
rect 226338 122168 226394 122224
rect 226430 120264 226486 120320
rect 226522 118360 226578 118416
rect 226338 114824 226394 114880
rect 226338 111288 226394 111344
rect 226522 110472 226578 110528
rect 225142 109656 225198 109712
rect 193218 104216 193274 104272
rect 193126 96328 193182 96384
rect 199106 93336 199162 93392
rect 205730 93336 205786 93392
rect 194690 85448 194746 85504
rect 195886 85448 195942 85504
rect 196530 92656 196586 92712
rect 196070 88204 196072 88224
rect 196072 88204 196124 88224
rect 196124 88204 196126 88224
rect 196070 88168 196126 88204
rect 197082 87896 197138 87952
rect 195886 78512 195942 78568
rect 200394 92792 200450 92848
rect 200210 92384 200266 92440
rect 200946 92384 201002 92440
rect 202602 92112 202658 92168
rect 200762 71712 200818 71768
rect 203338 92792 203394 92848
rect 208950 93336 209006 93392
rect 211710 93336 211766 93392
rect 224774 93336 224830 93392
rect 212446 92928 212502 92984
rect 203706 90480 203762 90536
rect 204442 90344 204498 90400
rect 205086 91024 205142 91080
rect 204994 89664 205050 89720
rect 204442 86808 204498 86864
rect 205546 79328 205602 79384
rect 205546 78648 205602 78704
rect 209226 88032 209282 88088
rect 210514 89392 210570 89448
rect 211066 89392 211122 89448
rect 210330 86672 210386 86728
rect 210238 85312 210294 85368
rect 212446 82048 212502 82104
rect 215298 90208 215354 90264
rect 216402 90208 216458 90264
rect 215206 62736 215262 62792
rect 218794 90888 218850 90944
rect 219622 81368 219678 81424
rect 220082 75792 220138 75848
rect 224038 92792 224094 92848
rect 224314 90616 224370 90672
rect 225050 104896 225106 104952
rect 225142 97144 225198 97200
rect 225142 92248 225198 92304
rect 226522 107752 226578 107808
rect 226522 104216 226578 104272
rect 226338 101496 226394 101552
rect 226338 100680 226394 100736
rect 226430 99592 226486 99648
rect 226338 98776 226394 98832
rect 225602 90888 225658 90944
rect 226338 82728 226394 82784
rect 226522 96056 226578 96112
rect 226522 95240 226578 95296
rect 231122 236680 231178 236736
rect 228362 230016 228418 230072
rect 227718 160112 227774 160168
rect 226706 137128 226762 137184
rect 226706 135496 226762 135552
rect 226706 134680 226762 134736
rect 226706 133592 226762 133648
rect 226706 130872 226762 130928
rect 226798 130056 226854 130112
rect 226706 128424 226762 128480
rect 226706 127336 226762 127392
rect 227718 125704 227774 125760
rect 226706 117544 226762 117600
rect 226706 115948 226708 115968
rect 226708 115948 226760 115968
rect 226760 115948 226762 115968
rect 226706 115912 226762 115948
rect 227626 113736 227682 113792
rect 229098 165688 229154 165744
rect 228362 160112 228418 160168
rect 227994 139848 228050 139904
rect 227994 129240 228050 129296
rect 230018 150456 230074 150512
rect 229742 144880 229798 144936
rect 230478 146512 230534 146568
rect 227902 116728 227958 116784
rect 226706 112104 226762 112160
rect 226706 106936 226762 106992
rect 226706 105848 226762 105904
rect 226706 103400 226762 103456
rect 226706 102312 226762 102368
rect 227074 108568 227130 108624
rect 226982 98776 227038 98832
rect 226614 94444 226670 94480
rect 226614 94424 226616 94444
rect 226616 94424 226668 94444
rect 226668 94424 226670 94444
rect 227626 93608 227682 93664
rect 226522 88168 226578 88224
rect 227902 98640 227958 98696
rect 227902 97960 227958 98016
rect 227902 89528 227958 89584
rect 228362 83408 228418 83464
rect 231950 229744 232006 229800
rect 231858 221992 231914 222048
rect 231214 142296 231270 142352
rect 234618 241304 234674 241360
rect 235538 241304 235594 241360
rect 233146 221992 233202 222048
rect 233882 213152 233938 213208
rect 231950 162832 232006 162888
rect 231858 92792 231914 92848
rect 231306 85312 231362 85368
rect 233330 153720 233386 153776
rect 233330 138896 233386 138952
rect 233330 138624 233386 138680
rect 237378 235728 237434 235784
rect 234618 158752 234674 158808
rect 234618 141344 234674 141400
rect 233882 117136 233938 117192
rect 235998 228248 236054 228304
rect 236642 226888 236698 226944
rect 236642 206896 236698 206952
rect 236090 162696 236146 162752
rect 236642 162696 236698 162752
rect 236090 161472 236146 161528
rect 237378 98676 237380 98696
rect 237380 98676 237432 98696
rect 237432 98676 237434 98696
rect 237378 98640 237434 98676
rect 240046 149096 240102 149152
rect 243542 240896 243598 240952
rect 239402 148280 239458 148336
rect 237654 85448 237710 85504
rect 238482 85448 238538 85504
rect 240322 156576 240378 156632
rect 240874 90616 240930 90672
rect 244370 153040 244426 153096
rect 244370 151816 244426 151872
rect 245014 153040 245070 153096
rect 246302 239536 246358 239592
rect 245106 146240 245162 146296
rect 247498 239400 247554 239456
rect 247038 234368 247094 234424
rect 248326 228384 248382 228440
rect 248326 224848 248382 224904
rect 249062 224848 249118 224904
rect 247038 217268 247040 217288
rect 247040 217268 247092 217288
rect 247092 217268 247094 217288
rect 247038 217232 247094 217268
rect 248326 217232 248382 217288
rect 248970 174528 249026 174584
rect 250166 241984 250222 242040
rect 251822 239808 251878 239864
rect 250534 239400 250590 239456
rect 250442 235184 250498 235240
rect 250534 210976 250590 211032
rect 252466 239672 252522 239728
rect 250442 92384 250498 92440
rect 253202 303592 253258 303648
rect 252926 301552 252982 301608
rect 254030 319368 254086 319424
rect 253018 299784 253074 299840
rect 253294 299784 253350 299840
rect 252834 298968 252890 299024
rect 252834 298016 252890 298072
rect 252834 293392 252890 293448
rect 253938 295604 253940 295624
rect 253940 295604 253992 295624
rect 253992 295604 253994 295624
rect 253938 295568 253994 295604
rect 253202 292848 253258 292904
rect 253018 244432 253074 244488
rect 252926 242800 252982 242856
rect 252926 241984 252982 242040
rect 254582 317328 254638 317384
rect 254122 315288 254178 315344
rect 254030 253952 254086 254008
rect 254030 251504 254086 251560
rect 254214 302232 254270 302288
rect 255318 296112 255374 296168
rect 255318 295432 255374 295488
rect 255318 294344 255374 294400
rect 256882 440408 256938 440464
rect 256882 394576 256938 394632
rect 255502 300736 255558 300792
rect 255594 300328 255650 300384
rect 255502 299104 255558 299160
rect 255870 298696 255926 298752
rect 255594 298560 255650 298616
rect 255502 298172 255558 298208
rect 255502 298152 255504 298172
rect 255504 298152 255556 298172
rect 255556 298152 255558 298172
rect 255502 296928 255558 296984
rect 255502 296556 255504 296576
rect 255504 296556 255556 296576
rect 255556 296556 255558 296576
rect 255502 296520 255558 296556
rect 255410 293972 255412 293992
rect 255412 293972 255464 293992
rect 255464 293972 255466 293992
rect 255410 293936 255466 293972
rect 255318 293120 255374 293176
rect 255410 292576 255466 292632
rect 255502 282376 255558 282432
rect 255410 281968 255466 282024
rect 255410 281460 255412 281480
rect 255412 281460 255464 281480
rect 255464 281460 255466 281480
rect 255410 281424 255466 281460
rect 255502 280200 255558 280256
rect 255410 278976 255466 279032
rect 255410 278432 255466 278488
rect 255502 277616 255558 277672
rect 255502 277208 255558 277264
rect 255410 276392 255466 276448
rect 255502 275440 255558 275496
rect 255410 275032 255466 275088
rect 255410 274216 255466 274272
rect 255502 273808 255558 273864
rect 255410 273128 255466 273184
rect 255502 272448 255558 272504
rect 255410 272040 255466 272096
rect 255502 271768 255558 271824
rect 255318 271632 255374 271688
rect 255410 271224 255466 271280
rect 255502 270816 255558 270872
rect 255318 270544 255374 270600
rect 255410 269864 255466 269920
rect 255502 269048 255558 269104
rect 255410 267844 255466 267880
rect 255410 267824 255412 267844
rect 255412 267824 255464 267844
rect 255464 267824 255466 267844
rect 255410 267416 255466 267472
rect 255318 266056 255374 266112
rect 255410 265648 255466 265704
rect 255502 264288 255558 264344
rect 255410 263880 255466 263936
rect 255502 263064 255558 263120
rect 255410 262268 255466 262304
rect 255410 262248 255412 262268
rect 255412 262248 255464 262268
rect 255464 262248 255466 262268
rect 255410 261840 255466 261896
rect 255318 261024 255374 261080
rect 255502 260888 255558 260944
rect 255410 260500 255466 260536
rect 255410 260480 255412 260500
rect 255412 260480 255464 260500
rect 255464 260480 255466 260500
rect 255318 259664 255374 259720
rect 255410 258304 255466 258360
rect 255318 257488 255374 257544
rect 255410 257080 255466 257136
rect 255502 256264 255558 256320
rect 255410 255332 255466 255368
rect 255410 255312 255412 255332
rect 255412 255312 255464 255332
rect 255464 255312 255466 255332
rect 255502 254904 255558 254960
rect 255410 254532 255412 254552
rect 255412 254532 255464 254552
rect 255464 254532 255466 254552
rect 255410 254496 255466 254532
rect 255502 253272 255558 253328
rect 255410 252748 255466 252784
rect 255410 252728 255412 252748
rect 255412 252728 255464 252748
rect 255464 252728 255466 252748
rect 254950 252456 255006 252512
rect 255410 251912 255466 251968
rect 254950 251504 255006 251560
rect 254214 249736 254270 249792
rect 255502 251096 255558 251152
rect 255410 250280 255466 250336
rect 255502 249328 255558 249384
rect 255410 248920 255466 248976
rect 255318 248512 255374 248568
rect 255502 248376 255558 248432
rect 255502 248104 255558 248160
rect 255410 247716 255466 247752
rect 255410 247696 255412 247716
rect 255412 247696 255464 247716
rect 255464 247696 255466 247716
rect 255502 246744 255558 246800
rect 254122 246336 254178 246392
rect 255318 246336 255374 246392
rect 254122 243752 254178 243808
rect 254214 242528 254270 242584
rect 254122 239536 254178 239592
rect 255410 245556 255412 245576
rect 255412 245556 255464 245576
rect 255464 245556 255466 245576
rect 255410 245520 255466 245556
rect 255410 245112 255466 245168
rect 255502 244160 255558 244216
rect 254214 237904 254270 237960
rect 256054 297744 256110 297800
rect 255870 297336 255926 297392
rect 255686 295432 255742 295488
rect 258262 525000 258318 525056
rect 257342 454008 257398 454064
rect 257066 353912 257122 353968
rect 258998 398520 259054 398576
rect 258170 390768 258226 390824
rect 259274 384784 259330 384840
rect 262218 598984 262274 599040
rect 259642 458496 259698 458552
rect 259550 383016 259606 383072
rect 259458 351736 259514 351792
rect 256698 295024 256754 295080
rect 256698 294752 256754 294808
rect 256790 293528 256846 293584
rect 256606 292168 256662 292224
rect 256606 291760 256662 291816
rect 256514 290944 256570 291000
rect 256514 290536 256570 290592
rect 256514 289584 256570 289640
rect 256606 289176 256662 289232
rect 255870 287952 255926 288008
rect 255962 287544 256018 287600
rect 255870 286592 255926 286648
rect 256514 286184 256570 286240
rect 256606 285368 256662 285424
rect 255778 283600 255834 283656
rect 256422 283192 256478 283248
rect 255778 271088 255834 271144
rect 255778 268232 255834 268288
rect 255870 243344 255926 243400
rect 256606 220088 256662 220144
rect 256606 219272 256662 219328
rect 252834 154536 252890 154592
rect 252742 114416 252798 114472
rect 253018 114416 253074 114472
rect 253018 113192 253074 113248
rect 256146 203496 256202 203552
rect 256974 305768 257030 305824
rect 256974 288360 257030 288416
rect 257986 288360 258042 288416
rect 257986 287680 258042 287736
rect 256882 278024 256938 278080
rect 259274 302368 259330 302424
rect 258722 302232 258778 302288
rect 259274 298016 259330 298072
rect 259458 302232 259514 302288
rect 258722 282240 258778 282296
rect 256882 266872 256938 266928
rect 256790 243208 256846 243264
rect 256790 242256 256846 242312
rect 258078 258168 258134 258224
rect 256790 236544 256846 236600
rect 258078 255720 258134 255776
rect 258170 246200 258226 246256
rect 258262 240760 258318 240816
rect 258170 228384 258226 228440
rect 256146 168952 256202 169008
rect 256698 95784 256754 95840
rect 259366 283464 259422 283520
rect 259366 282784 259422 282840
rect 259642 301416 259698 301472
rect 259458 282240 259514 282296
rect 260286 346976 260342 347032
rect 260194 319368 260250 319424
rect 260930 341400 260986 341456
rect 260286 311344 260342 311400
rect 259826 296656 259882 296712
rect 262310 452784 262366 452840
rect 262218 389000 262274 389056
rect 260102 282104 260158 282160
rect 259642 281016 259698 281072
rect 259458 279792 259514 279848
rect 259642 266464 259698 266520
rect 261022 300600 261078 300656
rect 260746 263472 260802 263528
rect 260746 260500 260802 260536
rect 260746 260480 260748 260500
rect 260748 260480 260800 260500
rect 260800 260480 260802 260500
rect 258722 113192 258778 113248
rect 261206 291216 261262 291272
rect 261114 253952 261170 254008
rect 261114 239400 261170 239456
rect 263782 460944 263838 461000
rect 262310 347792 262366 347848
rect 262218 285232 262274 285288
rect 262218 283872 262274 283928
rect 262494 303628 262496 303648
rect 262496 303628 262548 303648
rect 262548 303628 262550 303648
rect 262494 303592 262550 303628
rect 262862 299512 262918 299568
rect 263138 285232 263194 285288
rect 263138 284280 263194 284336
rect 262586 281016 262642 281072
rect 262310 277072 262366 277128
rect 262402 270544 262458 270600
rect 262218 270408 262274 270464
rect 262218 270136 262274 270192
rect 261482 262248 261538 262304
rect 262494 228248 262550 228304
rect 263690 284280 263746 284336
rect 265254 480800 265310 480856
rect 265162 387640 265218 387696
rect 265070 359352 265126 359408
rect 264978 318008 265034 318064
rect 263966 279656 264022 279712
rect 263874 262656 263930 262712
rect 263874 216552 263930 216608
rect 265714 387640 265770 387696
rect 266542 386144 266598 386200
rect 266450 335960 266506 336016
rect 267002 386144 267058 386200
rect 267738 369144 267794 369200
rect 267830 368328 267886 368384
rect 267738 334056 267794 334112
rect 265622 298016 265678 298072
rect 265254 260208 265310 260264
rect 265162 259120 265218 259176
rect 265070 252048 265126 252104
rect 265070 247716 265126 247752
rect 265070 247696 265072 247716
rect 265072 247696 265124 247716
rect 265124 247696 265126 247716
rect 262218 79464 262274 79520
rect 265070 206932 265072 206952
rect 265072 206932 265124 206952
rect 265124 206932 265126 206952
rect 265070 206896 265126 206932
rect 266450 295024 266506 295080
rect 266358 284280 266414 284336
rect 266634 285776 266690 285832
rect 267738 322088 267794 322144
rect 267738 306992 267794 307048
rect 267738 287680 267794 287736
rect 266726 284280 266782 284336
rect 266542 269320 266598 269376
rect 266634 252184 266690 252240
rect 266542 238584 266598 238640
rect 267094 235184 267150 235240
rect 266634 233144 266690 233200
rect 267094 204176 267150 204232
rect 268014 392536 268070 392592
rect 268014 341400 268070 341456
rect 267922 323584 267978 323640
rect 269394 465976 269450 466032
rect 269118 314064 269174 314120
rect 267002 140936 267058 140992
rect 267922 250008 267978 250064
rect 269118 285640 269174 285696
rect 268290 262384 268346 262440
rect 268382 142432 268438 142488
rect 271142 536560 271198 536616
rect 270590 451288 270646 451344
rect 269394 389816 269450 389872
rect 269762 311208 269818 311264
rect 269762 283600 269818 283656
rect 270774 362888 270830 362944
rect 270590 282104 270646 282160
rect 270590 281424 270646 281480
rect 270590 280608 270646 280664
rect 270498 274624 270554 274680
rect 269394 272448 269450 272504
rect 270406 244160 270462 244216
rect 269394 235864 269450 235920
rect 270682 273808 270738 273864
rect 270590 226208 270646 226264
rect 270590 222128 270646 222184
rect 271878 357992 271934 358048
rect 273350 465024 273406 465080
rect 273626 449928 273682 449984
rect 273442 379208 273498 379264
rect 273442 378936 273498 378992
rect 272062 346432 272118 346488
rect 270774 271088 270830 271144
rect 270774 248376 270830 248432
rect 273442 303864 273498 303920
rect 273258 281424 273314 281480
rect 273258 275984 273314 276040
rect 272062 273128 272118 273184
rect 273626 269320 273682 269376
rect 278042 601840 278098 601896
rect 276018 599120 276074 599176
rect 276018 468424 276074 468480
rect 276294 458360 276350 458416
rect 276110 382880 276166 382936
rect 276018 376624 276074 376680
rect 274914 331744 274970 331800
rect 276018 309032 276074 309088
rect 276018 307808 276074 307864
rect 274914 283464 274970 283520
rect 274822 279384 274878 279440
rect 276018 275984 276074 276040
rect 277490 369008 277546 369064
rect 276294 309032 276350 309088
rect 276110 271768 276166 271824
rect 274822 265512 274878 265568
rect 274730 257896 274786 257952
rect 270498 97416 270554 97472
rect 269026 3440 269082 3496
rect 273258 80688 273314 80744
rect 277858 386280 277914 386336
rect 278962 469240 279018 469296
rect 279330 416608 279386 416664
rect 278778 309168 278834 309224
rect 278778 298696 278834 298752
rect 277674 271768 277730 271824
rect 277674 209616 277730 209672
rect 277398 86808 277454 86864
rect 274822 3440 274878 3496
rect 278686 86808 278742 86864
rect 278686 85584 278742 85640
rect 278962 309168 279018 309224
rect 278962 262112 279018 262168
rect 280802 536424 280858 536480
rect 280434 380704 280490 380760
rect 280158 271088 280214 271144
rect 279422 246200 279478 246256
rect 280158 227568 280214 227624
rect 278778 77152 278834 77208
rect 280066 77152 280122 77208
rect 281814 456864 281870 456920
rect 283102 450064 283158 450120
rect 283010 385600 283066 385656
rect 282918 311072 282974 311128
rect 282918 273808 282974 273864
rect 281722 262792 281778 262848
rect 288714 604696 288770 604752
rect 289726 604696 289782 604752
rect 285678 466520 285734 466576
rect 285678 462848 285734 462904
rect 284482 456048 284538 456104
rect 284298 373224 284354 373280
rect 283102 253816 283158 253872
rect 284482 320184 284538 320240
rect 284482 262248 284538 262304
rect 284298 242120 284354 242176
rect 281630 151136 281686 151192
rect 284482 213152 284538 213208
rect 285126 263472 285182 263528
rect 285126 262248 285182 262304
rect 287610 472096 287666 472152
rect 287334 455504 287390 455560
rect 288346 455504 288402 455560
rect 287242 454688 287298 454744
rect 287150 301008 287206 301064
rect 285862 257216 285918 257272
rect 285126 216688 285182 216744
rect 285770 144064 285826 144120
rect 288530 463664 288586 463720
rect 287150 78512 287206 78568
rect 284942 74432 284998 74488
rect 284298 73208 284354 73264
rect 284942 73208 284998 73264
rect 289818 459584 289874 459640
rect 288622 377984 288678 378040
rect 288530 264152 288586 264208
rect 288714 263472 288770 263528
rect 289910 390496 289966 390552
rect 289910 389136 289966 389192
rect 291198 384920 291254 384976
rect 291382 471960 291438 472016
rect 291382 382200 291438 382256
rect 291198 311888 291254 311944
rect 288438 79328 288494 79384
rect 288346 78512 288402 78568
rect 291290 307944 291346 308000
rect 291474 376488 291530 376544
rect 296810 453192 296866 453248
rect 295338 437552 295394 437608
rect 293958 338680 294014 338736
rect 292670 282104 292726 282160
rect 291382 268504 291438 268560
rect 295522 309304 295578 309360
rect 295338 260072 295394 260128
rect 291290 117136 291346 117192
rect 291658 117136 291714 117192
rect 296718 306448 296774 306504
rect 582470 697176 582526 697232
rect 582378 617480 582434 617536
rect 582378 590960 582434 591016
rect 582378 577632 582434 577688
rect 582562 683848 582618 683904
rect 582654 644000 582710 644056
rect 582746 630808 582802 630864
rect 582930 670656 582986 670712
rect 582838 609184 582894 609240
rect 582746 607824 582802 607880
rect 582654 603608 582710 603664
rect 582746 601704 582802 601760
rect 582470 537784 582526 537840
rect 579802 484608 579858 484664
rect 299478 329024 299534 329080
rect 580170 458088 580226 458144
rect 582838 564304 582894 564360
rect 582930 538192 582986 538248
rect 582746 524456 582802 524512
rect 582654 511264 582710 511320
rect 582378 418240 582434 418296
rect 582654 471416 582710 471472
rect 582470 404912 582526 404968
rect 582378 378392 582434 378448
rect 582470 365064 582526 365120
rect 302330 304952 302386 305008
rect 582378 302776 582434 302832
rect 580170 272176 580226 272232
rect 580906 258848 580962 258904
rect 580170 232328 580226 232384
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192500 580226 192536
rect 580170 192480 580172 192500
rect 580172 192480 580224 192500
rect 580224 192480 580226 192500
rect 580170 179152 580226 179208
rect 316038 159296 316094 159352
rect 303618 157392 303674 157448
rect 299570 39208 299626 39264
rect 300858 26832 300914 26888
rect 302974 21256 303030 21312
rect 304262 3984 304318 4040
rect 307942 3984 307998 4040
rect 338118 87488 338174 87544
rect 335358 65456 335414 65512
rect 341522 3304 341578 3360
rect 350446 3304 350502 3360
rect 353298 82048 353354 82104
rect 580262 72936 580318 72992
rect 580170 46280 580226 46336
rect 582746 431568 582802 431624
rect 582746 390496 582802 390552
rect 582562 351872 582618 351928
rect 582654 312024 582710 312080
rect 582470 251776 582526 251832
rect 582470 248376 582526 248432
rect 582470 245520 582526 245576
rect 582654 152632 582710 152688
rect 582654 138624 582710 138680
rect 582838 165824 582894 165880
rect 583114 146376 583170 146432
rect 583022 139304 583078 139360
rect 582930 125976 582986 126032
rect 583114 112784 583170 112840
rect 583022 99456 583078 99512
rect 582746 59608 582802 59664
rect 582654 19760 582710 19816
rect 582930 33088 582986 33144
rect 582838 6568 582894 6624
<< metal3 >>
rect -960 697220 480 697460
rect 582465 697234 582531 697237
rect 583520 697234 584960 697324
rect 582465 697232 584960 697234
rect 582465 697176 582470 697232
rect 582526 697176 584960 697232
rect 582465 697174 584960 697176
rect 582465 697171 582531 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582557 683906 582623 683909
rect 583520 683906 584960 683996
rect 582557 683904 584960 683906
rect 582557 683848 582562 683904
rect 582618 683848 584960 683904
rect 582557 683846 584960 683848
rect 582557 683843 582623 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582925 670714 582991 670717
rect 583520 670714 584960 670804
rect 582925 670712 584960 670714
rect 582925 670656 582930 670712
rect 582986 670656 584960 670712
rect 582925 670654 584960 670656
rect 582925 670651 582991 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582649 644058 582715 644061
rect 583520 644058 584960 644148
rect 582649 644056 584960 644058
rect 582649 644000 582654 644056
rect 582710 644000 584960 644056
rect 582649 643998 584960 644000
rect 582649 643995 582715 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582741 630866 582807 630869
rect 583520 630866 584960 630956
rect 582741 630864 584960 630866
rect 582741 630808 582746 630864
rect 582802 630808 584960 630864
rect 582741 630806 584960 630808
rect 582741 630803 582807 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582373 617538 582439 617541
rect 583520 617538 584960 617628
rect 582373 617536 584960 617538
rect 582373 617480 582378 617536
rect 582434 617480 584960 617536
rect 582373 617478 584960 617480
rect 582373 617475 582439 617478
rect 583520 617388 584960 617478
rect 189717 612778 189783 612781
rect 222193 612778 222259 612781
rect 222837 612778 222903 612781
rect 189717 612776 222903 612778
rect 189717 612720 189722 612776
rect 189778 612720 222198 612776
rect 222254 612720 222842 612776
rect 222898 612720 222903 612776
rect 189717 612718 222903 612720
rect 189717 612715 189783 612718
rect 222193 612715 222259 612718
rect 222837 612715 222903 612718
rect 173801 611418 173867 611421
rect 204345 611418 204411 611421
rect 173801 611416 204411 611418
rect 173801 611360 173806 611416
rect 173862 611360 204350 611416
rect 204406 611360 204411 611416
rect 173801 611358 204411 611360
rect 173801 611355 173867 611358
rect 204345 611355 204411 611358
rect 143441 610058 143507 610061
rect 202873 610058 202939 610061
rect 143441 610056 202939 610058
rect 143441 610000 143446 610056
rect 143502 610000 202878 610056
rect 202934 610000 202939 610056
rect 143441 609998 202939 610000
rect 143441 609995 143507 609998
rect 202873 609995 202939 609998
rect 218237 609242 218303 609245
rect 582833 609242 582899 609245
rect 218237 609240 582899 609242
rect 218237 609184 218242 609240
rect 218298 609184 582838 609240
rect 582894 609184 582899 609240
rect 218237 609182 582899 609184
rect 218237 609179 218303 609182
rect 582833 609179 582899 609182
rect 160737 608698 160803 608701
rect 198733 608698 198799 608701
rect 160737 608696 198799 608698
rect 160737 608640 160742 608696
rect 160798 608640 198738 608696
rect 198794 608640 198799 608696
rect 160737 608638 198799 608640
rect 160737 608635 160803 608638
rect 198733 608635 198799 608638
rect 191649 607882 191715 607885
rect 582741 607882 582807 607885
rect 191649 607880 582807 607882
rect 191649 607824 191654 607880
rect 191710 607824 582746 607880
rect 582802 607824 582807 607880
rect 191649 607822 582807 607824
rect 191649 607819 191715 607822
rect 582741 607819 582807 607822
rect 155861 607338 155927 607341
rect 234061 607338 234127 607341
rect 155861 607336 234127 607338
rect 155861 607280 155866 607336
rect 155922 607280 234066 607336
rect 234122 607280 234127 607336
rect 155861 607278 234127 607280
rect 155861 607275 155927 607278
rect 234061 607275 234127 607278
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 239213 606114 239279 606117
rect 259494 606114 259500 606116
rect 239213 606112 259500 606114
rect 239213 606056 239218 606112
rect 239274 606056 259500 606112
rect 239213 606054 259500 606056
rect 239213 606051 239279 606054
rect 259494 606052 259500 606054
rect 259564 606052 259570 606116
rect 144729 605978 144795 605981
rect 245469 605978 245535 605981
rect 144729 605976 245535 605978
rect 144729 605920 144734 605976
rect 144790 605920 245474 605976
rect 245530 605920 245535 605976
rect 144729 605918 245535 605920
rect 144729 605915 144795 605918
rect 245469 605915 245535 605918
rect 196709 604754 196775 604757
rect 288709 604754 288775 604757
rect 289721 604754 289787 604757
rect 196709 604752 289787 604754
rect 196709 604696 196714 604752
rect 196770 604696 288714 604752
rect 288770 604696 289726 604752
rect 289782 604696 289787 604752
rect 196709 604694 289787 604696
rect 196709 604691 196775 604694
rect 288709 604691 288775 604694
rect 289721 604691 289787 604694
rect 188286 604556 188292 604620
rect 188356 604618 188362 604620
rect 199837 604618 199903 604621
rect 188356 604616 199903 604618
rect 188356 604560 199842 604616
rect 199898 604560 199903 604616
rect 188356 604558 199903 604560
rect 188356 604556 188362 604558
rect 199837 604555 199903 604558
rect 115289 604482 115355 604485
rect 238477 604482 238543 604485
rect 115289 604480 238543 604482
rect 115289 604424 115294 604480
rect 115350 604424 238482 604480
rect 238538 604424 238543 604480
rect 115289 604422 238543 604424
rect 115289 604419 115355 604422
rect 238477 604419 238543 604422
rect 583520 604060 584960 604300
rect 191189 603666 191255 603669
rect 582649 603666 582715 603669
rect 191189 603664 582715 603666
rect 191189 603608 191194 603664
rect 191250 603608 582654 603664
rect 582710 603608 582715 603664
rect 191189 603606 582715 603608
rect 191189 603603 191255 603606
rect 582649 603603 582715 603606
rect 155718 603196 155724 603260
rect 155788 603258 155794 603260
rect 208669 603258 208735 603261
rect 155788 603256 208735 603258
rect 155788 603200 208674 603256
rect 208730 603200 208735 603256
rect 155788 603198 208735 603200
rect 155788 603196 155794 603198
rect 208669 603195 208735 603198
rect 66161 603122 66227 603125
rect 255313 603122 255379 603125
rect 66161 603120 255379 603122
rect 66161 603064 66166 603120
rect 66222 603064 255318 603120
rect 255374 603064 255379 603120
rect 66161 603062 255379 603064
rect 66161 603059 66227 603062
rect 255313 603059 255379 603062
rect 185577 602034 185643 602037
rect 211613 602034 211679 602037
rect 185577 602032 211679 602034
rect 185577 601976 185582 602032
rect 185638 601976 211618 602032
rect 211674 601976 211679 602032
rect 185577 601974 211679 601976
rect 185577 601971 185643 601974
rect 211613 601971 211679 601974
rect 88977 601898 89043 601901
rect 229645 601898 229711 601901
rect 278037 601898 278103 601901
rect 88977 601896 278103 601898
rect 88977 601840 88982 601896
rect 89038 601840 229650 601896
rect 229706 601840 278042 601896
rect 278098 601840 278103 601896
rect 88977 601838 278103 601840
rect 88977 601835 89043 601838
rect 229645 601835 229711 601838
rect 278037 601835 278103 601838
rect 211613 601762 211679 601765
rect 582741 601762 582807 601765
rect 211613 601760 582807 601762
rect 211613 601704 211618 601760
rect 211674 601704 582746 601760
rect 582802 601704 582807 601760
rect 211613 601702 582807 601704
rect 211613 601699 211679 601702
rect 582741 601699 582807 601702
rect 211654 600748 211660 600812
rect 211724 600810 211730 600812
rect 219525 600810 219591 600813
rect 211724 600808 219591 600810
rect 211724 600752 219530 600808
rect 219586 600752 219591 600808
rect 211724 600750 219591 600752
rect 211724 600748 211730 600750
rect 219525 600747 219591 600750
rect 221365 600810 221431 600813
rect 246246 600810 246252 600812
rect 221365 600808 246252 600810
rect 221365 600752 221370 600808
rect 221426 600752 246252 600808
rect 221365 600750 246252 600752
rect 221365 600747 221431 600750
rect 246246 600748 246252 600750
rect 246316 600748 246322 600812
rect 186957 600674 187023 600677
rect 222285 600674 222351 600677
rect 222653 600674 222719 600677
rect 186957 600672 222719 600674
rect 186957 600616 186962 600672
rect 187018 600616 222290 600672
rect 222346 600616 222658 600672
rect 222714 600616 222719 600672
rect 186957 600614 222719 600616
rect 186957 600611 187023 600614
rect 222285 600611 222351 600614
rect 222653 600611 222719 600614
rect 243629 600674 243695 600677
rect 258390 600674 258396 600676
rect 243629 600672 258396 600674
rect 243629 600616 243634 600672
rect 243690 600616 258396 600672
rect 243629 600614 258396 600616
rect 243629 600611 243695 600614
rect 258390 600612 258396 600614
rect 258460 600612 258466 600676
rect 165521 600538 165587 600541
rect 198549 600538 198615 600541
rect 165521 600536 198615 600538
rect 165521 600480 165526 600536
rect 165582 600480 198554 600536
rect 198610 600480 198615 600536
rect 165521 600478 198615 600480
rect 165521 600475 165587 600478
rect 198549 600475 198615 600478
rect 209957 600538 210023 600541
rect 219934 600538 219940 600540
rect 209957 600536 219940 600538
rect 209957 600480 209962 600536
rect 210018 600480 219940 600536
rect 209957 600478 219940 600480
rect 209957 600475 210023 600478
rect 219934 600476 219940 600478
rect 220004 600476 220010 600540
rect 229686 600476 229692 600540
rect 229756 600538 229762 600540
rect 237557 600538 237623 600541
rect 229756 600536 237623 600538
rect 229756 600480 237562 600536
rect 237618 600480 237623 600536
rect 229756 600478 237623 600480
rect 229756 600476 229762 600478
rect 237557 600475 237623 600478
rect 237966 600476 237972 600540
rect 238036 600538 238042 600540
rect 244181 600538 244247 600541
rect 238036 600536 244247 600538
rect 238036 600480 244186 600536
rect 244242 600480 244247 600536
rect 238036 600478 244247 600480
rect 238036 600476 238042 600478
rect 244181 600475 244247 600478
rect 248781 600538 248847 600541
rect 253381 600538 253447 600541
rect 248781 600536 253447 600538
rect 248781 600480 248786 600536
rect 248842 600480 253386 600536
rect 253442 600480 253447 600536
rect 248781 600478 253447 600480
rect 248781 600475 248847 600478
rect 253381 600475 253447 600478
rect 192334 600340 192340 600404
rect 192404 600402 192410 600404
rect 194685 600402 194751 600405
rect 192404 600400 194751 600402
rect 192404 600344 194690 600400
rect 194746 600344 194751 600400
rect 192404 600342 194751 600344
rect 192404 600340 192410 600342
rect 194685 600339 194751 600342
rect 197353 600402 197419 600405
rect 201677 600402 201743 600405
rect 215293 600404 215359 600405
rect 215293 600402 215340 600404
rect 197353 600400 201743 600402
rect 197353 600344 197358 600400
rect 197414 600344 201682 600400
rect 201738 600344 201743 600400
rect 197353 600342 201743 600344
rect 215212 600400 215340 600402
rect 215404 600402 215410 600404
rect 216397 600402 216463 600405
rect 215404 600400 216463 600402
rect 215212 600344 215298 600400
rect 215404 600344 216402 600400
rect 216458 600344 216463 600400
rect 215212 600342 215340 600344
rect 197353 600339 197419 600342
rect 201677 600339 201743 600342
rect 215293 600340 215340 600342
rect 215404 600342 216463 600344
rect 215404 600340 215410 600342
rect 215293 600339 215359 600340
rect 216397 600339 216463 600342
rect 226926 600340 226932 600404
rect 226996 600402 227002 600404
rect 231485 600402 231551 600405
rect 226996 600400 231551 600402
rect 226996 600344 231490 600400
rect 231546 600344 231551 600400
rect 226996 600342 231551 600344
rect 226996 600340 227002 600342
rect 231485 600339 231551 600342
rect 236637 600402 236703 600405
rect 239254 600402 239260 600404
rect 236637 600400 239260 600402
rect 236637 600344 236642 600400
rect 236698 600344 239260 600400
rect 236637 600342 239260 600344
rect 236637 600339 236703 600342
rect 239254 600340 239260 600342
rect 239324 600340 239330 600404
rect 250069 600402 250135 600405
rect 253473 600402 253539 600405
rect 250069 600400 253539 600402
rect 250069 600344 250074 600400
rect 250130 600344 253478 600400
rect 253534 600344 253539 600400
rect 250069 600342 253539 600344
rect 250069 600339 250135 600342
rect 253473 600339 253539 600342
rect 187601 599586 187667 599589
rect 218237 599586 218303 599589
rect 187601 599584 218303 599586
rect 187601 599528 187606 599584
rect 187662 599528 218242 599584
rect 218298 599528 218303 599584
rect 187601 599526 218303 599528
rect 187601 599523 187667 599526
rect 218237 599523 218303 599526
rect 79317 599450 79383 599453
rect 248413 599450 248479 599453
rect 79317 599448 248479 599450
rect 79317 599392 79322 599448
rect 79378 599392 248418 599448
rect 248474 599392 248479 599448
rect 79317 599390 248479 599392
rect 79317 599387 79383 599390
rect 248370 599387 248479 599390
rect 192753 599314 192819 599317
rect 212533 599314 212599 599317
rect 192753 599312 212599 599314
rect 192753 599256 192758 599312
rect 192814 599256 212538 599312
rect 212594 599256 212599 599312
rect 192753 599254 212599 599256
rect 248370 599314 248430 599387
rect 249333 599314 249399 599317
rect 253565 599314 253631 599317
rect 248370 599312 253631 599314
rect 248370 599256 249338 599312
rect 249394 599256 253570 599312
rect 253626 599256 253631 599312
rect 248370 599254 253631 599256
rect 192753 599251 192819 599254
rect 212533 599251 212599 599254
rect 249333 599251 249399 599254
rect 253565 599251 253631 599254
rect 213361 599178 213427 599181
rect 222694 599178 222700 599180
rect 213361 599176 222700 599178
rect 213361 599120 213366 599176
rect 213422 599120 222700 599176
rect 213361 599118 222700 599120
rect 213361 599115 213427 599118
rect 222694 599116 222700 599118
rect 222764 599116 222770 599180
rect 223798 599116 223804 599180
rect 223868 599178 223874 599180
rect 224217 599178 224283 599181
rect 223868 599176 224283 599178
rect 223868 599120 224222 599176
rect 224278 599120 224283 599176
rect 223868 599118 224283 599120
rect 223868 599116 223874 599118
rect 224217 599115 224283 599118
rect 228633 599178 228699 599181
rect 276013 599178 276079 599181
rect 228633 599176 276079 599178
rect 228633 599120 228638 599176
rect 228694 599120 276018 599176
rect 276074 599120 276079 599176
rect 228633 599118 276079 599120
rect 228633 599115 228699 599118
rect 276013 599115 276079 599118
rect 191097 599042 191163 599045
rect 193630 599042 193690 599080
rect 197169 599044 197235 599045
rect 197118 599042 197124 599044
rect 191097 599040 193690 599042
rect 191097 598984 191102 599040
rect 191158 598984 193690 599040
rect 191097 598982 193690 598984
rect 197078 598982 197124 599042
rect 197188 599040 197235 599044
rect 197230 598984 197235 599040
rect 191097 598979 191163 598982
rect 197118 598980 197124 598982
rect 197188 598980 197235 598984
rect 197169 598979 197235 598980
rect 202597 599042 202663 599045
rect 207105 599044 207171 599045
rect 210417 599044 210483 599045
rect 203190 599042 203196 599044
rect 202597 599040 203196 599042
rect 202597 598984 202602 599040
rect 202658 598984 203196 599040
rect 202597 598982 203196 598984
rect 202597 598979 202663 598982
rect 203190 598980 203196 598982
rect 203260 598980 203266 599044
rect 207054 599042 207060 599044
rect 207014 598982 207060 599042
rect 207124 599040 207171 599044
rect 210366 599042 210372 599044
rect 207166 598984 207171 599040
rect 207054 598980 207060 598982
rect 207124 598980 207171 598984
rect 210326 598982 210372 599042
rect 210436 599040 210483 599044
rect 210478 598984 210483 599040
rect 210366 598980 210372 598982
rect 210436 598980 210483 598984
rect 207105 598979 207171 598980
rect 210417 598979 210483 598980
rect 214005 599042 214071 599045
rect 216673 599044 216739 599045
rect 218697 599044 218763 599045
rect 220905 599044 220971 599045
rect 224033 599044 224099 599045
rect 216438 599042 216444 599044
rect 214005 599040 216444 599042
rect 214005 598984 214010 599040
rect 214066 598984 216444 599040
rect 214005 598982 216444 598984
rect 214005 598979 214071 598982
rect 216438 598980 216444 598982
rect 216508 598980 216514 599044
rect 216622 598980 216628 599044
rect 216692 599042 216739 599044
rect 218646 599042 218652 599044
rect 216692 599040 216784 599042
rect 216734 598984 216784 599040
rect 216692 598982 216784 598984
rect 218606 598982 218652 599042
rect 218716 599040 218763 599044
rect 220854 599042 220860 599044
rect 218758 598984 218763 599040
rect 216692 598980 216739 598982
rect 218646 598980 218652 598982
rect 218716 598980 218763 598984
rect 220814 598982 220860 599042
rect 220924 599040 220971 599044
rect 223982 599042 223988 599044
rect 220966 598984 220971 599040
rect 220854 598980 220860 598982
rect 220924 598980 220971 598984
rect 223942 598982 223988 599042
rect 224052 599040 224099 599044
rect 224094 598984 224099 599040
rect 223982 598980 223988 598982
rect 224052 598980 224099 598984
rect 216673 598979 216739 598980
rect 218697 598979 218763 598980
rect 220905 598979 220971 598980
rect 224033 598979 224099 598980
rect 226057 599042 226123 599045
rect 226190 599042 226196 599044
rect 226057 599040 226196 599042
rect 226057 598984 226062 599040
rect 226118 598984 226196 599040
rect 226057 598982 226196 598984
rect 226057 598979 226123 598982
rect 226190 598980 226196 598982
rect 226260 598980 226266 599044
rect 226374 598980 226380 599044
rect 226444 599042 226450 599044
rect 226793 599042 226859 599045
rect 226444 599040 226859 599042
rect 226444 598984 226798 599040
rect 226854 598984 226859 599040
rect 226444 598982 226859 598984
rect 226444 598980 226450 598982
rect 226793 598979 226859 598982
rect 228214 598980 228220 599044
rect 228284 599042 228290 599044
rect 230013 599042 230079 599045
rect 228284 599040 230079 599042
rect 228284 598984 230018 599040
rect 230074 598984 230079 599040
rect 228284 598982 230079 598984
rect 228284 598980 228290 598982
rect 230013 598979 230079 598982
rect 232405 599042 232471 599045
rect 233233 599044 233299 599045
rect 234705 599044 234771 599045
rect 232998 599042 233004 599044
rect 232405 599040 233004 599042
rect 232405 598984 232410 599040
rect 232466 598984 233004 599040
rect 232405 598982 233004 598984
rect 232405 598979 232471 598982
rect 232998 598980 233004 598982
rect 233068 598980 233074 599044
rect 233182 599042 233188 599044
rect 233142 598982 233188 599042
rect 233252 599040 233299 599044
rect 234654 599042 234660 599044
rect 233294 598984 233299 599040
rect 233182 598980 233188 598982
rect 233252 598980 233299 598984
rect 234614 598982 234660 599042
rect 234724 599040 234771 599044
rect 234766 598984 234771 599040
rect 234654 598980 234660 598982
rect 234724 598980 234771 598984
rect 236494 598980 236500 599044
rect 236564 599042 236570 599044
rect 236821 599042 236887 599045
rect 236564 599040 236887 599042
rect 236564 598984 236826 599040
rect 236882 598984 236887 599040
rect 236564 598982 236887 598984
rect 236564 598980 236570 598982
rect 233233 598979 233299 598980
rect 234705 598979 234771 598980
rect 236821 598979 236887 598982
rect 240685 599044 240751 599045
rect 247769 599044 247835 599045
rect 240685 599040 240732 599044
rect 240796 599042 240802 599044
rect 247718 599042 247724 599044
rect 240685 598984 240690 599040
rect 240685 598980 240732 598984
rect 240796 598982 240842 599042
rect 247678 598982 247724 599042
rect 247788 599040 247835 599044
rect 247830 598984 247835 599040
rect 240796 598980 240802 598982
rect 247718 598980 247724 598982
rect 247788 598980 247835 598984
rect 240685 598979 240751 598980
rect 247769 598979 247835 598980
rect 250897 599042 250963 599045
rect 251030 599042 251036 599044
rect 250897 599040 251036 599042
rect 250897 598984 250902 599040
rect 250958 598984 251036 599040
rect 250897 598982 251036 598984
rect 250897 598979 250963 598982
rect 251030 598980 251036 598982
rect 251100 598980 251106 599044
rect 252502 598980 252508 599044
rect 252572 599042 252578 599044
rect 252829 599042 252895 599045
rect 252572 599040 252895 599042
rect 252572 598984 252834 599040
rect 252890 598984 252895 599040
rect 252572 598982 252895 598984
rect 252572 598980 252578 598982
rect 252829 598979 252895 598982
rect 253565 599042 253631 599045
rect 262213 599042 262279 599045
rect 253565 599040 262279 599042
rect 253565 598984 253570 599040
rect 253626 598984 262218 599040
rect 262274 598984 262279 599040
rect 253565 598982 262279 598984
rect 253565 598979 253631 598982
rect 262213 598979 262279 598982
rect 191741 598906 191807 598909
rect 255957 598906 256023 598909
rect 191741 598904 193690 598906
rect 191741 598848 191746 598904
rect 191802 598848 193690 598904
rect 191741 598846 193690 598848
rect 191741 598843 191807 598846
rect 193254 598436 193260 598500
rect 193324 598498 193330 598500
rect 193489 598498 193555 598501
rect 193324 598496 193555 598498
rect 193324 598440 193494 598496
rect 193550 598440 193555 598496
rect 193324 598438 193555 598440
rect 193324 598436 193330 598438
rect 193489 598435 193555 598438
rect 193630 598264 193690 598846
rect 253430 598904 256023 598906
rect 253430 598848 255962 598904
rect 256018 598848 256023 598904
rect 253430 598846 256023 598848
rect 253430 598808 253490 598846
rect 255957 598843 256023 598846
rect 184197 597818 184263 597821
rect 193305 597818 193371 597821
rect 184197 597816 193371 597818
rect 184197 597760 184202 597816
rect 184258 597760 193310 597816
rect 193366 597760 193371 597816
rect 184197 597758 193371 597760
rect 184197 597755 184263 597758
rect 193305 597755 193371 597758
rect 253430 597682 253490 597720
rect 255405 597682 255471 597685
rect 253430 597680 255471 597682
rect 253430 597624 255410 597680
rect 255466 597624 255471 597680
rect 253430 597622 255471 597624
rect 255405 597619 255471 597622
rect 170990 596804 170996 596868
rect 171060 596866 171066 596868
rect 191649 596866 191715 596869
rect 193630 596866 193690 597176
rect 171060 596864 193690 596866
rect 171060 596808 191654 596864
rect 191710 596808 193690 596864
rect 171060 596806 193690 596808
rect 171060 596804 171066 596806
rect 191649 596803 191715 596806
rect 253430 596594 253490 596904
rect 255405 596594 255471 596597
rect 253430 596592 255471 596594
rect 253430 596536 255410 596592
rect 255466 596536 255471 596592
rect 253430 596534 255471 596536
rect 255405 596531 255471 596534
rect 190637 596322 190703 596325
rect 193630 596322 193690 596360
rect 190637 596320 193690 596322
rect 190637 596264 190642 596320
rect 190698 596264 193690 596320
rect 190637 596262 193690 596264
rect 190637 596259 190703 596262
rect 190637 595234 190703 595237
rect 193630 595234 193690 595544
rect 190637 595232 193690 595234
rect 190637 595176 190642 595232
rect 190698 595176 193690 595232
rect 190637 595174 193690 595176
rect 253430 595234 253490 595816
rect 254526 595234 254532 595236
rect 253430 595174 254532 595234
rect 190637 595171 190703 595174
rect 254526 595172 254532 595174
rect 254596 595172 254602 595236
rect 253430 594962 253490 595000
rect 266302 594962 266308 594964
rect 253430 594902 266308 594962
rect 266302 594900 266308 594902
rect 266372 594900 266378 594964
rect 191741 594690 191807 594693
rect 191741 594688 193690 594690
rect 191741 594632 191746 594688
rect 191802 594632 193690 594688
rect 191741 594630 193690 594632
rect 191741 594627 191807 594630
rect 193630 594456 193690 594630
rect 255313 594282 255379 594285
rect 253430 594280 255379 594282
rect 253430 594224 255318 594280
rect 255374 594224 255379 594280
rect 253430 594222 255379 594224
rect 253430 594184 253490 594222
rect 255313 594219 255379 594222
rect 191649 593466 191715 593469
rect 193630 593466 193690 593640
rect 191649 593464 193690 593466
rect 191649 593408 191654 593464
rect 191710 593408 193690 593464
rect 191649 593406 193690 593408
rect 191649 593403 191715 593406
rect -960 592908 480 593148
rect 179270 592724 179276 592788
rect 179340 592786 179346 592788
rect 193397 592786 193463 592789
rect 179340 592784 193463 592786
rect 179340 592728 193402 592784
rect 193458 592728 193463 592784
rect 179340 592726 193463 592728
rect 253430 592786 253490 593096
rect 256325 592786 256391 592789
rect 253430 592784 256391 592786
rect 253430 592728 256330 592784
rect 256386 592728 256391 592784
rect 253430 592726 256391 592728
rect 179340 592724 179346 592726
rect 193397 592723 193463 592726
rect 256325 592723 256391 592726
rect 191741 592378 191807 592381
rect 193630 592378 193690 592552
rect 191741 592376 193690 592378
rect 191741 592320 191746 592376
rect 191802 592320 193690 592376
rect 191741 592318 193690 592320
rect 191741 592315 191807 592318
rect 253430 592109 253490 592280
rect 253381 592104 253490 592109
rect 253381 592048 253386 592104
rect 253442 592048 253490 592104
rect 253381 592046 253490 592048
rect 253381 592043 253447 592046
rect 191005 591290 191071 591293
rect 193630 591290 193690 591736
rect 191005 591288 193690 591290
rect 191005 591232 191010 591288
rect 191066 591232 193690 591288
rect 191005 591230 193690 591232
rect 191005 591227 191071 591230
rect 253430 591018 253490 591192
rect 255405 591018 255471 591021
rect 253430 591016 255471 591018
rect 253430 590960 255410 591016
rect 255466 590960 255471 591016
rect 253430 590958 255471 590960
rect 255405 590955 255471 590958
rect 582373 591018 582439 591021
rect 583520 591018 584960 591108
rect 582373 591016 584960 591018
rect 582373 590960 582378 591016
rect 582434 590960 584960 591016
rect 582373 590958 584960 590960
rect 582373 590955 582439 590958
rect 583520 590868 584960 590958
rect 191598 590684 191604 590748
rect 191668 590746 191674 590748
rect 191668 590686 193690 590746
rect 191668 590684 191674 590686
rect 193630 590648 193690 590686
rect 172329 589930 172395 589933
rect 193254 589930 193260 589932
rect 172329 589928 193260 589930
rect 172329 589872 172334 589928
rect 172390 589872 193260 589928
rect 172329 589870 193260 589872
rect 172329 589867 172395 589870
rect 193254 589868 193260 589870
rect 193324 589868 193330 589932
rect 253430 589930 253490 590376
rect 255405 589930 255471 589933
rect 253430 589928 255471 589930
rect 253430 589872 255410 589928
rect 255466 589872 255471 589928
rect 253430 589870 255471 589872
rect 255405 589867 255471 589870
rect 191281 589386 191347 589389
rect 193630 589386 193690 589832
rect 262254 589386 262260 589388
rect 191281 589384 193690 589386
rect 191281 589328 191286 589384
rect 191342 589328 193690 589384
rect 191281 589326 193690 589328
rect 253430 589326 262260 589386
rect 191281 589323 191347 589326
rect 253430 589288 253490 589326
rect 262254 589324 262260 589326
rect 262324 589324 262330 589388
rect 168230 588100 168236 588164
rect 168300 588162 168306 588164
rect 193630 588162 193690 588744
rect 168300 588102 193690 588162
rect 253430 588162 253490 588472
rect 255405 588162 255471 588165
rect 253430 588160 255471 588162
rect 253430 588104 255410 588160
rect 255466 588104 255471 588160
rect 253430 588102 255471 588104
rect 168300 588100 168306 588102
rect 255405 588099 255471 588102
rect 162710 587964 162716 588028
rect 162780 588026 162786 588028
rect 162780 587966 193690 588026
rect 162780 587964 162786 587966
rect 193630 587928 193690 587966
rect 253933 587414 253999 587417
rect 253460 587412 253999 587414
rect 253460 587356 253938 587412
rect 253994 587356 253999 587412
rect 253460 587354 253999 587356
rect 253933 587351 253999 587354
rect 190453 586530 190519 586533
rect 190453 586528 190562 586530
rect 190453 586472 190458 586528
rect 190514 586472 190562 586528
rect 190453 586467 190562 586472
rect 190502 586394 190562 586467
rect 193630 586394 193690 587112
rect 190502 586334 193690 586394
rect 253430 586394 253490 586568
rect 256734 586468 256740 586532
rect 256804 586468 256810 586532
rect 256742 586394 256802 586468
rect 253430 586334 256802 586394
rect 191189 586258 191255 586261
rect 191189 586256 193690 586258
rect 191189 586200 191194 586256
rect 191250 586200 193690 586256
rect 191189 586198 193690 586200
rect 191189 586195 191255 586198
rect 193630 586024 193690 586198
rect 191741 585170 191807 585173
rect 193630 585170 193690 585208
rect 191741 585168 193690 585170
rect 191741 585112 191746 585168
rect 191802 585112 193690 585168
rect 191741 585110 193690 585112
rect 253430 585170 253490 585480
rect 255405 585170 255471 585173
rect 253430 585168 255471 585170
rect 253430 585112 255410 585168
rect 255466 585112 255471 585168
rect 253430 585110 255471 585112
rect 191741 585107 191807 585110
rect 255405 585107 255471 585110
rect 118693 585034 118759 585037
rect 119337 585034 119403 585037
rect 188337 585034 188403 585037
rect 118693 585032 188403 585034
rect 118693 584976 118698 585032
rect 118754 584976 119342 585032
rect 119398 584976 188342 585032
rect 188398 584976 188403 585032
rect 118693 584974 188403 584976
rect 118693 584971 118759 584974
rect 119337 584971 119403 584974
rect 188337 584971 188403 584974
rect 253430 584354 253490 584664
rect 253430 584294 258090 584354
rect 255313 584218 255379 584221
rect 253430 584216 255379 584218
rect 253430 584160 255318 584216
rect 255374 584160 255379 584216
rect 253430 584158 255379 584160
rect 191741 583946 191807 583949
rect 193630 583946 193690 584120
rect 191741 583944 193690 583946
rect 191741 583888 191746 583944
rect 191802 583888 193690 583944
rect 191741 583886 193690 583888
rect 191741 583883 191807 583886
rect 253430 583848 253490 584158
rect 255313 584155 255379 584158
rect 258030 584082 258090 584294
rect 280286 584082 280292 584084
rect 258030 584022 280292 584082
rect 280286 584020 280292 584022
rect 280356 584020 280362 584084
rect 82721 582722 82787 582725
rect 122097 582722 122163 582725
rect 82721 582720 122163 582722
rect 82721 582664 82726 582720
rect 82782 582664 122102 582720
rect 122158 582664 122163 582720
rect 82721 582662 122163 582664
rect 82721 582659 82787 582662
rect 122097 582659 122163 582662
rect 191741 582722 191807 582725
rect 193630 582722 193690 583304
rect 255405 583266 255471 583269
rect 253430 583264 255471 583266
rect 253430 583208 255410 583264
rect 255466 583208 255471 583264
rect 253430 583206 255471 583208
rect 253430 582760 253490 583206
rect 255405 583203 255471 583206
rect 191741 582720 193690 582722
rect 191741 582664 191746 582720
rect 191802 582664 193690 582720
rect 191741 582662 193690 582664
rect 191741 582659 191807 582662
rect 55029 582586 55095 582589
rect 82997 582586 83063 582589
rect 55029 582584 83063 582586
rect 55029 582528 55034 582584
rect 55090 582528 83002 582584
rect 83058 582528 83063 582584
rect 55029 582526 83063 582528
rect 55029 582523 55095 582526
rect 82997 582523 83063 582526
rect 254025 582314 254091 582317
rect 253430 582312 254091 582314
rect 253430 582256 254030 582312
rect 254086 582256 254091 582312
rect 253430 582254 254091 582256
rect 191741 581634 191807 581637
rect 193630 581634 193690 582216
rect 253430 581944 253490 582254
rect 254025 582251 254091 582254
rect 191741 581632 193690 581634
rect 191741 581576 191746 581632
rect 191802 581576 193690 581632
rect 191741 581574 193690 581576
rect 191741 581571 191807 581574
rect 74257 581226 74323 581229
rect 79961 581228 80027 581229
rect 79910 581226 79916 581228
rect 74257 581224 79426 581226
rect 74257 581168 74262 581224
rect 74318 581168 79426 581224
rect 74257 581166 79426 581168
rect 79834 581166 79916 581226
rect 79980 581226 80027 581228
rect 98545 581226 98611 581229
rect 79980 581224 98611 581226
rect 80022 581168 98550 581224
rect 98606 581168 98611 581224
rect 74257 581163 74323 581166
rect 75361 581090 75427 581093
rect 75678 581090 75684 581092
rect 75361 581088 75684 581090
rect 75361 581032 75366 581088
rect 75422 581032 75684 581088
rect 75361 581030 75684 581032
rect 75361 581027 75427 581030
rect 75678 581028 75684 581030
rect 75748 581028 75754 581092
rect 79366 581090 79426 581166
rect 79910 581164 79916 581166
rect 79980 581166 98611 581168
rect 79980 581164 80027 581166
rect 79961 581163 80027 581164
rect 98545 581163 98611 581166
rect 105537 581090 105603 581093
rect 79366 581088 105603 581090
rect 79366 581032 105542 581088
rect 105598 581032 105603 581088
rect 79366 581030 105603 581032
rect 105537 581027 105603 581030
rect 173157 581090 173223 581093
rect 193630 581090 193690 581400
rect 173157 581088 193690 581090
rect 173157 581032 173162 581088
rect 173218 581032 193690 581088
rect 173157 581030 193690 581032
rect 173157 581027 173223 581030
rect 71497 580818 71563 580821
rect 71630 580818 71636 580820
rect 71497 580816 71636 580818
rect 71497 580760 71502 580816
rect 71558 580760 71636 580816
rect 71497 580758 71636 580760
rect 71497 580755 71563 580758
rect 71630 580756 71636 580758
rect 71700 580756 71706 580820
rect 80881 580818 80947 580821
rect 81014 580818 81020 580820
rect 80881 580816 81020 580818
rect 80881 580760 80886 580816
rect 80942 580760 81020 580816
rect 80881 580758 81020 580760
rect 80881 580755 80947 580758
rect 81014 580756 81020 580758
rect 81084 580756 81090 580820
rect 83958 580756 83964 580820
rect 84028 580818 84034 580820
rect 84193 580818 84259 580821
rect 84028 580816 84259 580818
rect 84028 580760 84198 580816
rect 84254 580760 84259 580816
rect 84028 580758 84259 580760
rect 84028 580756 84034 580758
rect 84193 580755 84259 580758
rect 89253 580820 89319 580821
rect 89253 580816 89300 580820
rect 89364 580818 89370 580820
rect 89253 580760 89258 580816
rect 89253 580756 89300 580760
rect 89364 580758 89410 580818
rect 89364 580756 89370 580758
rect 89253 580755 89319 580756
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 66621 580002 66687 580005
rect 68878 580002 68938 580584
rect 66621 580000 68938 580002
rect 66621 579944 66626 580000
rect 66682 579944 68938 580000
rect 66621 579942 68938 579944
rect 66621 579939 66687 579942
rect 169109 579730 169175 579733
rect 193630 579730 193690 580312
rect 253430 580274 253490 580856
rect 263542 580274 263548 580276
rect 253430 580214 263548 580274
rect 263542 580212 263548 580214
rect 263612 580212 263618 580276
rect 169109 579728 193690 579730
rect 169109 579672 169114 579728
rect 169170 579672 193690 579728
rect 169109 579670 193690 579672
rect 253430 579730 253490 580040
rect 255405 579730 255471 579733
rect 253430 579728 255471 579730
rect 253430 579672 255410 579728
rect 255466 579672 255471 579728
rect 253430 579670 255471 579672
rect 169109 579667 169175 579670
rect 255405 579667 255471 579670
rect 66437 578642 66503 578645
rect 68878 578642 68938 579224
rect 94638 578914 94698 579496
rect 96797 578914 96863 578917
rect 94638 578912 96863 578914
rect 94638 578856 96802 578912
rect 96858 578856 96863 578912
rect 94638 578854 96863 578856
rect 96797 578851 96863 578854
rect 191741 578914 191807 578917
rect 193630 578914 193690 579496
rect 191741 578912 193690 578914
rect 191741 578856 191746 578912
rect 191802 578856 193690 578912
rect 191741 578854 193690 578856
rect 191741 578851 191807 578854
rect 66437 578640 68938 578642
rect 66437 578584 66442 578640
rect 66498 578584 68938 578640
rect 66437 578582 68938 578584
rect 66437 578579 66503 578582
rect 186221 578370 186287 578373
rect 191097 578370 191163 578373
rect 186221 578368 191163 578370
rect 186221 578312 186226 578368
rect 186282 578312 191102 578368
rect 191158 578312 191163 578368
rect 186221 578310 191163 578312
rect 186221 578307 186287 578310
rect 191097 578307 191163 578310
rect 191557 578370 191623 578373
rect 193630 578370 193690 578408
rect 191557 578368 193690 578370
rect 191557 578312 191562 578368
rect 191618 578312 193690 578368
rect 191557 578310 193690 578312
rect 253430 578370 253490 578952
rect 267774 578370 267780 578372
rect 253430 578310 267780 578370
rect 191557 578307 191623 578310
rect 267774 578308 267780 578310
rect 267844 578308 267850 578372
rect 67173 577418 67239 577421
rect 68878 577418 68938 577864
rect 94638 577554 94698 578136
rect 191741 578098 191807 578101
rect 191741 578096 193690 578098
rect 191741 578040 191746 578096
rect 191802 578040 193690 578096
rect 191741 578038 193690 578040
rect 191741 578035 191807 578038
rect 193630 577592 193690 578038
rect 97901 577554 97967 577557
rect 94638 577552 97967 577554
rect 94638 577496 97906 577552
rect 97962 577496 97967 577552
rect 94638 577494 97967 577496
rect 253430 577554 253490 578136
rect 582373 577690 582439 577693
rect 583520 577690 584960 577780
rect 582373 577688 584960 577690
rect 582373 577632 582378 577688
rect 582434 577632 584960 577688
rect 582373 577630 584960 577632
rect 582373 577627 582439 577630
rect 254025 577554 254091 577557
rect 253430 577552 254091 577554
rect 253430 577496 254030 577552
rect 254086 577496 254091 577552
rect 583520 577540 584960 577630
rect 253430 577494 254091 577496
rect 97901 577491 97967 577494
rect 254025 577491 254091 577494
rect 67173 577416 68938 577418
rect 67173 577360 67178 577416
rect 67234 577360 68938 577416
rect 67173 577358 68938 577360
rect 67173 577355 67239 577358
rect 253430 577010 253490 577048
rect 255405 577010 255471 577013
rect 253430 577008 255471 577010
rect 253430 576952 255410 577008
rect 255466 576952 255471 577008
rect 253430 576950 255471 576952
rect 255405 576947 255471 576950
rect 94638 576738 94698 576776
rect 97901 576738 97967 576741
rect 94638 576736 97967 576738
rect 94638 576680 97906 576736
rect 97962 576680 97967 576736
rect 94638 576678 97967 576680
rect 97901 576675 97967 576678
rect 67541 576466 67607 576469
rect 68878 576466 68938 576504
rect 67541 576464 68938 576466
rect 67541 576408 67546 576464
rect 67602 576408 68938 576464
rect 67541 576406 68938 576408
rect 67541 576403 67607 576406
rect 191005 576194 191071 576197
rect 193630 576194 193690 576776
rect 191005 576192 193690 576194
rect 191005 576136 191010 576192
rect 191066 576136 193690 576192
rect 191005 576134 193690 576136
rect 191005 576131 191071 576134
rect 253430 575922 253490 576232
rect 255405 575922 255471 575925
rect 253430 575920 255471 575922
rect 253430 575864 255410 575920
rect 255466 575864 255471 575920
rect 253430 575862 255471 575864
rect 255405 575859 255471 575862
rect 191189 575650 191255 575653
rect 193630 575650 193690 575688
rect 191189 575648 193690 575650
rect 191189 575592 191194 575648
rect 191250 575592 193690 575648
rect 191189 575590 193690 575592
rect 191189 575587 191255 575590
rect 191598 575452 191604 575516
rect 191668 575514 191674 575516
rect 193438 575514 193444 575516
rect 191668 575454 193444 575514
rect 191668 575452 191674 575454
rect 193438 575452 193444 575454
rect 193508 575452 193514 575516
rect 67357 575378 67423 575381
rect 67357 575376 68938 575378
rect 67357 575320 67362 575376
rect 67418 575320 68938 575376
rect 67357 575318 68938 575320
rect 67357 575315 67423 575318
rect 68878 575144 68938 575318
rect 94638 574834 94698 575416
rect 96797 574834 96863 574837
rect 94638 574832 96863 574834
rect 94638 574776 96802 574832
rect 96858 574776 96863 574832
rect 94638 574774 96863 574776
rect 96797 574771 96863 574774
rect 191281 574562 191347 574565
rect 193630 574562 193690 574872
rect 253430 574698 253490 575144
rect 255405 574698 255471 574701
rect 253430 574696 255471 574698
rect 253430 574640 255410 574696
rect 255466 574640 255471 574696
rect 253430 574638 255471 574640
rect 255405 574635 255471 574638
rect 191281 574560 193690 574562
rect 191281 574504 191286 574560
rect 191342 574504 193690 574560
rect 191281 574502 193690 574504
rect 191281 574499 191347 574502
rect 253430 574154 253490 574328
rect 255589 574154 255655 574157
rect 253430 574152 255655 574154
rect 253430 574096 255594 574152
rect 255650 574096 255655 574152
rect 253430 574094 255655 574096
rect 255589 574091 255655 574094
rect 66621 573202 66687 573205
rect 68878 573202 68938 573784
rect 94638 573474 94698 574056
rect 96889 573474 96955 573477
rect 94638 573472 96955 573474
rect 94638 573416 96894 573472
rect 96950 573416 96955 573472
rect 94638 573414 96955 573416
rect 96889 573411 96955 573414
rect 191005 573338 191071 573341
rect 193630 573338 193690 573784
rect 191005 573336 193690 573338
rect 191005 573280 191010 573336
rect 191066 573280 193690 573336
rect 191005 573278 193690 573280
rect 191005 573275 191071 573278
rect 66621 573200 68938 573202
rect 66621 573144 66626 573200
rect 66682 573144 68938 573200
rect 66621 573142 68938 573144
rect 66621 573139 66687 573142
rect 191557 572794 191623 572797
rect 193630 572794 193690 572968
rect 253430 572930 253490 573512
rect 255497 572930 255563 572933
rect 253430 572928 255563 572930
rect 253430 572872 255502 572928
rect 255558 572872 255563 572928
rect 253430 572870 255563 572872
rect 255497 572867 255563 572870
rect 191557 572792 193690 572794
rect 191557 572736 191562 572792
rect 191618 572736 193690 572792
rect 191557 572734 193690 572736
rect 191557 572731 191623 572734
rect 94638 572658 94698 572696
rect 97901 572658 97967 572661
rect 255405 572658 255471 572661
rect 94638 572656 97967 572658
rect 94638 572600 97906 572656
rect 97962 572600 97967 572656
rect 94638 572598 97967 572600
rect 97901 572595 97967 572598
rect 253430 572656 255471 572658
rect 253430 572600 255410 572656
rect 255466 572600 255471 572656
rect 253430 572598 255471 572600
rect 253430 572424 253490 572598
rect 255405 572595 255471 572598
rect 66621 571842 66687 571845
rect 68878 571842 68938 572424
rect 191281 572250 191347 572253
rect 191281 572248 193690 572250
rect 191281 572192 191286 572248
rect 191342 572192 193690 572248
rect 191281 572190 193690 572192
rect 191281 572187 191347 572190
rect 193630 571880 193690 572190
rect 66621 571840 68938 571842
rect 66621 571784 66626 571840
rect 66682 571784 68938 571840
rect 66621 571782 68938 571784
rect 66621 571779 66687 571782
rect 253430 571570 253490 571608
rect 255405 571570 255471 571573
rect 253430 571568 255471 571570
rect 253430 571512 255410 571568
rect 255466 571512 255471 571568
rect 253430 571510 255471 571512
rect 255405 571507 255471 571510
rect 97717 571434 97783 571437
rect 94638 571432 97783 571434
rect 94638 571376 97722 571432
rect 97778 571376 97783 571432
rect 94638 571374 97783 571376
rect 94638 571336 94698 571374
rect 97717 571371 97783 571374
rect 191557 570890 191623 570893
rect 193630 570890 193690 571064
rect 191557 570888 193690 570890
rect 191557 570832 191562 570888
rect 191618 570832 193690 570888
rect 191557 570830 193690 570832
rect 191557 570827 191623 570830
rect 66621 570210 66687 570213
rect 68878 570210 68938 570792
rect 192334 570754 192340 570756
rect 180750 570694 192340 570754
rect 153929 570618 153995 570621
rect 180750 570618 180810 570694
rect 192334 570692 192340 570694
rect 192404 570692 192410 570756
rect 153929 570616 180810 570618
rect 153929 570560 153934 570616
rect 153990 570560 180810 570616
rect 153929 570558 180810 570560
rect 190913 570618 190979 570621
rect 255405 570618 255471 570621
rect 190913 570616 193690 570618
rect 190913 570560 190918 570616
rect 190974 570560 193690 570616
rect 190913 570558 193690 570560
rect 153929 570555 153995 570558
rect 190913 570555 190979 570558
rect 66621 570208 68938 570210
rect 66621 570152 66626 570208
rect 66682 570152 68938 570208
rect 66621 570150 68938 570152
rect 66621 570147 66687 570150
rect 97901 570074 97967 570077
rect 94638 570072 97967 570074
rect 94638 570016 97906 570072
rect 97962 570016 97967 570072
rect 94638 570014 97967 570016
rect 94638 569976 94698 570014
rect 97901 570011 97967 570014
rect 193630 569976 193690 570558
rect 253430 570616 255471 570618
rect 253430 570560 255410 570616
rect 255466 570560 255471 570616
rect 253430 570558 255471 570560
rect 253430 570520 253490 570558
rect 255405 570555 255471 570558
rect 67449 569938 67515 569941
rect 67449 569936 68938 569938
rect 67449 569880 67454 569936
rect 67510 569880 68938 569936
rect 67449 569878 68938 569880
rect 67449 569875 67515 569878
rect 68878 569432 68938 569878
rect 253430 569394 253490 569704
rect 255405 569394 255471 569397
rect 253430 569392 255471 569394
rect 253430 569336 255410 569392
rect 255466 569336 255471 569392
rect 253430 569334 255471 569336
rect 255405 569331 255471 569334
rect 96705 569122 96771 569125
rect 97441 569122 97507 569125
rect 94638 569120 97507 569122
rect 94638 569064 96710 569120
rect 96766 569064 97446 569120
rect 97502 569064 97507 569120
rect 94638 569062 97507 569064
rect 94638 568616 94698 569062
rect 96705 569059 96771 569062
rect 97441 569059 97507 569062
rect 190361 568714 190427 568717
rect 193630 568714 193690 569160
rect 255405 568714 255471 568717
rect 190361 568712 193690 568714
rect 190361 568656 190366 568712
rect 190422 568656 193690 568712
rect 190361 568654 193690 568656
rect 253430 568712 255471 568714
rect 253430 568656 255410 568712
rect 255466 568656 255471 568712
rect 253430 568654 255471 568656
rect 190361 568651 190427 568654
rect 253430 568616 253490 568654
rect 255405 568651 255471 568654
rect 67449 567626 67515 567629
rect 68878 567626 68938 568072
rect 96797 567898 96863 567901
rect 67449 567624 68938 567626
rect 67449 567568 67454 567624
rect 67510 567568 68938 567624
rect 67449 567566 68938 567568
rect 94638 567896 96863 567898
rect 94638 567840 96802 567896
rect 96858 567840 96863 567896
rect 94638 567838 96863 567840
rect 67449 567563 67515 567566
rect 94638 567256 94698 567838
rect 96797 567835 96863 567838
rect 190453 567626 190519 567629
rect 193630 567626 193690 568072
rect 190453 567624 193690 567626
rect 190453 567568 190458 567624
rect 190514 567568 193690 567624
rect 190453 567566 193690 567568
rect 253430 567626 253490 567800
rect 255773 567626 255839 567629
rect 253430 567624 255839 567626
rect 253430 567568 255778 567624
rect 255834 567568 255839 567624
rect 253430 567566 255839 567568
rect 190453 567563 190519 567566
rect 255773 567563 255839 567566
rect 191741 567218 191807 567221
rect 193630 567218 193690 567256
rect 191741 567216 193690 567218
rect 191741 567160 191746 567216
rect 191802 567160 193690 567216
rect 191741 567158 193690 567160
rect 191741 567155 191807 567158
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67633 566674 67699 566677
rect 68878 566674 68938 566712
rect 67633 566672 68938 566674
rect 67633 566616 67638 566672
rect 67694 566616 68938 566672
rect 67633 566614 68938 566616
rect 67633 566611 67699 566614
rect 94638 565858 94698 565896
rect 95417 565858 95483 565861
rect 94638 565856 95483 565858
rect 94638 565800 95422 565856
rect 95478 565800 95483 565856
rect 94638 565798 95483 565800
rect 95417 565795 95483 565798
rect 159950 565796 159956 565860
rect 160020 565858 160026 565860
rect 193630 565858 193690 566440
rect 253430 566402 253490 566712
rect 255681 566402 255747 566405
rect 253430 566400 255747 566402
rect 253430 566344 255686 566400
rect 255742 566344 255747 566400
rect 253430 566342 255747 566344
rect 255681 566339 255747 566342
rect 160020 565798 193690 565858
rect 253430 565858 253490 565896
rect 255589 565858 255655 565861
rect 253430 565856 255655 565858
rect 253430 565800 255594 565856
rect 255650 565800 255655 565856
rect 253430 565798 255655 565800
rect 160020 565796 160026 565798
rect 255589 565795 255655 565798
rect 66805 564770 66871 564773
rect 68878 564770 68938 565352
rect 158621 565042 158687 565045
rect 190453 565042 190519 565045
rect 158621 565040 190519 565042
rect 158621 564984 158626 565040
rect 158682 564984 190458 565040
rect 190514 564984 190519 565040
rect 158621 564982 190519 564984
rect 158621 564979 158687 564982
rect 190453 564979 190519 564982
rect 191097 564906 191163 564909
rect 193630 564906 193690 565352
rect 191097 564904 193690 564906
rect 191097 564848 191102 564904
rect 191158 564848 193690 564904
rect 191097 564846 193690 564848
rect 191097 564843 191163 564846
rect 66805 564768 68938 564770
rect 66805 564712 66810 564768
rect 66866 564712 68938 564768
rect 66805 564710 68938 564712
rect 190821 564770 190887 564773
rect 253430 564770 253490 565080
rect 255589 564770 255655 564773
rect 190821 564768 193690 564770
rect 190821 564712 190826 564768
rect 190882 564712 193690 564768
rect 190821 564710 193690 564712
rect 253430 564768 255655 564770
rect 253430 564712 255594 564768
rect 255650 564712 255655 564768
rect 253430 564710 255655 564712
rect 66805 564707 66871 564710
rect 190821 564707 190887 564710
rect 193630 564536 193690 564710
rect 255589 564707 255655 564710
rect 582833 564362 582899 564365
rect 583520 564362 584960 564452
rect 582833 564360 584960 564362
rect 582833 564304 582838 564360
rect 582894 564304 584960 564360
rect 582833 564302 584960 564304
rect 582833 564299 582899 564302
rect 66713 563410 66779 563413
rect 68878 563410 68938 563992
rect 94638 563682 94698 564264
rect 583520 564212 584960 564302
rect 95233 563682 95299 563685
rect 94638 563680 95299 563682
rect 94638 563624 95238 563680
rect 95294 563624 95299 563680
rect 94638 563622 95299 563624
rect 95233 563619 95299 563622
rect 191005 563682 191071 563685
rect 191005 563680 193690 563682
rect 191005 563624 191010 563680
rect 191066 563624 193690 563680
rect 191005 563622 193690 563624
rect 191005 563619 191071 563622
rect 193630 563448 193690 563622
rect 66713 563408 68938 563410
rect 66713 563352 66718 563408
rect 66774 563352 68938 563408
rect 66713 563350 68938 563352
rect 253430 563410 253490 563992
rect 267958 563410 267964 563412
rect 253430 563350 267964 563410
rect 66713 563347 66779 563350
rect 267958 563348 267964 563350
rect 268028 563348 268034 563412
rect 253430 563138 253490 563176
rect 255589 563138 255655 563141
rect 253430 563136 255655 563138
rect 253430 563080 255594 563136
rect 255650 563080 255655 563136
rect 253430 563078 255655 563080
rect 255589 563075 255655 563078
rect 67725 562050 67791 562053
rect 68878 562050 68938 562632
rect 94638 562322 94698 562904
rect 98085 562322 98151 562325
rect 94638 562320 98151 562322
rect 94638 562264 98090 562320
rect 98146 562264 98151 562320
rect 94638 562262 98151 562264
rect 98085 562259 98151 562262
rect 67725 562048 68938 562050
rect 67725 561992 67730 562048
rect 67786 561992 68938 562048
rect 67725 561990 68938 561992
rect 191741 562050 191807 562053
rect 193630 562050 193690 562632
rect 191741 562048 193690 562050
rect 191741 561992 191746 562048
rect 191802 561992 193690 562048
rect 191741 561990 193690 561992
rect 67725 561987 67791 561990
rect 191741 561987 191807 561990
rect 253430 561914 253490 562088
rect 255589 561914 255655 561917
rect 253430 561912 255655 561914
rect 253430 561856 255594 561912
rect 255650 561856 255655 561912
rect 253430 561854 255655 561856
rect 255589 561851 255655 561854
rect 66161 561642 66227 561645
rect 66161 561640 68938 561642
rect 66161 561584 66166 561640
rect 66222 561584 68938 561640
rect 66161 561582 68938 561584
rect 66161 561579 66227 561582
rect 68878 561272 68938 561582
rect 94638 561098 94698 561544
rect 96889 561098 96955 561101
rect 94638 561096 96955 561098
rect 94638 561040 96894 561096
rect 96950 561040 96955 561096
rect 94638 561038 96955 561040
rect 96889 561035 96955 561038
rect 191189 560962 191255 560965
rect 193630 560962 193690 561544
rect 191189 560960 193690 560962
rect 191189 560904 191194 560960
rect 191250 560904 193690 560960
rect 191189 560902 193690 560904
rect 191189 560899 191255 560902
rect 253430 560826 253490 561272
rect 255589 560826 255655 560829
rect 253430 560824 255655 560826
rect 253430 560768 255594 560824
rect 255650 560768 255655 560824
rect 253430 560766 255655 560768
rect 255589 560763 255655 560766
rect 191097 560690 191163 560693
rect 193630 560690 193690 560728
rect 191097 560688 193690 560690
rect 191097 560632 191102 560688
rect 191158 560632 193690 560688
rect 191097 560630 193690 560632
rect 191097 560627 191163 560630
rect 66805 559330 66871 559333
rect 68878 559330 68938 559912
rect 94638 559602 94698 560184
rect 96981 559602 97047 559605
rect 94638 559600 97047 559602
rect 94638 559544 96986 559600
rect 97042 559544 97047 559600
rect 94638 559542 97047 559544
rect 96981 559539 97047 559542
rect 66805 559328 68938 559330
rect 66805 559272 66810 559328
rect 66866 559272 68938 559328
rect 66805 559270 68938 559272
rect 66805 559267 66871 559270
rect 161238 558996 161244 559060
rect 161308 559058 161314 559060
rect 193630 559058 193690 559640
rect 253430 559602 253490 560184
rect 255589 559602 255655 559605
rect 253430 559600 255655 559602
rect 253430 559544 255594 559600
rect 255650 559544 255655 559600
rect 253430 559542 255655 559544
rect 255589 559539 255655 559542
rect 161308 558998 193690 559058
rect 253430 559058 253490 559368
rect 269062 559058 269068 559060
rect 253430 558998 269068 559058
rect 161308 558996 161314 558998
rect 269062 558996 269068 558998
rect 269132 558996 269138 559060
rect 95325 558922 95391 558925
rect 94638 558920 95391 558922
rect 94638 558864 95330 558920
rect 95386 558864 95391 558920
rect 94638 558862 95391 558864
rect 94638 558653 94698 558862
rect 95325 558859 95391 558862
rect 94638 558648 94747 558653
rect 94638 558592 94686 558648
rect 94742 558592 94747 558648
rect 94638 558590 94747 558592
rect 94681 558587 94747 558590
rect 66161 558106 66227 558109
rect 68878 558106 68938 558552
rect 190913 558242 190979 558245
rect 193630 558242 193690 558824
rect 190913 558240 193690 558242
rect 190913 558184 190918 558240
rect 190974 558184 193690 558240
rect 190913 558182 193690 558184
rect 190913 558179 190979 558182
rect 66161 558104 68938 558106
rect 66161 558048 66166 558104
rect 66222 558048 68938 558104
rect 66161 558046 68938 558048
rect 66161 558043 66227 558046
rect 191741 557834 191807 557837
rect 193630 557834 193690 558008
rect 253430 557970 253490 558280
rect 255589 557970 255655 557973
rect 253430 557968 255655 557970
rect 253430 557912 255594 557968
rect 255650 557912 255655 557968
rect 253430 557910 255655 557912
rect 255589 557907 255655 557910
rect 191741 557832 193690 557834
rect 191741 557776 191746 557832
rect 191802 557776 193690 557832
rect 191741 557774 193690 557776
rect 191741 557771 191807 557774
rect 67633 556610 67699 556613
rect 68878 556610 68938 557192
rect 94638 556882 94698 557464
rect 96705 556882 96771 556885
rect 97901 556882 97967 556885
rect 94638 556880 97967 556882
rect 94638 556824 96710 556880
rect 96766 556824 97906 556880
rect 97962 556824 97967 556880
rect 94638 556822 97967 556824
rect 96705 556819 96771 556822
rect 97901 556819 97967 556822
rect 67633 556608 68938 556610
rect 67633 556552 67638 556608
rect 67694 556552 68938 556608
rect 67633 556550 68938 556552
rect 67633 556547 67699 556550
rect 191741 556474 191807 556477
rect 193630 556474 193690 556920
rect 253430 556882 253490 557464
rect 255589 556882 255655 556885
rect 253430 556880 255655 556882
rect 253430 556824 255594 556880
rect 255650 556824 255655 556880
rect 253430 556822 255655 556824
rect 255589 556819 255655 556822
rect 191741 556472 193690 556474
rect 191741 556416 191746 556472
rect 191802 556416 193690 556472
rect 191741 556414 193690 556416
rect 191741 556411 191807 556414
rect 253430 556205 253490 556376
rect 253381 556200 253490 556205
rect 253381 556144 253386 556200
rect 253442 556144 253490 556200
rect 253381 556142 253490 556144
rect 253381 556139 253447 556142
rect 67357 555250 67423 555253
rect 68878 555250 68938 555832
rect 94638 555522 94698 556104
rect 94773 555522 94839 555525
rect 94638 555520 94839 555522
rect 94638 555464 94778 555520
rect 94834 555464 94839 555520
rect 94638 555462 94839 555464
rect 94773 555459 94839 555462
rect 67357 555248 68938 555250
rect 67357 555192 67362 555248
rect 67418 555192 68938 555248
rect 67357 555190 68938 555192
rect 187325 555250 187391 555253
rect 193630 555250 193690 556104
rect 187325 555248 193690 555250
rect 187325 555192 187330 555248
rect 187386 555192 193690 555248
rect 187325 555190 193690 555192
rect 67357 555187 67423 555190
rect 187325 555187 187391 555190
rect 190821 554842 190887 554845
rect 193630 554842 193690 555016
rect 253430 554978 253490 555560
rect 256601 554978 256667 554981
rect 253430 554976 256667 554978
rect 253430 554920 256606 554976
rect 256662 554920 256667 554976
rect 253430 554918 256667 554920
rect 256601 554915 256667 554918
rect 190821 554840 193690 554842
rect 190821 554784 190826 554840
rect 190882 554784 193690 554840
rect 190821 554782 193690 554784
rect 190821 554779 190887 554782
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 66713 553618 66779 553621
rect 68878 553618 68938 554200
rect 94638 554162 94698 554744
rect 96981 554162 97047 554165
rect 94638 554160 97047 554162
rect 94638 554104 96986 554160
rect 97042 554104 97047 554160
rect 94638 554102 97047 554104
rect 96981 554099 97047 554102
rect 116209 554026 116275 554029
rect 173157 554026 173223 554029
rect 66713 553616 68938 553618
rect 66713 553560 66718 553616
rect 66774 553560 68938 553616
rect 66713 553558 68938 553560
rect 103470 554024 173223 554026
rect 103470 553968 116214 554024
rect 116270 553968 173162 554024
rect 173218 553968 173223 554024
rect 103470 553966 173223 553968
rect 66713 553555 66779 553558
rect 96654 553420 96660 553484
rect 96724 553482 96730 553484
rect 103470 553482 103530 553966
rect 116209 553963 116275 553966
rect 173157 553963 173223 553966
rect 190913 553890 190979 553893
rect 193630 553890 193690 554200
rect 253430 554162 253490 554744
rect 255681 554162 255747 554165
rect 253430 554160 255747 554162
rect 253430 554104 255686 554160
rect 255742 554104 255747 554160
rect 253430 554102 255747 554104
rect 255681 554099 255747 554102
rect 190913 553888 193690 553890
rect 190913 553832 190918 553888
rect 190974 553832 193690 553888
rect 190913 553830 193690 553832
rect 190913 553827 190979 553830
rect 253430 553618 253490 553656
rect 255589 553618 255655 553621
rect 253430 553616 255655 553618
rect 253430 553560 255594 553616
rect 255650 553560 255655 553616
rect 253430 553558 255655 553560
rect 255589 553555 255655 553558
rect 96724 553422 103530 553482
rect 96724 553420 96730 553422
rect 67265 552258 67331 552261
rect 68878 552258 68938 552840
rect 94638 552802 94698 553384
rect 193121 553142 193187 553145
rect 193121 553140 193660 553142
rect 193121 553084 193126 553140
rect 193182 553084 193660 553140
rect 193121 553082 193660 553084
rect 193121 553079 193187 553082
rect 97901 552802 97967 552805
rect 94638 552800 97967 552802
rect 94638 552744 97906 552800
rect 97962 552744 97967 552800
rect 94638 552742 97967 552744
rect 253430 552802 253490 552840
rect 255589 552802 255655 552805
rect 253430 552800 255655 552802
rect 253430 552744 255594 552800
rect 255650 552744 255655 552800
rect 253430 552742 255655 552744
rect 97901 552739 97967 552742
rect 255589 552739 255655 552742
rect 67265 552256 68938 552258
rect 67265 552200 67270 552256
rect 67326 552200 68938 552256
rect 67265 552198 68938 552200
rect 67265 552195 67331 552198
rect 96613 552122 96679 552125
rect 97901 552122 97967 552125
rect 94638 552120 97967 552122
rect 94638 552064 96618 552120
rect 96674 552064 97906 552120
rect 97962 552064 97967 552120
rect 94638 552062 97967 552064
rect 94638 552024 94698 552062
rect 96613 552059 96679 552062
rect 97901 552059 97967 552062
rect 191741 552122 191807 552125
rect 193630 552122 193690 552296
rect 191741 552120 193690 552122
rect 191741 552064 191746 552120
rect 191802 552064 193690 552120
rect 191741 552062 193690 552064
rect 191741 552059 191807 552062
rect 101397 551986 101463 551989
rect 104934 551986 104940 551988
rect 101397 551984 104940 551986
rect 101397 551928 101402 551984
rect 101458 551928 104940 551984
rect 101397 551926 104940 551928
rect 101397 551923 101463 551926
rect 104934 551924 104940 551926
rect 105004 551924 105010 551988
rect 69246 550900 69306 551480
rect 96654 551306 96660 551308
rect 94638 551246 96660 551306
rect 69238 550836 69244 550900
rect 69308 550836 69314 550900
rect 94638 550664 94698 551246
rect 96654 551244 96660 551246
rect 96724 551244 96730 551308
rect 191373 550762 191439 550765
rect 193630 550762 193690 551208
rect 253430 551170 253490 551752
rect 256785 551170 256851 551173
rect 253430 551168 256851 551170
rect 253430 551112 256790 551168
rect 256846 551112 256851 551168
rect 253430 551110 256851 551112
rect 256785 551107 256851 551110
rect 583520 551020 584960 551260
rect 253430 550898 253490 550936
rect 255589 550898 255655 550901
rect 253430 550896 255655 550898
rect 253430 550840 255594 550896
rect 255650 550840 255655 550896
rect 253430 550838 255655 550840
rect 255589 550835 255655 550838
rect 191373 550760 193690 550762
rect 191373 550704 191378 550760
rect 191434 550704 193690 550760
rect 191373 550702 193690 550704
rect 191373 550699 191439 550702
rect 67766 549476 67772 549540
rect 67836 549538 67842 549540
rect 68878 549538 68938 550120
rect 191557 549810 191623 549813
rect 193630 549810 193690 550392
rect 255589 550218 255655 550221
rect 253430 550216 255655 550218
rect 253430 550160 255594 550216
rect 255650 550160 255655 550216
rect 253430 550158 255655 550160
rect 253430 549848 253490 550158
rect 255589 550155 255655 550158
rect 191557 549808 193690 549810
rect 191557 549752 191562 549808
rect 191618 549752 193690 549808
rect 191557 549750 193690 549752
rect 191557 549747 191623 549750
rect 67836 549478 68938 549538
rect 67836 549476 67842 549478
rect 100702 549402 100708 549404
rect 94638 549342 100708 549402
rect 94638 549304 94698 549342
rect 100702 549340 100708 549342
rect 100772 549340 100778 549404
rect 191741 549402 191807 549405
rect 191741 549400 193690 549402
rect 191741 549344 191746 549400
rect 191802 549344 193690 549400
rect 191741 549342 193690 549344
rect 191741 549339 191807 549342
rect 193630 549304 193690 549342
rect 65793 548314 65859 548317
rect 68878 548314 68938 548760
rect 65793 548312 68938 548314
rect 65793 548256 65798 548312
rect 65854 548256 68938 548312
rect 65793 548254 68938 548256
rect 65793 548251 65859 548254
rect 191557 548042 191623 548045
rect 193630 548042 193690 548488
rect 253430 548450 253490 549032
rect 255589 548450 255655 548453
rect 253430 548448 255655 548450
rect 253430 548392 255594 548448
rect 255650 548392 255655 548448
rect 253430 548390 255655 548392
rect 255589 548387 255655 548390
rect 191557 548040 193690 548042
rect 191557 547984 191562 548040
rect 191618 547984 193690 548040
rect 191557 547982 193690 547984
rect 191557 547979 191623 547982
rect 253430 547906 253490 547944
rect 254117 547906 254183 547909
rect 253430 547904 254183 547906
rect 253430 547848 254122 547904
rect 254178 547848 254183 547904
rect 253430 547846 254183 547848
rect 254117 547843 254183 547846
rect 65885 546818 65951 546821
rect 68878 546818 68938 547400
rect 94638 547090 94698 547672
rect 96838 547090 96844 547092
rect 94638 547030 96844 547090
rect 96838 547028 96844 547030
rect 96908 547028 96914 547092
rect 151670 547028 151676 547092
rect 151740 547090 151746 547092
rect 178769 547090 178835 547093
rect 151740 547088 178835 547090
rect 151740 547032 178774 547088
rect 178830 547032 178835 547088
rect 151740 547030 178835 547032
rect 151740 547028 151746 547030
rect 178769 547027 178835 547030
rect 191281 547090 191347 547093
rect 193630 547090 193690 547672
rect 191281 547088 193690 547090
rect 191281 547032 191286 547088
rect 191342 547032 193690 547088
rect 191281 547030 193690 547032
rect 191281 547027 191347 547030
rect 65885 546816 68938 546818
rect 65885 546760 65890 546816
rect 65946 546760 68938 546816
rect 65885 546758 68938 546760
rect 253430 546818 253490 547128
rect 255589 546818 255655 546821
rect 253430 546816 255655 546818
rect 253430 546760 255594 546816
rect 255650 546760 255655 546816
rect 253430 546758 255655 546760
rect 65885 546755 65951 546758
rect 255589 546755 255655 546758
rect 191557 546546 191623 546549
rect 193630 546546 193690 546584
rect 191557 546544 193690 546546
rect 191557 546488 191562 546544
rect 191618 546488 193690 546544
rect 191557 546486 193690 546488
rect 191557 546483 191623 546486
rect 66069 546410 66135 546413
rect 66069 546408 68938 546410
rect 66069 546352 66074 546408
rect 66130 546352 68938 546408
rect 66069 546350 68938 546352
rect 66069 546347 66135 546350
rect 68878 546040 68938 546350
rect 94638 545730 94698 546312
rect 253430 545866 253490 546312
rect 255589 545866 255655 545869
rect 253430 545864 255655 545866
rect 253430 545808 255594 545864
rect 255650 545808 255655 545864
rect 253430 545806 255655 545808
rect 255589 545803 255655 545806
rect 95325 545730 95391 545733
rect 94638 545728 95391 545730
rect 94638 545672 95330 545728
rect 95386 545672 95391 545728
rect 94638 545670 95391 545672
rect 95325 545667 95391 545670
rect 191189 545458 191255 545461
rect 193630 545458 193690 545768
rect 191189 545456 193690 545458
rect 191189 545400 191194 545456
rect 191250 545400 193690 545456
rect 191189 545398 193690 545400
rect 191189 545395 191255 545398
rect 253430 545186 253490 545224
rect 255681 545186 255747 545189
rect 253430 545184 255747 545186
rect 253430 545128 255686 545184
rect 255742 545128 255747 545184
rect 253430 545126 255747 545128
rect 255681 545123 255747 545126
rect 66805 544098 66871 544101
rect 68878 544098 68938 544680
rect 94638 544370 94698 544952
rect 97533 544370 97599 544373
rect 94638 544368 97599 544370
rect 94638 544312 97538 544368
rect 97594 544312 97599 544368
rect 94638 544310 97599 544312
rect 97533 544307 97599 544310
rect 191097 544234 191163 544237
rect 193630 544234 193690 544680
rect 191097 544232 193690 544234
rect 191097 544176 191102 544232
rect 191158 544176 193690 544232
rect 191097 544174 193690 544176
rect 191097 544171 191163 544174
rect 66805 544096 68938 544098
rect 66805 544040 66810 544096
rect 66866 544040 68938 544096
rect 66805 544038 68938 544040
rect 190637 544098 190703 544101
rect 253430 544098 253490 544408
rect 255589 544098 255655 544101
rect 190637 544096 193690 544098
rect 190637 544040 190642 544096
rect 190698 544040 193690 544096
rect 190637 544038 193690 544040
rect 253430 544096 255655 544098
rect 253430 544040 255594 544096
rect 255650 544040 255655 544096
rect 253430 544038 255655 544040
rect 66805 544035 66871 544038
rect 190637 544035 190703 544038
rect 193630 543864 193690 544038
rect 255589 544035 255655 544038
rect 66529 543146 66595 543149
rect 68878 543146 68938 543320
rect 66529 543144 68938 543146
rect 66529 543088 66534 543144
rect 66590 543088 68938 543144
rect 66529 543086 68938 543088
rect 66529 543083 66595 543086
rect 94638 543010 94698 543592
rect 97533 543010 97599 543013
rect 94638 543008 97599 543010
rect 94638 542952 97538 543008
rect 97594 542952 97599 543008
rect 94638 542950 97599 542952
rect 97533 542947 97599 542950
rect 191557 542602 191623 542605
rect 193630 542602 193690 542776
rect 253430 542738 253490 543320
rect 270534 542738 270540 542740
rect 253430 542678 270540 542738
rect 270534 542676 270540 542678
rect 270604 542676 270610 542740
rect 191557 542600 193690 542602
rect 191557 542544 191562 542600
rect 191618 542544 193690 542600
rect 191557 542542 193690 542544
rect 191557 542539 191623 542542
rect 253430 542466 253490 542504
rect 254209 542466 254275 542469
rect 253430 542464 254275 542466
rect 253430 542408 254214 542464
rect 254270 542408 254275 542464
rect 253430 542406 254275 542408
rect 254209 542403 254275 542406
rect 69422 542132 69428 542196
rect 69492 542132 69498 542196
rect 15837 541106 15903 541109
rect 69430 541106 69490 542132
rect 94638 541786 94698 542232
rect 96889 541786 96955 541789
rect 97901 541786 97967 541789
rect 94638 541784 97967 541786
rect 94638 541728 96894 541784
rect 96950 541728 97906 541784
rect 97962 541728 97967 541784
rect 94638 541726 97967 541728
rect 96889 541723 96955 541726
rect 97901 541723 97967 541726
rect 190821 541514 190887 541517
rect 193630 541514 193690 541960
rect 190821 541512 193690 541514
rect 190821 541456 190826 541512
rect 190882 541456 193690 541512
rect 190821 541454 193690 541456
rect 190821 541451 190887 541454
rect 253430 541242 253490 541416
rect 255589 541242 255655 541245
rect 253430 541240 255655 541242
rect 253430 541184 255594 541240
rect 255650 541184 255655 541240
rect 253430 541182 255655 541184
rect 255589 541179 255655 541182
rect 15837 541104 69490 541106
rect 15837 541048 15842 541104
rect 15898 541048 69490 541104
rect 15837 541046 69490 541048
rect 15837 541043 15903 541046
rect -960 540684 480 540924
rect 66621 540018 66687 540021
rect 68878 540018 68938 540600
rect 66621 540016 68938 540018
rect 66621 539960 66626 540016
rect 66682 539960 68938 540016
rect 66621 539958 68938 539960
rect 66621 539955 66687 539958
rect 94270 539885 94330 540872
rect 191465 540290 191531 540293
rect 193630 540290 193690 540872
rect 191465 540288 193690 540290
rect 191465 540232 191470 540288
rect 191526 540232 193690 540288
rect 191465 540230 193690 540232
rect 191465 540227 191531 540230
rect 191557 540154 191623 540157
rect 191557 540152 193690 540154
rect 191557 540096 191562 540152
rect 191618 540096 193690 540152
rect 191557 540094 193690 540096
rect 191557 540091 191623 540094
rect 193630 540056 193690 540094
rect 94270 539880 94379 539885
rect 94270 539824 94318 539880
rect 94374 539824 94379 539880
rect 94270 539822 94379 539824
rect 253430 539882 253490 540600
rect 253430 539822 258090 539882
rect 94313 539819 94379 539822
rect 89713 539746 89779 539749
rect 180609 539746 180675 539749
rect 89713 539744 180675 539746
rect 89713 539688 89718 539744
rect 89774 539688 180614 539744
rect 180670 539688 180675 539744
rect 89713 539686 180675 539688
rect 258030 539746 258090 539822
rect 276238 539746 276244 539748
rect 258030 539686 276244 539746
rect 89713 539683 89779 539686
rect 180609 539683 180675 539686
rect 276238 539684 276244 539686
rect 276308 539684 276314 539748
rect 94638 538933 94698 539512
rect 94589 538928 94698 538933
rect 94589 538872 94594 538928
rect 94650 538872 94698 538928
rect 94589 538870 94698 538872
rect 253430 538930 253490 539512
rect 255589 538930 255655 538933
rect 253430 538928 255655 538930
rect 253430 538872 255594 538928
rect 255650 538872 255655 538928
rect 253430 538870 255655 538872
rect 94589 538867 94655 538870
rect 255589 538867 255655 538870
rect 67766 538732 67772 538796
rect 67836 538794 67842 538796
rect 82854 538794 82860 538796
rect 67836 538734 82860 538794
rect 67836 538732 67842 538734
rect 82854 538732 82860 538734
rect 82924 538732 82930 538796
rect 243537 538794 243603 538797
rect 253933 538794 253999 538797
rect 243537 538792 253999 538794
rect 243537 538736 243542 538792
rect 243598 538736 253938 538792
rect 253994 538736 253999 538792
rect 243537 538734 253999 538736
rect 243537 538731 243603 538734
rect 253933 538731 253999 538734
rect 80145 538386 80211 538389
rect 179505 538386 179571 538389
rect 80145 538384 180810 538386
rect 80145 538328 80150 538384
rect 80206 538328 179510 538384
rect 179566 538328 180810 538384
rect 80145 538326 180810 538328
rect 80145 538323 80211 538326
rect 179505 538323 179571 538326
rect 180750 538250 180810 538326
rect 207381 538250 207447 538253
rect 180750 538248 207447 538250
rect 180750 538192 207386 538248
rect 207442 538192 207447 538248
rect 180750 538190 207447 538192
rect 207381 538187 207447 538190
rect 223573 538250 223639 538253
rect 224677 538250 224743 538253
rect 582925 538250 582991 538253
rect 223573 538248 582991 538250
rect 223573 538192 223578 538248
rect 223634 538192 224682 538248
rect 224738 538192 582930 538248
rect 582986 538192 582991 538248
rect 223573 538190 582991 538192
rect 223573 538187 223639 538190
rect 224677 538187 224743 538190
rect 582925 538187 582991 538190
rect 84009 538114 84075 538117
rect 202965 538114 203031 538117
rect 84009 538112 203031 538114
rect 84009 538056 84014 538112
rect 84070 538056 202970 538112
rect 203026 538056 203031 538112
rect 84009 538054 203031 538056
rect 84009 538051 84075 538054
rect 202965 538051 203031 538054
rect 188429 537978 188495 537981
rect 255497 537978 255563 537981
rect 188429 537976 255563 537978
rect 188429 537920 188434 537976
rect 188490 537920 255502 537976
rect 255558 537920 255563 537976
rect 188429 537918 255563 537920
rect 188429 537915 188495 537918
rect 255497 537915 255563 537918
rect 582465 537842 582531 537845
rect 583520 537842 584960 537932
rect 582465 537840 584960 537842
rect 582465 537784 582470 537840
rect 582526 537784 584960 537840
rect 582465 537782 584960 537784
rect 582465 537779 582531 537782
rect 583520 537692 584960 537782
rect 202965 536890 203031 536893
rect 203517 536890 203583 536893
rect 202965 536888 203583 536890
rect 202965 536832 202970 536888
rect 203026 536832 203522 536888
rect 203578 536832 203583 536888
rect 202965 536830 203583 536832
rect 202965 536827 203031 536830
rect 203517 536827 203583 536830
rect 87689 536754 87755 536757
rect 215385 536754 215451 536757
rect 87689 536752 215451 536754
rect 87689 536696 87694 536752
rect 87750 536696 215390 536752
rect 215446 536696 215451 536752
rect 87689 536694 215451 536696
rect 87689 536691 87755 536694
rect 215385 536691 215451 536694
rect 199377 536618 199443 536621
rect 271137 536618 271203 536621
rect 199377 536616 271203 536618
rect 199377 536560 199382 536616
rect 199438 536560 271142 536616
rect 271198 536560 271203 536616
rect 199377 536558 271203 536560
rect 199377 536555 199443 536558
rect 271137 536555 271203 536558
rect 212441 536482 212507 536485
rect 280797 536482 280863 536485
rect 212441 536480 280863 536482
rect 212441 536424 212446 536480
rect 212502 536424 280802 536480
rect 280858 536424 280863 536480
rect 212441 536422 280863 536424
rect 212441 536419 212507 536422
rect 280797 536419 280863 536422
rect 188337 536074 188403 536077
rect 195421 536074 195487 536077
rect 188337 536072 195487 536074
rect 188337 536016 188342 536072
rect 188398 536016 195426 536072
rect 195482 536016 195487 536072
rect 188337 536014 195487 536016
rect 188337 536011 188403 536014
rect 195421 536011 195487 536014
rect 253197 536074 253263 536077
rect 262438 536074 262444 536076
rect 253197 536072 262444 536074
rect 253197 536016 253202 536072
rect 253258 536016 262444 536072
rect 253197 536014 262444 536016
rect 253197 536011 253263 536014
rect 262438 536012 262444 536014
rect 262508 536012 262514 536076
rect 194133 535530 194199 535533
rect 197445 535530 197511 535533
rect 194133 535528 197511 535530
rect 194133 535472 194138 535528
rect 194194 535472 197450 535528
rect 197506 535472 197511 535528
rect 194133 535470 197511 535472
rect 194133 535467 194199 535470
rect 197445 535467 197511 535470
rect 206134 535468 206140 535532
rect 206204 535530 206210 535532
rect 208117 535530 208183 535533
rect 206204 535528 208183 535530
rect 206204 535472 208122 535528
rect 208178 535472 208183 535528
rect 206204 535470 208183 535472
rect 206204 535468 206210 535470
rect 208117 535467 208183 535470
rect 222837 535530 222903 535533
rect 226517 535530 226583 535533
rect 222837 535528 226583 535530
rect 222837 535472 222842 535528
rect 222898 535472 226522 535528
rect 226578 535472 226583 535528
rect 222837 535470 226583 535472
rect 222837 535467 222903 535470
rect 226517 535467 226583 535470
rect 242934 535468 242940 535532
rect 243004 535530 243010 535532
rect 243629 535530 243695 535533
rect 243004 535528 243695 535530
rect 243004 535472 243634 535528
rect 243690 535472 243695 535528
rect 243004 535470 243695 535472
rect 243004 535468 243010 535470
rect 243629 535467 243695 535470
rect 151077 535394 151143 535397
rect 199377 535394 199443 535397
rect 151077 535392 199443 535394
rect 151077 535336 151082 535392
rect 151138 535336 199382 535392
rect 199438 535336 199443 535392
rect 151077 535334 199443 535336
rect 151077 535331 151143 535334
rect 199377 535331 199443 535334
rect 65885 534714 65951 534717
rect 104198 534714 104204 534716
rect 65885 534712 104204 534714
rect 65885 534656 65890 534712
rect 65946 534656 104204 534712
rect 65885 534654 104204 534656
rect 65885 534651 65951 534654
rect 104198 534652 104204 534654
rect 104268 534652 104274 534716
rect 222929 534034 222995 534037
rect 229645 534034 229711 534037
rect 222929 534032 229711 534034
rect 222929 533976 222934 534032
rect 222990 533976 229650 534032
rect 229706 533976 229711 534032
rect 222929 533974 229711 533976
rect 222929 533971 222995 533974
rect 229645 533971 229711 533974
rect 66110 533292 66116 533356
rect 66180 533354 66186 533356
rect 84285 533354 84351 533357
rect 66180 533352 84351 533354
rect 66180 533296 84290 533352
rect 84346 533296 84351 533352
rect 66180 533294 84351 533296
rect 66180 533292 66186 533294
rect 84285 533291 84351 533294
rect 96429 533354 96495 533357
rect 111742 533354 111748 533356
rect 96429 533352 111748 533354
rect 96429 533296 96434 533352
rect 96490 533296 111748 533352
rect 96429 533294 111748 533296
rect 96429 533291 96495 533294
rect 111742 533292 111748 533294
rect 111812 533292 111818 533356
rect 152457 533354 152523 533357
rect 212625 533354 212691 533357
rect 152457 533352 212691 533354
rect 152457 533296 152462 533352
rect 152518 533296 212630 533352
rect 212686 533296 212691 533352
rect 152457 533294 212691 533296
rect 152457 533291 152523 533294
rect 212625 533291 212691 533294
rect 213269 533354 213335 533357
rect 218973 533354 219039 533357
rect 213269 533352 219039 533354
rect 213269 533296 213274 533352
rect 213330 533296 218978 533352
rect 219034 533296 219039 533352
rect 213269 533294 219039 533296
rect 213269 533291 213335 533294
rect 218973 533291 219039 533294
rect 220077 533354 220143 533357
rect 223941 533354 224007 533357
rect 220077 533352 224007 533354
rect 220077 533296 220082 533352
rect 220138 533296 223946 533352
rect 224002 533296 224007 533352
rect 220077 533294 224007 533296
rect 220077 533291 220143 533294
rect 223941 533291 224007 533294
rect 232497 533354 232563 533357
rect 235349 533354 235415 533357
rect 232497 533352 235415 533354
rect 232497 533296 232502 533352
rect 232558 533296 235354 533352
rect 235410 533296 235415 533352
rect 232497 533294 235415 533296
rect 232497 533291 232563 533294
rect 235349 533291 235415 533294
rect 250069 533354 250135 533357
rect 257061 533354 257127 533357
rect 250069 533352 257127 533354
rect 250069 533296 250074 533352
rect 250130 533296 257066 533352
rect 257122 533296 257127 533352
rect 250069 533294 257127 533296
rect 250069 533291 250135 533294
rect 257061 533291 257127 533294
rect 194685 531994 194751 531997
rect 244406 531994 244412 531996
rect 194685 531992 244412 531994
rect 194685 531936 194690 531992
rect 194746 531936 244412 531992
rect 194685 531934 244412 531936
rect 194685 531931 194751 531934
rect 244406 531932 244412 531934
rect 244476 531932 244482 531996
rect 249006 531252 249012 531316
rect 249076 531314 249082 531316
rect 256785 531314 256851 531317
rect 249076 531312 256851 531314
rect 249076 531256 256790 531312
rect 256846 531256 256851 531312
rect 249076 531254 256851 531256
rect 249076 531252 249082 531254
rect 256785 531251 256851 531254
rect 88333 530770 88399 530773
rect 106774 530770 106780 530772
rect 88333 530768 106780 530770
rect 88333 530712 88338 530768
rect 88394 530712 106780 530768
rect 88333 530710 106780 530712
rect 88333 530707 88399 530710
rect 106774 530708 106780 530710
rect 106844 530708 106850 530772
rect 69790 530572 69796 530636
rect 69860 530634 69866 530636
rect 88926 530634 88932 530636
rect 69860 530574 88932 530634
rect 69860 530572 69866 530574
rect 88926 530572 88932 530574
rect 88996 530572 89002 530636
rect 177798 530572 177804 530636
rect 177868 530634 177874 530636
rect 204437 530634 204503 530637
rect 177868 530632 204503 530634
rect 177868 530576 204442 530632
rect 204498 530576 204503 530632
rect 177868 530574 204503 530576
rect 177868 530572 177874 530574
rect 204437 530571 204503 530574
rect 205081 530634 205147 530637
rect 219525 530634 219591 530637
rect 205081 530632 219591 530634
rect 205081 530576 205086 530632
rect 205142 530576 219530 530632
rect 219586 530576 219591 530632
rect 205081 530574 219591 530576
rect 205081 530571 205147 530574
rect 219525 530571 219591 530574
rect 168189 529138 168255 529141
rect 198733 529138 198799 529141
rect 168189 529136 198799 529138
rect 168189 529080 168194 529136
rect 168250 529080 198738 529136
rect 198794 529080 198799 529136
rect 168189 529078 198799 529080
rect 168189 529075 168255 529078
rect 198733 529075 198799 529078
rect 232998 529076 233004 529140
rect 233068 529138 233074 529140
rect 249742 529138 249748 529140
rect 233068 529078 249748 529138
rect 233068 529076 233074 529078
rect 249742 529076 249748 529078
rect 249812 529076 249818 529140
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 67817 527778 67883 527781
rect 97022 527778 97028 527780
rect 67817 527776 97028 527778
rect 67817 527720 67822 527776
rect 67878 527720 97028 527776
rect 67817 527718 97028 527720
rect 67817 527715 67883 527718
rect 97022 527716 97028 527718
rect 97092 527716 97098 527780
rect 249793 527098 249859 527101
rect 84150 527096 249859 527098
rect 84150 527040 249798 527096
rect 249854 527040 249859 527096
rect 84150 527038 249859 527040
rect 81014 526764 81020 526828
rect 81084 526826 81090 526828
rect 84150 526826 84210 527038
rect 249793 527035 249859 527038
rect 81084 526766 84210 526826
rect 81084 526764 81090 526766
rect 81014 525812 81020 525876
rect 81084 525874 81090 525876
rect 81341 525874 81407 525877
rect 81084 525872 81407 525874
rect 81084 525816 81346 525872
rect 81402 525816 81407 525872
rect 81084 525814 81407 525816
rect 81084 525812 81090 525814
rect 81341 525811 81407 525814
rect 65977 525058 66043 525061
rect 68921 525058 68987 525061
rect 258257 525058 258323 525061
rect 65977 525056 258323 525058
rect 65977 525000 65982 525056
rect 66038 525000 68926 525056
rect 68982 525000 258262 525056
rect 258318 525000 258323 525056
rect 65977 524998 258323 525000
rect 65977 524995 66043 524998
rect 68921 524995 68987 524998
rect 258257 524995 258323 524998
rect 582741 524514 582807 524517
rect 583520 524514 584960 524604
rect 582741 524512 584960 524514
rect 582741 524456 582746 524512
rect 582802 524456 584960 524512
rect 582741 524454 584960 524456
rect 582741 524451 582807 524454
rect 583520 524364 584960 524454
rect 77150 523636 77156 523700
rect 77220 523698 77226 523700
rect 94773 523698 94839 523701
rect 77220 523696 94839 523698
rect 77220 523640 94778 523696
rect 94834 523640 94839 523696
rect 77220 523638 94839 523640
rect 77220 523636 77226 523638
rect 94773 523635 94839 523638
rect 148869 523698 148935 523701
rect 213269 523698 213335 523701
rect 148869 523696 213335 523698
rect 148869 523640 148874 523696
rect 148930 523640 213274 523696
rect 213330 523640 213335 523696
rect 148869 523638 213335 523640
rect 148869 523635 148935 523638
rect 213269 523635 213335 523638
rect 226190 523636 226196 523700
rect 226260 523698 226266 523700
rect 245694 523698 245700 523700
rect 226260 523638 245700 523698
rect 226260 523636 226266 523638
rect 245694 523636 245700 523638
rect 245764 523636 245770 523700
rect 219934 522276 219940 522340
rect 220004 522338 220010 522340
rect 231117 522338 231183 522341
rect 220004 522336 231183 522338
rect 220004 522280 231122 522336
rect 231178 522280 231183 522336
rect 220004 522278 231183 522280
rect 220004 522276 220010 522278
rect 231117 522275 231183 522278
rect 72734 520916 72740 520980
rect 72804 520978 72810 520980
rect 95233 520978 95299 520981
rect 72804 520976 95299 520978
rect 72804 520920 95238 520976
rect 95294 520920 95299 520976
rect 72804 520918 95299 520920
rect 72804 520916 72810 520918
rect 95233 520915 95299 520918
rect 60549 519482 60615 519485
rect 96838 519482 96844 519484
rect 60549 519480 96844 519482
rect 60549 519424 60554 519480
rect 60610 519424 96844 519480
rect 60549 519422 96844 519424
rect 60549 519419 60615 519422
rect 96838 519420 96844 519422
rect 96908 519420 96914 519484
rect 222694 518060 222700 518124
rect 222764 518122 222770 518124
rect 244273 518122 244339 518125
rect 222764 518120 244339 518122
rect 222764 518064 244278 518120
rect 244334 518064 244339 518120
rect 222764 518062 244339 518064
rect 222764 518060 222770 518062
rect 244273 518059 244339 518062
rect 69606 516700 69612 516764
rect 69676 516762 69682 516764
rect 115289 516762 115355 516765
rect 69676 516760 115355 516762
rect 69676 516704 115294 516760
rect 115350 516704 115355 516760
rect 69676 516702 115355 516704
rect 69676 516700 69682 516702
rect 115289 516699 115355 516702
rect 147489 516762 147555 516765
rect 249006 516762 249012 516764
rect 147489 516760 249012 516762
rect 147489 516704 147494 516760
rect 147550 516704 249012 516760
rect 147489 516702 249012 516704
rect 147489 516699 147555 516702
rect 249006 516700 249012 516702
rect 249076 516700 249082 516764
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 169201 513362 169267 513365
rect 169334 513362 169340 513364
rect 169201 513360 169340 513362
rect 169201 513304 169206 513360
rect 169262 513304 169340 513360
rect 169201 513302 169340 513304
rect 169201 513299 169267 513302
rect 169334 513300 169340 513302
rect 169404 513300 169410 513364
rect 203517 512682 203583 512685
rect 218646 512682 218652 512684
rect 203517 512680 218652 512682
rect 203517 512624 203522 512680
rect 203578 512624 218652 512680
rect 203517 512622 218652 512624
rect 203517 512619 203583 512622
rect 218646 512620 218652 512622
rect 218716 512620 218722 512684
rect 163630 511260 163636 511324
rect 163700 511322 163706 511324
rect 188337 511322 188403 511325
rect 163700 511320 188403 511322
rect 163700 511264 188342 511320
rect 188398 511264 188403 511320
rect 163700 511262 188403 511264
rect 163700 511260 163706 511262
rect 188337 511259 188403 511262
rect 582649 511322 582715 511325
rect 583520 511322 584960 511412
rect 582649 511320 584960 511322
rect 582649 511264 582654 511320
rect 582710 511264 584960 511320
rect 582649 511262 584960 511264
rect 582649 511259 582715 511262
rect 583520 511172 584960 511262
rect 202137 509826 202203 509829
rect 216622 509826 216628 509828
rect 202137 509824 216628 509826
rect 202137 509768 202142 509824
rect 202198 509768 216628 509824
rect 202137 509766 216628 509768
rect 202137 509763 202203 509766
rect 216622 509764 216628 509766
rect 216692 509764 216698 509828
rect 203190 508404 203196 508468
rect 203260 508466 203266 508468
rect 254710 508466 254716 508468
rect 203260 508406 254716 508466
rect 203260 508404 203266 508406
rect 254710 508404 254716 508406
rect 254780 508404 254786 508468
rect 253933 507922 253999 507925
rect 254526 507922 254532 507924
rect 253933 507920 254532 507922
rect 253933 507864 253938 507920
rect 253994 507864 254532 507920
rect 253933 507862 254532 507864
rect 253933 507859 253999 507862
rect 254526 507860 254532 507862
rect 254596 507860 254602 507924
rect 159766 502964 159772 503028
rect 159836 503026 159842 503028
rect 170397 503026 170463 503029
rect 159836 503024 170463 503026
rect 159836 502968 170402 503024
rect 170458 502968 170463 503024
rect 159836 502966 170463 502968
rect 159836 502964 159842 502966
rect 170397 502963 170463 502966
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 234613 500170 234679 500173
rect 244774 500170 244780 500172
rect 234613 500168 244780 500170
rect 234613 500112 234618 500168
rect 234674 500112 244780 500168
rect 234613 500110 244780 500112
rect 234613 500107 234679 500110
rect 244774 500108 244780 500110
rect 244844 500108 244850 500172
rect 195421 498810 195487 498813
rect 229686 498810 229692 498812
rect 195421 498808 229692 498810
rect 195421 498752 195426 498808
rect 195482 498752 229692 498808
rect 195421 498750 229692 498752
rect 195421 498747 195487 498750
rect 229686 498748 229692 498750
rect 229756 498748 229762 498812
rect 583520 497844 584960 498084
rect 235901 496090 235967 496093
rect 252502 496090 252508 496092
rect 235901 496088 252508 496090
rect 235901 496032 235906 496088
rect 235962 496032 252508 496088
rect 235901 496030 252508 496032
rect 235901 496027 235967 496030
rect 252502 496028 252508 496030
rect 252572 496028 252578 496092
rect 216438 493444 216444 493508
rect 216508 493506 216514 493508
rect 228449 493506 228515 493509
rect 216508 493504 228515 493506
rect 216508 493448 228454 493504
rect 228510 493448 228515 493504
rect 216508 493446 228515 493448
rect 216508 493444 216514 493446
rect 228449 493443 228515 493446
rect 197118 493308 197124 493372
rect 197188 493370 197194 493372
rect 252502 493370 252508 493372
rect 197188 493310 252508 493370
rect 197188 493308 197194 493310
rect 252502 493308 252508 493310
rect 252572 493308 252578 493372
rect 210233 492826 210299 492829
rect 210366 492826 210372 492828
rect 210233 492824 210372 492826
rect 210233 492768 210238 492824
rect 210294 492768 210372 492824
rect 210233 492766 210372 492768
rect 210233 492763 210299 492766
rect 210366 492764 210372 492766
rect 210436 492764 210442 492828
rect 251030 492628 251036 492692
rect 251100 492690 251106 492692
rect 251357 492690 251423 492693
rect 251100 492688 251423 492690
rect 251100 492632 251362 492688
rect 251418 492632 251423 492688
rect 251100 492630 251423 492632
rect 251100 492628 251106 492630
rect 251357 492627 251423 492630
rect 195329 491874 195395 491877
rect 226926 491874 226932 491876
rect 195329 491872 226932 491874
rect 195329 491816 195334 491872
rect 195390 491816 226932 491872
rect 195329 491814 226932 491816
rect 195329 491811 195395 491814
rect 226926 491812 226932 491814
rect 226996 491812 227002 491876
rect 231209 491194 231275 491197
rect 237966 491194 237972 491196
rect 231209 491192 237972 491194
rect 231209 491136 231214 491192
rect 231270 491136 237972 491192
rect 231209 491134 237972 491136
rect 231209 491131 231275 491134
rect 237966 491132 237972 491134
rect 238036 491132 238042 491196
rect 197997 490650 198063 490653
rect 223798 490650 223804 490652
rect 197997 490648 223804 490650
rect 197997 490592 198002 490648
rect 198058 490592 223804 490648
rect 197997 490590 223804 490592
rect 197997 490587 198063 490590
rect 223798 490588 223804 490590
rect 223868 490588 223874 490652
rect 169518 490452 169524 490516
rect 169588 490514 169594 490516
rect 227713 490514 227779 490517
rect 169588 490512 227779 490514
rect 169588 490456 227718 490512
rect 227774 490456 227779 490512
rect 169588 490454 227779 490456
rect 169588 490452 169594 490454
rect 227713 490451 227779 490454
rect 203609 489290 203675 489293
rect 226374 489290 226380 489292
rect 203609 489288 226380 489290
rect 203609 489232 203614 489288
rect 203670 489232 226380 489288
rect 203609 489230 226380 489232
rect 203609 489227 203675 489230
rect 226374 489228 226380 489230
rect 226444 489228 226450 489292
rect 158478 489092 158484 489156
rect 158548 489154 158554 489156
rect 169109 489154 169175 489157
rect 158548 489152 169175 489154
rect 158548 489096 169114 489152
rect 169170 489096 169175 489152
rect 158548 489094 169175 489096
rect 158548 489092 158554 489094
rect 169109 489091 169175 489094
rect 172094 489092 172100 489156
rect 172164 489154 172170 489156
rect 209037 489154 209103 489157
rect 172164 489152 209103 489154
rect 172164 489096 209042 489152
rect 209098 489096 209103 489152
rect 172164 489094 209103 489096
rect 172164 489092 172170 489094
rect 209037 489091 209103 489094
rect -960 488596 480 488836
rect 180190 485828 180196 485892
rect 180260 485890 180266 485892
rect 180609 485890 180675 485893
rect 250437 485890 250503 485893
rect 180260 485888 250503 485890
rect 180260 485832 180614 485888
rect 180670 485832 250442 485888
rect 250498 485832 250503 485888
rect 180260 485830 250503 485832
rect 180260 485828 180266 485830
rect 180609 485827 180675 485830
rect 250437 485827 250503 485830
rect 183001 485074 183067 485077
rect 218697 485074 218763 485077
rect 183001 485072 218763 485074
rect 183001 485016 183006 485072
rect 183062 485016 218702 485072
rect 218758 485016 218763 485072
rect 183001 485014 218763 485016
rect 183001 485011 183067 485014
rect 218697 485011 218763 485014
rect 239254 485012 239260 485076
rect 239324 485074 239330 485076
rect 247125 485074 247191 485077
rect 239324 485072 247191 485074
rect 239324 485016 247130 485072
rect 247186 485016 247191 485072
rect 239324 485014 247191 485016
rect 239324 485012 239330 485014
rect 247125 485011 247191 485014
rect 579797 484666 579863 484669
rect 583520 484666 584960 484756
rect 579797 484664 584960 484666
rect 579797 484608 579802 484664
rect 579858 484608 584960 484664
rect 579797 484606 584960 484608
rect 579797 484603 579863 484606
rect 583520 484516 584960 484606
rect 88977 484394 89043 484397
rect 89294 484394 89300 484396
rect 88977 484392 89300 484394
rect 88977 484336 88982 484392
rect 89038 484336 89300 484392
rect 88977 484334 89300 484336
rect 88977 484331 89043 484334
rect 89294 484332 89300 484334
rect 89364 484332 89370 484396
rect 156638 483652 156644 483716
rect 156708 483714 156714 483716
rect 167637 483714 167703 483717
rect 156708 483712 167703 483714
rect 156708 483656 167642 483712
rect 167698 483656 167703 483712
rect 156708 483654 167703 483656
rect 156708 483652 156714 483654
rect 167637 483651 167703 483654
rect 202873 483714 202939 483717
rect 215334 483714 215340 483716
rect 202873 483712 215340 483714
rect 202873 483656 202878 483712
rect 202934 483656 215340 483712
rect 202873 483654 215340 483656
rect 202873 483651 202939 483654
rect 215334 483652 215340 483654
rect 215404 483652 215410 483716
rect 88977 483034 89043 483037
rect 209037 483034 209103 483037
rect 88977 483032 209103 483034
rect 88977 482976 88982 483032
rect 89038 482976 209042 483032
rect 209098 482976 209103 483032
rect 88977 482974 209103 482976
rect 88977 482971 89043 482974
rect 209037 482971 209103 482974
rect 75678 482156 75684 482220
rect 75748 482218 75754 482220
rect 94589 482218 94655 482221
rect 75748 482216 94655 482218
rect 75748 482160 94594 482216
rect 94650 482160 94655 482216
rect 75748 482158 94655 482160
rect 75748 482156 75754 482158
rect 94589 482155 94655 482158
rect 175089 482218 175155 482221
rect 206134 482218 206140 482220
rect 175089 482216 206140 482218
rect 175089 482160 175094 482216
rect 175150 482160 206140 482216
rect 175089 482158 206140 482160
rect 175089 482155 175155 482158
rect 206134 482156 206140 482158
rect 206204 482156 206210 482220
rect 218697 482218 218763 482221
rect 236494 482218 236500 482220
rect 218697 482216 236500 482218
rect 218697 482160 218702 482216
rect 218758 482160 236500 482216
rect 218697 482158 236500 482160
rect 218697 482155 218763 482158
rect 236494 482156 236500 482158
rect 236564 482156 236570 482220
rect 240777 481540 240843 481541
rect 240726 481476 240732 481540
rect 240796 481538 240843 481540
rect 240796 481536 240888 481538
rect 240838 481480 240888 481536
rect 240796 481478 240888 481480
rect 240796 481476 240843 481478
rect 249006 481476 249012 481540
rect 249076 481538 249082 481540
rect 253381 481538 253447 481541
rect 249076 481536 253447 481538
rect 249076 481480 253386 481536
rect 253442 481480 253447 481536
rect 249076 481478 253447 481480
rect 249076 481476 249082 481478
rect 240777 481475 240843 481476
rect 253381 481475 253447 481478
rect 166206 480796 166212 480860
rect 166276 480858 166282 480860
rect 185669 480858 185735 480861
rect 166276 480856 185735 480858
rect 166276 480800 185674 480856
rect 185730 480800 185735 480856
rect 166276 480798 185735 480800
rect 166276 480796 166282 480798
rect 185669 480795 185735 480798
rect 231945 480858 232011 480861
rect 265249 480858 265315 480861
rect 231945 480856 265315 480858
rect 231945 480800 231950 480856
rect 232006 480800 265254 480856
rect 265310 480800 265315 480856
rect 231945 480798 265315 480800
rect 231945 480795 232011 480798
rect 265249 480795 265315 480798
rect 162526 479436 162532 479500
rect 162596 479498 162602 479500
rect 231853 479498 231919 479501
rect 162596 479496 231919 479498
rect 162596 479440 231858 479496
rect 231914 479440 231919 479496
rect 162596 479438 231919 479440
rect 162596 479436 162602 479438
rect 231853 479435 231919 479438
rect 195237 478138 195303 478141
rect 234654 478138 234660 478140
rect 195237 478136 234660 478138
rect 195237 478080 195242 478136
rect 195298 478080 234660 478136
rect 195237 478078 234660 478080
rect 195237 478075 195303 478078
rect 234654 478076 234660 478078
rect 234724 478076 234730 478140
rect 176510 476716 176516 476780
rect 176580 476778 176586 476780
rect 195329 476778 195395 476781
rect 176580 476776 195395 476778
rect 176580 476720 195334 476776
rect 195390 476720 195395 476776
rect 176580 476718 195395 476720
rect 176580 476716 176586 476718
rect 195329 476715 195395 476718
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 186221 475418 186287 475421
rect 207054 475418 207060 475420
rect 186221 475416 207060 475418
rect 186221 475360 186226 475416
rect 186282 475360 207060 475416
rect 186221 475358 207060 475360
rect 186221 475355 186287 475358
rect 207054 475356 207060 475358
rect 207124 475356 207130 475420
rect 142889 475282 142955 475285
rect 143349 475282 143415 475285
rect 142889 475280 143415 475282
rect 142889 475224 142894 475280
rect 142950 475224 143354 475280
rect 143410 475224 143415 475280
rect 142889 475222 143415 475224
rect 142889 475219 142955 475222
rect 143349 475219 143415 475222
rect 143349 474874 143415 474877
rect 231301 474874 231367 474877
rect 143349 474872 231367 474874
rect 143349 474816 143354 474872
rect 143410 474816 231306 474872
rect 231362 474816 231367 474872
rect 143349 474814 231367 474816
rect 143349 474811 143415 474814
rect 231301 474811 231367 474814
rect 181478 473996 181484 474060
rect 181548 474058 181554 474060
rect 220854 474058 220860 474060
rect 181548 473998 220860 474058
rect 181548 473996 181554 473998
rect 220854 473996 220860 473998
rect 220924 473996 220930 474060
rect 133137 473242 133203 473245
rect 133689 473242 133755 473245
rect 133137 473240 133755 473242
rect 133137 473184 133142 473240
rect 133198 473184 133694 473240
rect 133750 473184 133755 473240
rect 133137 473182 133755 473184
rect 133137 473179 133203 473182
rect 133689 473179 133755 473182
rect 253933 472154 253999 472157
rect 287094 472154 287100 472156
rect 253933 472152 287100 472154
rect 253933 472096 253938 472152
rect 253994 472096 287100 472152
rect 253933 472094 287100 472096
rect 253933 472091 253999 472094
rect 287094 472092 287100 472094
rect 287164 472154 287170 472156
rect 287605 472154 287671 472157
rect 287164 472152 287671 472154
rect 287164 472096 287610 472152
rect 287666 472096 287671 472152
rect 287164 472094 287671 472096
rect 287164 472092 287170 472094
rect 287605 472091 287671 472094
rect 133137 472018 133203 472021
rect 291377 472018 291443 472021
rect 133137 472016 291443 472018
rect 133137 471960 133142 472016
rect 133198 471960 291382 472016
rect 291438 471960 291443 472016
rect 133137 471958 291443 471960
rect 133137 471955 133203 471958
rect 291377 471955 291443 471958
rect 582649 471474 582715 471477
rect 583520 471474 584960 471564
rect 582649 471472 584960 471474
rect 582649 471416 582654 471472
rect 582710 471416 584960 471472
rect 582649 471414 584960 471416
rect 582649 471411 582715 471414
rect 583520 471324 584960 471414
rect 161289 471202 161355 471205
rect 170489 471202 170555 471205
rect 161289 471200 170555 471202
rect 161289 471144 161294 471200
rect 161350 471144 170494 471200
rect 170550 471144 170555 471200
rect 161289 471142 170555 471144
rect 161289 471139 161355 471142
rect 170489 471139 170555 471142
rect 170857 471202 170923 471205
rect 206369 471202 206435 471205
rect 170857 471200 206435 471202
rect 170857 471144 170862 471200
rect 170918 471144 206374 471200
rect 206430 471144 206435 471200
rect 170857 471142 206435 471144
rect 170857 471139 170923 471142
rect 206369 471139 206435 471142
rect 209037 471202 209103 471205
rect 253933 471202 253999 471205
rect 209037 471200 253999 471202
rect 209037 471144 209042 471200
rect 209098 471144 253938 471200
rect 253994 471144 253999 471200
rect 209037 471142 253999 471144
rect 209037 471139 209103 471142
rect 209730 470661 209790 471142
rect 253933 471139 253999 471142
rect 209730 470656 209839 470661
rect 209730 470600 209778 470656
rect 209834 470600 209839 470656
rect 209730 470598 209839 470600
rect 209773 470595 209839 470598
rect 67725 469842 67791 469845
rect 91318 469842 91324 469844
rect 67725 469840 91324 469842
rect 67725 469784 67730 469840
rect 67786 469784 91324 469840
rect 67725 469782 91324 469784
rect 67725 469779 67791 469782
rect 91318 469780 91324 469782
rect 91388 469780 91394 469844
rect 165470 469780 165476 469844
rect 165540 469842 165546 469844
rect 228357 469842 228423 469845
rect 165540 469840 228423 469842
rect 165540 469784 228362 469840
rect 228418 469784 228423 469840
rect 165540 469782 228423 469784
rect 165540 469780 165546 469782
rect 228357 469779 228423 469782
rect 90357 469298 90423 469301
rect 91001 469298 91067 469301
rect 182909 469298 182975 469301
rect 90357 469296 182975 469298
rect 90357 469240 90362 469296
rect 90418 469240 91006 469296
rect 91062 469240 182914 469296
rect 182970 469240 182975 469296
rect 90357 469238 182975 469240
rect 90357 469235 90423 469238
rect 91001 469235 91067 469238
rect 182909 469235 182975 469238
rect 189717 469298 189783 469301
rect 278957 469298 279023 469301
rect 189717 469296 279023 469298
rect 189717 469240 189722 469296
rect 189778 469240 278962 469296
rect 279018 469240 279023 469296
rect 189717 469238 279023 469240
rect 189717 469235 189783 469238
rect 278957 469235 279023 469238
rect 173750 468556 173756 468620
rect 173820 468618 173826 468620
rect 184197 468618 184263 468621
rect 173820 468616 184263 468618
rect 173820 468560 184202 468616
rect 184258 468560 184263 468616
rect 173820 468558 184263 468560
rect 173820 468556 173826 468558
rect 184197 468555 184263 468558
rect 187141 468618 187207 468621
rect 196617 468618 196683 468621
rect 187141 468616 196683 468618
rect 187141 468560 187146 468616
rect 187202 468560 196622 468616
rect 196678 468560 196683 468616
rect 187141 468558 196683 468560
rect 187141 468555 187207 468558
rect 196617 468555 196683 468558
rect 115289 468482 115355 468485
rect 276013 468482 276079 468485
rect 115289 468480 276079 468482
rect 115289 468424 115294 468480
rect 115350 468424 276018 468480
rect 276074 468424 276079 468480
rect 115289 468422 276079 468424
rect 115289 468419 115355 468422
rect 276013 468419 276079 468422
rect 180006 467740 180012 467804
rect 180076 467802 180082 467804
rect 183001 467802 183067 467805
rect 180076 467800 183067 467802
rect 180076 467744 183006 467800
rect 183062 467744 183067 467800
rect 180076 467742 183067 467744
rect 180076 467740 180082 467742
rect 183001 467739 183067 467742
rect 186814 467196 186820 467260
rect 186884 467258 186890 467260
rect 203609 467258 203675 467261
rect 186884 467256 203675 467258
rect 186884 467200 203614 467256
rect 203670 467200 203675 467256
rect 186884 467198 203675 467200
rect 186884 467196 186890 467198
rect 203609 467195 203675 467198
rect 174670 467060 174676 467124
rect 174740 467122 174746 467124
rect 231209 467122 231275 467125
rect 174740 467120 231275 467122
rect 174740 467064 231214 467120
rect 231270 467064 231275 467120
rect 174740 467062 231275 467064
rect 174740 467060 174746 467062
rect 231209 467059 231275 467062
rect 255497 466714 255563 466717
rect 256550 466714 256556 466716
rect 255497 466712 256556 466714
rect 255497 466656 255502 466712
rect 255558 466656 256556 466712
rect 255497 466654 256556 466656
rect 255497 466651 255563 466654
rect 256550 466652 256556 466654
rect 256620 466652 256626 466716
rect 251081 466578 251147 466581
rect 285673 466580 285739 466581
rect 285622 466578 285628 466580
rect 251081 466576 285628 466578
rect 285692 466578 285739 466580
rect 285692 466576 285784 466578
rect 251081 466520 251086 466576
rect 251142 466520 285628 466576
rect 285734 466520 285784 466576
rect 251081 466518 285628 466520
rect 251081 466515 251147 466518
rect 285622 466516 285628 466518
rect 285692 466518 285784 466520
rect 285692 466516 285739 466518
rect 285673 466515 285739 466516
rect 246246 465972 246252 466036
rect 246316 466034 246322 466036
rect 269389 466034 269455 466037
rect 246316 466032 269455 466034
rect 246316 465976 269394 466032
rect 269450 465976 269455 466032
rect 246316 465974 269455 465976
rect 246316 465972 246322 465974
rect 269389 465971 269455 465974
rect 202781 465898 202847 465901
rect 251081 465898 251147 465901
rect 202781 465896 251147 465898
rect 202781 465840 202786 465896
rect 202842 465840 251086 465896
rect 251142 465840 251147 465896
rect 202781 465838 251147 465840
rect 202781 465835 202847 465838
rect 251081 465835 251147 465838
rect 169661 465762 169727 465765
rect 170949 465762 171015 465765
rect 255497 465762 255563 465765
rect 169661 465760 255563 465762
rect 169661 465704 169666 465760
rect 169722 465704 170954 465760
rect 171010 465704 255502 465760
rect 255558 465704 255563 465760
rect 169661 465702 255563 465704
rect 169661 465699 169727 465702
rect 170949 465699 171015 465702
rect 255497 465699 255563 465702
rect 273345 465082 273411 465085
rect 273478 465082 273484 465084
rect 273345 465080 273484 465082
rect 273345 465024 273350 465080
rect 273406 465024 273484 465080
rect 273345 465022 273484 465024
rect 273345 465019 273411 465022
rect 273478 465020 273484 465022
rect 273548 465020 273554 465084
rect 209865 464674 209931 464677
rect 227805 464674 227871 464677
rect 209865 464672 227871 464674
rect 209865 464616 209870 464672
rect 209926 464616 227810 464672
rect 227866 464616 227871 464672
rect 209865 464614 227871 464616
rect 209865 464611 209931 464614
rect 227805 464611 227871 464614
rect 181437 464538 181503 464541
rect 214557 464538 214623 464541
rect 181437 464536 214623 464538
rect 181437 464480 181442 464536
rect 181498 464480 214562 464536
rect 214618 464480 214623 464536
rect 181437 464478 214623 464480
rect 181437 464475 181503 464478
rect 214557 464475 214623 464478
rect 169334 464340 169340 464404
rect 169404 464402 169410 464404
rect 213913 464402 213979 464405
rect 169404 464400 213979 464402
rect 169404 464344 213918 464400
rect 213974 464344 213979 464400
rect 169404 464342 213979 464344
rect 169404 464340 169410 464342
rect 213913 464339 213979 464342
rect 213913 463722 213979 463725
rect 288525 463722 288591 463725
rect 213913 463720 288591 463722
rect 213913 463664 213918 463720
rect 213974 463664 288530 463720
rect 288586 463664 288591 463720
rect 213913 463662 288591 463664
rect 213913 463659 213979 463662
rect 288525 463659 288591 463662
rect 82670 463524 82676 463588
rect 82740 463586 82746 463588
rect 83958 463586 83964 463588
rect 82740 463526 83964 463586
rect 82740 463524 82746 463526
rect 83958 463524 83964 463526
rect 84028 463524 84034 463588
rect 171777 462906 171843 462909
rect 211654 462906 211660 462908
rect 171777 462904 211660 462906
rect 171777 462848 171782 462904
rect 171838 462848 211660 462904
rect 171777 462846 211660 462848
rect 171777 462843 171843 462846
rect 211654 462844 211660 462846
rect 211724 462844 211730 462908
rect 235993 462906 236059 462909
rect 244273 462906 244339 462909
rect 285673 462906 285739 462909
rect 235993 462904 285739 462906
rect 235993 462848 235998 462904
rect 236054 462848 244278 462904
rect 244334 462848 285678 462904
rect 285734 462848 285739 462904
rect 235993 462846 285739 462848
rect 235993 462843 236059 462846
rect 244273 462843 244339 462846
rect 285673 462843 285739 462846
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 98729 462362 98795 462365
rect 201493 462362 201559 462365
rect 202781 462362 202847 462365
rect 98729 462360 202847 462362
rect 98729 462304 98734 462360
rect 98790 462304 201498 462360
rect 201554 462304 202786 462360
rect 202842 462304 202847 462360
rect 98729 462302 202847 462304
rect 98729 462299 98795 462302
rect 201493 462299 201559 462302
rect 202781 462299 202847 462302
rect 193121 461682 193187 461685
rect 215385 461682 215451 461685
rect 193121 461680 215451 461682
rect 193121 461624 193126 461680
rect 193182 461624 215390 461680
rect 215446 461624 215451 461680
rect 193121 461622 215451 461624
rect 193121 461619 193187 461622
rect 215385 461619 215451 461622
rect 170806 461484 170812 461548
rect 170876 461546 170882 461548
rect 204897 461546 204963 461549
rect 170876 461544 204963 461546
rect 170876 461488 204902 461544
rect 204958 461488 204963 461544
rect 170876 461486 204963 461488
rect 170876 461484 170882 461486
rect 204897 461483 204963 461486
rect 117313 461002 117379 461005
rect 263777 461002 263843 461005
rect 117313 461000 263843 461002
rect 117313 460944 117318 461000
rect 117374 460944 263782 461000
rect 263838 460944 263843 461000
rect 117313 460942 263843 460944
rect 117313 460939 117379 460942
rect 263777 460939 263843 460942
rect 188337 460322 188403 460325
rect 208393 460322 208459 460325
rect 188337 460320 208459 460322
rect 188337 460264 188342 460320
rect 188398 460264 208398 460320
rect 208454 460264 208459 460320
rect 188337 460262 208459 460264
rect 188337 460259 188403 460262
rect 208393 460259 208459 460262
rect 215385 460322 215451 460325
rect 223982 460322 223988 460324
rect 215385 460320 223988 460322
rect 215385 460264 215390 460320
rect 215446 460264 223988 460320
rect 215385 460262 223988 460264
rect 215385 460259 215451 460262
rect 223982 460260 223988 460262
rect 224052 460260 224058 460324
rect 240777 460322 240843 460325
rect 255589 460322 255655 460325
rect 240777 460320 255655 460322
rect 240777 460264 240782 460320
rect 240838 460264 255594 460320
rect 255650 460264 255655 460320
rect 240777 460262 255655 460264
rect 240777 460259 240843 460262
rect 255589 460259 255655 460262
rect 166441 460186 166507 460189
rect 244917 460186 244983 460189
rect 166441 460184 244983 460186
rect 166441 460128 166446 460184
rect 166502 460128 244922 460184
rect 244978 460128 244983 460184
rect 166441 460126 244983 460128
rect 166441 460123 166507 460126
rect 244917 460123 244983 460126
rect 231117 459642 231183 459645
rect 289813 459642 289879 459645
rect 231117 459640 289879 459642
rect 231117 459584 231122 459640
rect 231178 459584 289818 459640
rect 289874 459584 289879 459640
rect 231117 459582 289879 459584
rect 231117 459579 231183 459582
rect 289813 459579 289879 459582
rect 201401 458962 201467 458965
rect 233182 458962 233188 458964
rect 201401 458960 233188 458962
rect 201401 458904 201406 458960
rect 201462 458904 233188 458960
rect 201401 458902 233188 458904
rect 201401 458899 201467 458902
rect 233182 458900 233188 458902
rect 233252 458900 233258 458964
rect 80053 458826 80119 458829
rect 113214 458826 113220 458828
rect 80053 458824 113220 458826
rect 80053 458768 80058 458824
rect 80114 458768 113220 458824
rect 80053 458766 113220 458768
rect 80053 458763 80119 458766
rect 113214 458764 113220 458766
rect 113284 458764 113290 458828
rect 135161 458826 135227 458829
rect 184657 458826 184723 458829
rect 135161 458824 184723 458826
rect 135161 458768 135166 458824
rect 135222 458768 184662 458824
rect 184718 458768 184723 458824
rect 135161 458766 184723 458768
rect 135161 458763 135227 458766
rect 184657 458763 184723 458766
rect 191649 458826 191715 458829
rect 228214 458826 228220 458828
rect 191649 458824 228220 458826
rect 191649 458768 191654 458824
rect 191710 458768 228220 458824
rect 191649 458766 228220 458768
rect 191649 458763 191715 458766
rect 228214 458764 228220 458766
rect 228284 458764 228290 458828
rect 187601 458554 187667 458557
rect 259637 458554 259703 458557
rect 187601 458552 259703 458554
rect 187601 458496 187606 458552
rect 187662 458496 259642 458552
rect 259698 458496 259703 458552
rect 187601 458494 259703 458496
rect 187601 458491 187667 458494
rect 259637 458491 259703 458494
rect 232129 458418 232195 458421
rect 276289 458418 276355 458421
rect 232129 458416 276355 458418
rect 232129 458360 232134 458416
rect 232190 458360 276294 458416
rect 276350 458360 276355 458416
rect 232129 458358 276355 458360
rect 232129 458355 232195 458358
rect 276289 458355 276355 458358
rect 184790 458220 184796 458284
rect 184860 458282 184866 458284
rect 187785 458282 187851 458285
rect 184860 458280 187851 458282
rect 184860 458224 187790 458280
rect 187846 458224 187851 458280
rect 184860 458222 187851 458224
rect 184860 458220 184866 458222
rect 187785 458219 187851 458222
rect 148910 458084 148916 458148
rect 148980 458146 148986 458148
rect 153929 458146 153995 458149
rect 148980 458144 153995 458146
rect 148980 458088 153934 458144
rect 153990 458088 153995 458144
rect 148980 458086 153995 458088
rect 148980 458084 148986 458086
rect 153929 458083 153995 458086
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 172329 457602 172395 457605
rect 202965 457602 203031 457605
rect 172329 457600 203031 457602
rect 172329 457544 172334 457600
rect 172390 457544 202970 457600
rect 203026 457544 203031 457600
rect 172329 457542 203031 457544
rect 172329 457539 172395 457542
rect 202965 457539 203031 457542
rect 81341 457466 81407 457469
rect 96838 457466 96844 457468
rect 81341 457464 96844 457466
rect 81341 457408 81346 457464
rect 81402 457408 96844 457464
rect 81341 457406 96844 457408
rect 81341 457403 81407 457406
rect 96838 457404 96844 457406
rect 96908 457404 96914 457468
rect 164141 457466 164207 457469
rect 206461 457466 206527 457469
rect 164141 457464 206527 457466
rect 164141 457408 164146 457464
rect 164202 457408 206466 457464
rect 206522 457408 206527 457464
rect 164141 457406 206527 457408
rect 164141 457403 164207 457406
rect 206461 457403 206527 457406
rect 223665 457466 223731 457469
rect 284334 457466 284340 457468
rect 223665 457464 284340 457466
rect 223665 457408 223670 457464
rect 223726 457408 284340 457464
rect 223665 457406 284340 457408
rect 223665 457403 223731 457406
rect 284334 457404 284340 457406
rect 284404 457404 284410 457468
rect 52361 456922 52427 456925
rect 150934 456922 150940 456924
rect 52361 456920 150940 456922
rect 52361 456864 52366 456920
rect 52422 456864 150940 456920
rect 52361 456862 150940 456864
rect 52361 456859 52427 456862
rect 150934 456860 150940 456862
rect 151004 456860 151010 456924
rect 190361 456922 190427 456925
rect 219433 456922 219499 456925
rect 219801 456922 219867 456925
rect 190361 456920 219867 456922
rect 190361 456864 190366 456920
rect 190422 456864 219438 456920
rect 219494 456864 219806 456920
rect 219862 456864 219867 456920
rect 190361 456862 219867 456864
rect 190361 456859 190427 456862
rect 219433 456859 219499 456862
rect 219801 456859 219867 456862
rect 223481 456922 223547 456925
rect 223665 456922 223731 456925
rect 223481 456920 223731 456922
rect 223481 456864 223486 456920
rect 223542 456864 223670 456920
rect 223726 456864 223731 456920
rect 223481 456862 223731 456864
rect 223481 456859 223547 456862
rect 223665 456859 223731 456862
rect 241421 456922 241487 456925
rect 281809 456922 281875 456925
rect 241421 456920 281875 456922
rect 241421 456864 241426 456920
rect 241482 456864 281814 456920
rect 281870 456864 281875 456920
rect 241421 456862 281875 456864
rect 241421 456859 241487 456862
rect 281809 456859 281875 456862
rect 168966 456180 168972 456244
rect 169036 456242 169042 456244
rect 200205 456242 200271 456245
rect 169036 456240 200271 456242
rect 169036 456184 200210 456240
rect 200266 456184 200271 456240
rect 169036 456182 200271 456184
rect 169036 456180 169042 456182
rect 200205 456179 200271 456182
rect 106774 456044 106780 456108
rect 106844 456106 106850 456108
rect 153837 456106 153903 456109
rect 106844 456104 153903 456106
rect 106844 456048 153842 456104
rect 153898 456048 153903 456104
rect 106844 456046 153903 456048
rect 106844 456044 106850 456046
rect 153837 456043 153903 456046
rect 191465 456106 191531 456109
rect 247718 456106 247724 456108
rect 191465 456104 247724 456106
rect 191465 456048 191470 456104
rect 191526 456048 247724 456104
rect 191465 456046 247724 456048
rect 191465 456043 191531 456046
rect 247718 456044 247724 456046
rect 247788 456044 247794 456108
rect 249057 456106 249123 456109
rect 284477 456106 284543 456109
rect 249057 456104 284543 456106
rect 249057 456048 249062 456104
rect 249118 456048 284482 456104
rect 284538 456048 284543 456104
rect 249057 456046 284543 456048
rect 249057 456043 249123 456046
rect 284477 456043 284543 456046
rect 230565 455970 230631 455973
rect 231301 455970 231367 455973
rect 230565 455968 231367 455970
rect 230565 455912 230570 455968
rect 230626 455912 231306 455968
rect 231362 455912 231367 455968
rect 230565 455910 231367 455912
rect 230565 455907 230631 455910
rect 231301 455907 231367 455910
rect 150157 455562 150223 455565
rect 215385 455562 215451 455565
rect 150157 455560 215451 455562
rect 150157 455504 150162 455560
rect 150218 455504 215390 455560
rect 215446 455504 215451 455560
rect 150157 455502 215451 455504
rect 150157 455499 150223 455502
rect 215385 455499 215451 455502
rect 231301 455562 231367 455565
rect 287329 455562 287395 455565
rect 288341 455562 288407 455565
rect 231301 455560 288407 455562
rect 231301 455504 231306 455560
rect 231362 455504 287334 455560
rect 287390 455504 288346 455560
rect 288402 455504 288407 455560
rect 231301 455502 288407 455504
rect 231301 455499 231367 455502
rect 287329 455499 287395 455502
rect 288341 455499 288407 455502
rect 182909 454882 182975 454885
rect 193397 454882 193463 454885
rect 182909 454880 193463 454882
rect 182909 454824 182914 454880
rect 182970 454824 193402 454880
rect 193458 454824 193463 454880
rect 182909 454822 193463 454824
rect 182909 454819 182975 454822
rect 193397 454819 193463 454822
rect 179086 454684 179092 454748
rect 179156 454746 179162 454748
rect 202137 454746 202203 454749
rect 179156 454744 202203 454746
rect 179156 454688 202142 454744
rect 202198 454688 202203 454744
rect 179156 454686 202203 454688
rect 179156 454684 179162 454686
rect 202137 454683 202203 454686
rect 212625 454746 212691 454749
rect 222193 454746 222259 454749
rect 287237 454746 287303 454749
rect 212625 454744 287303 454746
rect 212625 454688 212630 454744
rect 212686 454688 222198 454744
rect 222254 454688 287242 454744
rect 287298 454688 287303 454744
rect 212625 454686 287303 454688
rect 212625 454683 212691 454686
rect 222193 454683 222259 454686
rect 287237 454683 287303 454686
rect 112989 454068 113055 454069
rect 112989 454064 113036 454068
rect 113100 454066 113106 454068
rect 112989 454008 112994 454064
rect 112989 454004 113036 454008
rect 113100 454006 113146 454066
rect 113100 454004 113106 454006
rect 147438 454004 147444 454068
rect 147508 454066 147514 454068
rect 197905 454066 197971 454069
rect 147508 454064 197971 454066
rect 147508 454008 197910 454064
rect 197966 454008 197971 454064
rect 147508 454006 197971 454008
rect 147508 454004 147514 454006
rect 112989 454003 113055 454004
rect 197905 454003 197971 454006
rect 202965 454066 203031 454069
rect 222101 454066 222167 454069
rect 202965 454064 222167 454066
rect 202965 454008 202970 454064
rect 203026 454008 222106 454064
rect 222162 454008 222167 454064
rect 202965 454006 222167 454008
rect 202965 454003 203031 454006
rect 222101 454003 222167 454006
rect 234889 454066 234955 454069
rect 235901 454066 235967 454069
rect 257337 454066 257403 454069
rect 234889 454064 257403 454066
rect 234889 454008 234894 454064
rect 234950 454008 235906 454064
rect 235962 454008 257342 454064
rect 257398 454008 257403 454064
rect 234889 454006 257403 454008
rect 234889 454003 234955 454006
rect 235901 454003 235967 454006
rect 257337 454003 257403 454006
rect 232497 453930 232563 453933
rect 233509 453930 233575 453933
rect 232497 453928 233575 453930
rect 232497 453872 232502 453928
rect 232558 453872 233514 453928
rect 233570 453872 233575 453928
rect 232497 453870 233575 453872
rect 232497 453867 232563 453870
rect 233509 453867 233575 453870
rect 239397 453930 239463 453933
rect 241646 453930 241652 453932
rect 239397 453928 241652 453930
rect 239397 453872 239402 453928
rect 239458 453872 241652 453928
rect 239397 453870 241652 453872
rect 239397 453867 239463 453870
rect 241646 453868 241652 453870
rect 241716 453868 241722 453932
rect 166441 453250 166507 453253
rect 198825 453250 198891 453253
rect 166441 453248 198891 453250
rect 166441 453192 166446 453248
rect 166502 453192 198830 453248
rect 198886 453192 198891 453248
rect 166441 453190 198891 453192
rect 166441 453187 166507 453190
rect 198825 453187 198891 453190
rect 222101 453250 222167 453253
rect 296805 453250 296871 453253
rect 222101 453248 296871 453250
rect 222101 453192 222106 453248
rect 222162 453192 296810 453248
rect 296866 453192 296871 453248
rect 222101 453190 296871 453192
rect 222101 453187 222167 453190
rect 296805 453187 296871 453190
rect 242157 452842 242223 452845
rect 262305 452842 262371 452845
rect 242157 452840 262371 452842
rect 242157 452784 242162 452840
rect 242218 452784 262310 452840
rect 262366 452784 262371 452840
rect 242157 452782 262371 452784
rect 242157 452779 242223 452782
rect 262305 452779 262371 452782
rect 74441 452706 74507 452709
rect 200849 452706 200915 452709
rect 201401 452706 201467 452709
rect 74441 452704 201467 452706
rect 74441 452648 74446 452704
rect 74502 452648 200854 452704
rect 200910 452648 201406 452704
rect 201462 452648 201467 452704
rect 74441 452646 201467 452648
rect 74441 452643 74507 452646
rect 200849 452643 200915 452646
rect 201401 452643 201467 452646
rect 244917 452706 244983 452709
rect 277158 452706 277164 452708
rect 244917 452704 277164 452706
rect 244917 452648 244922 452704
rect 244978 452648 277164 452704
rect 244917 452646 277164 452648
rect 244917 452643 244983 452646
rect 277158 452644 277164 452646
rect 277228 452644 277234 452708
rect 193305 452570 193371 452573
rect 197445 452570 197511 452573
rect 193305 452568 197511 452570
rect 193305 452512 193310 452568
rect 193366 452512 197450 452568
rect 197506 452512 197511 452568
rect 193305 452510 197511 452512
rect 193305 452507 193371 452510
rect 197445 452507 197511 452510
rect 250437 452162 250503 452165
rect 253974 452162 253980 452164
rect 250437 452160 253980 452162
rect 250437 452104 250442 452160
rect 250498 452104 253980 452160
rect 250437 452102 253980 452104
rect 250437 452099 250503 452102
rect 253974 452100 253980 452102
rect 254044 452100 254050 452164
rect 98637 451890 98703 451893
rect 122741 451890 122807 451893
rect 98637 451888 122807 451890
rect 98637 451832 98642 451888
rect 98698 451832 122746 451888
rect 122802 451832 122807 451888
rect 98637 451830 122807 451832
rect 98637 451827 98703 451830
rect 122741 451827 122807 451830
rect 158805 451890 158871 451893
rect 159909 451890 159975 451893
rect 239213 451890 239279 451893
rect 158805 451888 239279 451890
rect 158805 451832 158810 451888
rect 158866 451832 159914 451888
rect 159970 451832 239218 451888
rect 239274 451832 239279 451888
rect 158805 451830 239279 451832
rect 158805 451827 158871 451830
rect 159909 451827 159975 451830
rect 239213 451827 239279 451830
rect 233509 451482 233575 451485
rect 251909 451482 251975 451485
rect 233509 451480 251975 451482
rect 233509 451424 233514 451480
rect 233570 451424 251914 451480
rect 251970 451424 251975 451480
rect 233509 451422 251975 451424
rect 233509 451419 233575 451422
rect 251909 451419 251975 451422
rect 122741 451346 122807 451349
rect 122925 451346 122991 451349
rect 122741 451344 122991 451346
rect 122741 451288 122746 451344
rect 122802 451288 122930 451344
rect 122986 451288 122991 451344
rect 122741 451286 122991 451288
rect 122741 451283 122807 451286
rect 122925 451283 122991 451286
rect 239213 451346 239279 451349
rect 270585 451346 270651 451349
rect 239213 451344 270651 451346
rect 239213 451288 239218 451344
rect 239274 451288 270590 451344
rect 270646 451288 270651 451344
rect 239213 451286 270651 451288
rect 239213 451283 239279 451286
rect 270585 451283 270651 451286
rect 202873 450530 202939 450533
rect 204069 450530 204135 450533
rect 202873 450528 204135 450530
rect 202873 450472 202878 450528
rect 202934 450472 204074 450528
rect 204130 450472 204135 450528
rect 202873 450470 204135 450472
rect 202873 450467 202939 450470
rect 204069 450467 204135 450470
rect 192661 450394 192727 450397
rect 197537 450394 197603 450397
rect 192661 450392 197603 450394
rect 192661 450336 192666 450392
rect 192722 450336 197542 450392
rect 197598 450336 197603 450392
rect 192661 450334 197603 450336
rect 192661 450331 192727 450334
rect 197537 450331 197603 450334
rect 174997 450258 175063 450261
rect 207289 450258 207355 450261
rect 207565 450258 207631 450261
rect 245929 450260 245995 450261
rect 174997 450256 207631 450258
rect 174997 450200 175002 450256
rect 175058 450200 207294 450256
rect 207350 450200 207570 450256
rect 207626 450200 207631 450256
rect 174997 450198 207631 450200
rect 174997 450195 175063 450198
rect 207289 450195 207355 450198
rect 207565 450195 207631 450198
rect 245878 450196 245884 450260
rect 245948 450258 245995 450260
rect 245948 450256 246040 450258
rect 245990 450200 246040 450256
rect 245948 450198 246040 450200
rect 245948 450196 245995 450198
rect 245929 450195 245995 450196
rect 151629 450122 151695 450125
rect 205633 450122 205699 450125
rect 151629 450120 205699 450122
rect 151629 450064 151634 450120
rect 151690 450064 205638 450120
rect 205694 450064 205699 450120
rect 151629 450062 205699 450064
rect 151629 450059 151695 450062
rect 205633 450059 205699 450062
rect 228817 450122 228883 450125
rect 283097 450122 283163 450125
rect 228817 450120 283163 450122
rect 228817 450064 228822 450120
rect 228878 450064 283102 450120
rect 283158 450064 283163 450120
rect 228817 450062 283163 450064
rect 228817 450059 228883 450062
rect 283097 450059 283163 450062
rect 204161 449986 204227 449989
rect 273621 449986 273687 449989
rect 204161 449984 273687 449986
rect 204161 449928 204166 449984
rect 204222 449928 273626 449984
rect 273682 449928 273687 449984
rect 204161 449926 273687 449928
rect 204161 449923 204227 449926
rect 273621 449923 273687 449926
rect -960 449578 480 449668
rect 245694 449652 245700 449716
rect 245764 449714 245770 449716
rect 246113 449714 246179 449717
rect 245764 449712 246179 449714
rect 245764 449656 246118 449712
rect 246174 449656 246179 449712
rect 245764 449654 246179 449656
rect 245764 449652 245770 449654
rect 246113 449651 246179 449654
rect 247125 449714 247191 449717
rect 247718 449714 247724 449716
rect 247125 449712 247724 449714
rect 247125 449656 247130 449712
rect 247186 449656 247724 449712
rect 247125 449654 247724 449656
rect 247125 449651 247191 449654
rect 247718 449652 247724 449654
rect 247788 449652 247794 449716
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 186129 449442 186195 449445
rect 193213 449442 193279 449445
rect 186129 449440 193279 449442
rect 186129 449384 186134 449440
rect 186190 449384 193218 449440
rect 193274 449384 193279 449440
rect 186129 449382 193279 449384
rect 186129 449379 186195 449382
rect 193213 449379 193279 449382
rect 144637 449170 144703 449173
rect 184841 449170 184907 449173
rect 144637 449168 184907 449170
rect 144637 449112 144642 449168
rect 144698 449112 184846 449168
rect 184902 449112 184907 449168
rect 144637 449110 184907 449112
rect 144637 449107 144703 449110
rect 184841 449107 184907 449110
rect 191557 449170 191623 449173
rect 191557 449168 193660 449170
rect 191557 449112 191562 449168
rect 191618 449112 193660 449168
rect 191557 449110 193660 449112
rect 191557 449107 191623 449110
rect 255589 448898 255655 448901
rect 253460 448896 255655 448898
rect 253460 448840 255594 448896
rect 255650 448840 255655 448896
rect 253460 448838 255655 448840
rect 255589 448835 255655 448838
rect 192753 448628 192819 448629
rect 192702 448626 192708 448628
rect 192662 448566 192708 448626
rect 192772 448624 192819 448628
rect 192814 448568 192819 448624
rect 192702 448564 192708 448566
rect 192772 448564 192819 448568
rect 192753 448563 192819 448564
rect 69657 448490 69723 448493
rect 182173 448490 182239 448493
rect 69657 448488 182239 448490
rect 69657 448432 69662 448488
rect 69718 448432 182178 448488
rect 182234 448432 182239 448488
rect 69657 448430 182239 448432
rect 69657 448427 69723 448430
rect 182173 448427 182239 448430
rect 253565 448082 253631 448085
rect 253430 448080 253631 448082
rect 253430 448024 253570 448080
rect 253626 448024 253631 448080
rect 253430 448022 253631 448024
rect 191557 447810 191623 447813
rect 191557 447808 193660 447810
rect 191557 447752 191562 447808
rect 191618 447752 193660 447808
rect 191557 447750 193660 447752
rect 191557 447747 191623 447750
rect 253430 447538 253490 448022
rect 253565 448019 253631 448022
rect 255589 447810 255655 447813
rect 271086 447810 271092 447812
rect 255589 447808 271092 447810
rect 255589 447752 255594 447808
rect 255650 447752 271092 447808
rect 255589 447750 271092 447752
rect 255589 447747 255655 447750
rect 271086 447748 271092 447750
rect 271156 447748 271162 447812
rect 255589 447538 255655 447541
rect 253430 447536 255655 447538
rect 253430 447508 255594 447536
rect 253460 447480 255594 447508
rect 255650 447480 255655 447536
rect 253460 447478 255655 447480
rect 255589 447475 255655 447478
rect 188838 447340 188844 447404
rect 188908 447402 188914 447404
rect 192661 447402 192727 447405
rect 188908 447400 192727 447402
rect 188908 447344 192666 447400
rect 192722 447344 192727 447400
rect 188908 447342 192727 447344
rect 188908 447340 188914 447342
rect 192661 447339 192727 447342
rect 187601 446450 187667 446453
rect 188286 446450 188292 446452
rect 187601 446448 188292 446450
rect 187601 446392 187606 446448
rect 187662 446392 188292 446448
rect 187601 446390 188292 446392
rect 187601 446387 187667 446390
rect 188286 446388 188292 446390
rect 188356 446388 188362 446452
rect 191005 446450 191071 446453
rect 191005 446448 193660 446450
rect 191005 446392 191010 446448
rect 191066 446392 193660 446448
rect 191005 446390 193660 446392
rect 191005 446387 191071 446390
rect 253974 446178 253980 446180
rect 253460 446118 253980 446178
rect 253974 446116 253980 446118
rect 254044 446178 254050 446180
rect 255957 446178 256023 446181
rect 254044 446176 256023 446178
rect 254044 446120 255962 446176
rect 256018 446120 256023 446176
rect 254044 446118 256023 446120
rect 254044 446116 254050 446118
rect 255957 446115 256023 446118
rect 191005 445090 191071 445093
rect 191005 445088 193660 445090
rect 191005 445032 191010 445088
rect 191066 445032 193660 445088
rect 191005 445030 193660 445032
rect 191005 445027 191071 445030
rect 66662 444892 66668 444956
rect 66732 444954 66738 444956
rect 95325 444954 95391 444957
rect 66732 444952 95391 444954
rect 66732 444896 95330 444952
rect 95386 444896 95391 444952
rect 66732 444894 95391 444896
rect 66732 444892 66738 444894
rect 95325 444891 95391 444894
rect 255497 444818 255563 444821
rect 253460 444816 255563 444818
rect 253460 444760 255502 444816
rect 255558 444760 255563 444816
rect 253460 444758 255563 444760
rect 255497 444755 255563 444758
rect 583520 444668 584960 444908
rect 193029 443730 193095 443733
rect 193029 443728 193660 443730
rect 193029 443672 193034 443728
rect 193090 443672 193660 443728
rect 193029 443670 193660 443672
rect 193029 443667 193095 443670
rect 255497 443458 255563 443461
rect 253460 443456 255563 443458
rect 253460 443400 255502 443456
rect 255558 443400 255563 443456
rect 253460 443398 255563 443400
rect 255497 443395 255563 443398
rect 60641 443050 60707 443053
rect 76557 443050 76623 443053
rect 60641 443048 76623 443050
rect 60641 442992 60646 443048
rect 60702 442992 76562 443048
rect 76618 442992 76623 443048
rect 60641 442990 76623 442992
rect 60641 442987 60707 442990
rect 76557 442987 76623 442990
rect 159909 443050 159975 443053
rect 163589 443050 163655 443053
rect 159909 443048 163655 443050
rect 159909 442992 159914 443048
rect 159970 442992 163594 443048
rect 163650 442992 163655 443048
rect 159909 442990 163655 442992
rect 159909 442987 159975 442990
rect 163589 442987 163655 442990
rect 191557 442098 191623 442101
rect 255497 442098 255563 442101
rect 191557 442096 193660 442098
rect 191557 442040 191562 442096
rect 191618 442040 193660 442096
rect 191557 442038 193660 442040
rect 253460 442096 255563 442098
rect 253460 442040 255502 442096
rect 255558 442040 255563 442096
rect 253460 442038 255563 442040
rect 191557 442035 191623 442038
rect 255497 442035 255563 442038
rect 69422 440812 69428 440876
rect 69492 440874 69498 440876
rect 173617 440874 173683 440877
rect 69492 440872 173683 440874
rect 69492 440816 173622 440872
rect 173678 440816 173683 440872
rect 69492 440814 173683 440816
rect 69492 440812 69498 440814
rect 173617 440811 173683 440814
rect 191557 440738 191623 440741
rect 191557 440736 193660 440738
rect 191557 440680 191562 440736
rect 191618 440680 193660 440736
rect 191557 440678 193660 440680
rect 191557 440675 191623 440678
rect 254526 440466 254532 440468
rect 253460 440406 254532 440466
rect 254526 440404 254532 440406
rect 254596 440466 254602 440468
rect 256877 440466 256943 440469
rect 254596 440464 256943 440466
rect 254596 440408 256882 440464
rect 256938 440408 256943 440464
rect 254596 440406 256943 440408
rect 254596 440404 254602 440406
rect 256877 440403 256943 440406
rect 68134 439452 68140 439516
rect 68204 439514 68210 439516
rect 170765 439514 170831 439517
rect 68204 439512 171150 439514
rect 68204 439456 170770 439512
rect 170826 439456 171150 439512
rect 68204 439454 171150 439456
rect 68204 439452 68210 439454
rect 170765 439451 170831 439454
rect 70710 438908 70716 438972
rect 70780 438970 70786 438972
rect 71630 438970 71636 438972
rect 70780 438910 71636 438970
rect 70780 438908 70786 438910
rect 71630 438908 71636 438910
rect 71700 438970 71706 438972
rect 128997 438970 129063 438973
rect 71700 438968 129063 438970
rect 71700 438912 129002 438968
rect 129058 438912 129063 438968
rect 71700 438910 129063 438912
rect 171090 438970 171150 439454
rect 193630 438970 193690 439348
rect 255497 439106 255563 439109
rect 253460 439104 255563 439106
rect 253460 439048 255502 439104
rect 255558 439048 255563 439104
rect 253460 439046 255563 439048
rect 255497 439043 255563 439046
rect 171090 438910 193690 438970
rect 71700 438908 71706 438910
rect 128997 438907 129063 438910
rect 68921 438154 68987 438157
rect 90357 438154 90423 438157
rect 68921 438152 90423 438154
rect 68921 438096 68926 438152
rect 68982 438096 90362 438152
rect 90418 438096 90423 438152
rect 68921 438094 90423 438096
rect 68921 438091 68987 438094
rect 90357 438091 90423 438094
rect 191649 438018 191715 438021
rect 191649 438016 193660 438018
rect 191649 437960 191654 438016
rect 191710 437960 193660 438016
rect 191649 437958 193660 437960
rect 191649 437955 191715 437958
rect 255497 437746 255563 437749
rect 253460 437744 255563 437746
rect 253460 437688 255502 437744
rect 255558 437688 255563 437744
rect 253460 437686 255563 437688
rect 255497 437683 255563 437686
rect 42701 437610 42767 437613
rect 77385 437610 77451 437613
rect 79317 437610 79383 437613
rect 42701 437608 79383 437610
rect 42701 437552 42706 437608
rect 42762 437552 77390 437608
rect 77446 437552 79322 437608
rect 79378 437552 79383 437608
rect 42701 437550 79383 437552
rect 42701 437547 42767 437550
rect 77385 437547 77451 437550
rect 79317 437547 79383 437550
rect 255865 437610 255931 437613
rect 256550 437610 256556 437612
rect 255865 437608 256556 437610
rect 255865 437552 255870 437608
rect 255926 437552 256556 437608
rect 255865 437550 256556 437552
rect 255865 437547 255931 437550
rect 256550 437548 256556 437550
rect 256620 437610 256626 437612
rect 295333 437610 295399 437613
rect 256620 437608 295399 437610
rect 256620 437552 295338 437608
rect 295394 437552 295399 437608
rect 256620 437550 295399 437552
rect 256620 437548 256626 437550
rect 295333 437547 295399 437550
rect 89345 436794 89411 436797
rect 98637 436794 98703 436797
rect 89345 436792 98703 436794
rect -960 436508 480 436748
rect 89345 436736 89350 436792
rect 89406 436736 98642 436792
rect 98698 436736 98703 436792
rect 89345 436734 98703 436736
rect 89345 436731 89411 436734
rect 98637 436731 98703 436734
rect 191649 436658 191715 436661
rect 191649 436656 193660 436658
rect 191649 436600 191654 436656
rect 191710 436600 193660 436656
rect 191649 436598 193660 436600
rect 191649 436595 191715 436598
rect 73470 436324 73476 436388
rect 73540 436386 73546 436388
rect 80237 436386 80303 436389
rect 255865 436386 255931 436389
rect 73540 436384 80303 436386
rect 73540 436328 80242 436384
rect 80298 436328 80303 436384
rect 73540 436326 80303 436328
rect 253460 436384 255931 436386
rect 253460 436328 255870 436384
rect 255926 436328 255931 436384
rect 253460 436326 255931 436328
rect 73540 436324 73546 436326
rect 80237 436323 80303 436326
rect 255865 436323 255931 436326
rect 70485 436250 70551 436253
rect 70853 436250 70919 436253
rect 75177 436250 75243 436253
rect 70485 436248 75243 436250
rect 70485 436192 70490 436248
rect 70546 436192 70858 436248
rect 70914 436192 75182 436248
rect 75238 436192 75243 436248
rect 70485 436190 75243 436192
rect 70485 436187 70551 436190
rect 70853 436187 70919 436190
rect 75177 436187 75243 436190
rect 78254 436188 78260 436252
rect 78324 436250 78330 436252
rect 80053 436250 80119 436253
rect 78324 436248 80119 436250
rect 78324 436192 80058 436248
rect 80114 436192 80119 436248
rect 78324 436190 80119 436192
rect 78324 436188 78330 436190
rect 80053 436187 80119 436190
rect 102726 436188 102732 436252
rect 102796 436250 102802 436252
rect 107653 436250 107719 436253
rect 102796 436248 107719 436250
rect 102796 436192 107658 436248
rect 107714 436192 107719 436248
rect 102796 436190 107719 436192
rect 102796 436188 102802 436190
rect 107653 436187 107719 436190
rect 108941 436250 109007 436253
rect 118693 436250 118759 436253
rect 108941 436248 118759 436250
rect 108941 436192 108946 436248
rect 109002 436192 118698 436248
rect 118754 436192 118759 436248
rect 108941 436190 118759 436192
rect 108941 436187 109007 436190
rect 118693 436187 118759 436190
rect 79726 436052 79732 436116
rect 79796 436114 79802 436116
rect 82077 436114 82143 436117
rect 79796 436112 82143 436114
rect 79796 436056 82082 436112
rect 82138 436056 82143 436112
rect 79796 436054 82143 436056
rect 79796 436052 79802 436054
rect 82077 436051 82143 436054
rect 84694 436052 84700 436116
rect 84764 436114 84770 436116
rect 91093 436114 91159 436117
rect 84764 436112 91159 436114
rect 84764 436056 91098 436112
rect 91154 436056 91159 436112
rect 84764 436054 91159 436056
rect 84764 436052 84770 436054
rect 91093 436051 91159 436054
rect 94446 436052 94452 436116
rect 94516 436114 94522 436116
rect 96889 436114 96955 436117
rect 94516 436112 96955 436114
rect 94516 436056 96894 436112
rect 96950 436056 96955 436112
rect 94516 436054 96955 436056
rect 94516 436052 94522 436054
rect 96889 436051 96955 436054
rect 180517 435978 180583 435981
rect 182817 435978 182883 435981
rect 180517 435976 182883 435978
rect 180517 435920 180522 435976
rect 180578 435920 182822 435976
rect 182878 435920 182883 435976
rect 180517 435918 182883 435920
rect 180517 435915 180583 435918
rect 182817 435915 182883 435918
rect 191649 435298 191715 435301
rect 191649 435296 193660 435298
rect 191649 435240 191654 435296
rect 191710 435240 193660 435296
rect 191649 435238 193660 435240
rect 191649 435235 191715 435238
rect 255497 435026 255563 435029
rect 253460 435024 255563 435026
rect 253460 434968 255502 435024
rect 255558 434968 255563 435024
rect 253460 434966 255563 434968
rect 255497 434963 255563 434966
rect 72601 434890 72667 434893
rect 72601 434888 84210 434890
rect 72601 434832 72606 434888
rect 72662 434832 84210 434888
rect 72601 434830 84210 434832
rect 72601 434827 72667 434830
rect 53465 434754 53531 434757
rect 69841 434754 69907 434757
rect 53465 434752 69907 434754
rect 53465 434696 53470 434752
rect 53526 434696 69846 434752
rect 69902 434696 69907 434752
rect 53465 434694 69907 434696
rect 84150 434754 84210 434830
rect 132493 434754 132559 434757
rect 84150 434752 132559 434754
rect 84150 434696 132498 434752
rect 132554 434696 132559 434752
rect 84150 434694 132559 434696
rect 53465 434691 53531 434694
rect 69841 434691 69907 434694
rect 132493 434691 132559 434694
rect 66069 434618 66135 434621
rect 67398 434618 67404 434620
rect 66069 434616 67404 434618
rect 66069 434560 66074 434616
rect 66130 434560 67404 434616
rect 66069 434558 67404 434560
rect 66069 434555 66135 434558
rect 67398 434556 67404 434558
rect 67468 434556 67474 434620
rect 83038 434420 83044 434484
rect 83108 434482 83114 434484
rect 83733 434482 83799 434485
rect 83108 434480 83799 434482
rect 83108 434424 83738 434480
rect 83794 434424 83799 434480
rect 83108 434422 83799 434424
rect 83108 434420 83114 434422
rect 83733 434419 83799 434422
rect 69054 434284 69060 434348
rect 69124 434346 69130 434348
rect 69197 434346 69263 434349
rect 69124 434344 69263 434346
rect 69124 434288 69202 434344
rect 69258 434288 69263 434344
rect 69124 434286 69263 434288
rect 69124 434284 69130 434286
rect 69197 434283 69263 434286
rect 80094 434284 80100 434348
rect 80164 434346 80170 434348
rect 80973 434346 81039 434349
rect 84561 434348 84627 434349
rect 85849 434348 85915 434349
rect 84510 434346 84516 434348
rect 80164 434344 81039 434346
rect 80164 434288 80978 434344
rect 81034 434288 81039 434344
rect 80164 434286 81039 434288
rect 84470 434286 84516 434346
rect 84580 434344 84627 434348
rect 85798 434346 85804 434348
rect 84622 434288 84627 434344
rect 80164 434284 80170 434286
rect 80973 434283 81039 434286
rect 84510 434284 84516 434286
rect 84580 434284 84627 434288
rect 85758 434286 85804 434346
rect 85868 434344 85915 434348
rect 85910 434288 85915 434344
rect 85798 434284 85804 434286
rect 85868 434284 85915 434288
rect 95182 434284 95188 434348
rect 95252 434346 95258 434348
rect 95693 434346 95759 434349
rect 100201 434348 100267 434349
rect 100150 434346 100156 434348
rect 95252 434344 95759 434346
rect 95252 434288 95698 434344
rect 95754 434288 95759 434344
rect 95252 434286 95759 434288
rect 100110 434286 100156 434346
rect 100220 434344 100267 434348
rect 100262 434288 100267 434344
rect 95252 434284 95258 434286
rect 84561 434283 84627 434284
rect 85849 434283 85915 434284
rect 95693 434283 95759 434286
rect 100150 434284 100156 434286
rect 100220 434284 100267 434288
rect 100201 434283 100267 434284
rect 92657 434212 92723 434213
rect 92606 434210 92612 434212
rect 92566 434150 92612 434210
rect 92676 434208 92723 434212
rect 92718 434152 92723 434208
rect 92606 434148 92612 434150
rect 92676 434148 92723 434152
rect 92657 434147 92723 434148
rect 67398 433876 67404 433940
rect 67468 433938 67474 433940
rect 90633 433938 90699 433941
rect 67468 433936 90699 433938
rect 67468 433880 90638 433936
rect 90694 433880 90699 433936
rect 67468 433878 90699 433880
rect 67468 433876 67474 433878
rect 90633 433875 90699 433878
rect 74942 433740 74948 433804
rect 75012 433802 75018 433804
rect 75453 433802 75519 433805
rect 75012 433800 75519 433802
rect 75012 433744 75458 433800
rect 75514 433744 75519 433800
rect 75012 433742 75519 433744
rect 75012 433740 75018 433742
rect 75453 433739 75519 433742
rect 98494 433740 98500 433804
rect 98564 433802 98570 433804
rect 101213 433802 101279 433805
rect 98564 433800 101279 433802
rect 98564 433744 101218 433800
rect 101274 433744 101279 433800
rect 98564 433742 101279 433744
rect 98564 433740 98570 433742
rect 101213 433739 101279 433742
rect 70669 433668 70735 433669
rect 70669 433666 70716 433668
rect 70624 433664 70716 433666
rect 70624 433608 70674 433664
rect 70624 433606 70716 433608
rect 70669 433604 70716 433606
rect 70780 433604 70786 433668
rect 73654 433604 73660 433668
rect 73724 433666 73730 433668
rect 74073 433666 74139 433669
rect 74809 433668 74875 433669
rect 73724 433664 74139 433666
rect 73724 433608 74078 433664
rect 74134 433608 74139 433664
rect 73724 433606 74139 433608
rect 73724 433604 73730 433606
rect 70669 433603 70735 433604
rect 74073 433603 74139 433606
rect 74758 433604 74764 433668
rect 74828 433666 74875 433668
rect 74828 433664 74920 433666
rect 74870 433608 74920 433664
rect 74828 433606 74920 433608
rect 74828 433604 74875 433606
rect 76046 433604 76052 433668
rect 76116 433666 76122 433668
rect 76189 433666 76255 433669
rect 76116 433664 76255 433666
rect 76116 433608 76194 433664
rect 76250 433608 76255 433664
rect 76116 433606 76255 433608
rect 76116 433604 76122 433606
rect 74809 433603 74875 433604
rect 76189 433603 76255 433606
rect 78121 433666 78187 433669
rect 78438 433666 78444 433668
rect 78121 433664 78444 433666
rect 78121 433608 78126 433664
rect 78182 433608 78444 433664
rect 78121 433606 78444 433608
rect 78121 433603 78187 433606
rect 78438 433604 78444 433606
rect 78508 433604 78514 433668
rect 85849 433666 85915 433669
rect 86718 433666 86724 433668
rect 85849 433664 86724 433666
rect 85849 433608 85854 433664
rect 85910 433608 86724 433664
rect 85849 433606 86724 433608
rect 85849 433603 85915 433606
rect 86718 433604 86724 433606
rect 86788 433604 86794 433668
rect 87086 433604 87092 433668
rect 87156 433666 87162 433668
rect 87321 433666 87387 433669
rect 87156 433664 87387 433666
rect 87156 433608 87326 433664
rect 87382 433608 87387 433664
rect 87156 433606 87387 433608
rect 87156 433604 87162 433606
rect 87321 433603 87387 433606
rect 87454 433604 87460 433668
rect 87524 433666 87530 433668
rect 87965 433666 88031 433669
rect 87524 433664 88031 433666
rect 87524 433608 87970 433664
rect 88026 433608 88031 433664
rect 87524 433606 88031 433608
rect 87524 433604 87530 433606
rect 87965 433603 88031 433606
rect 89621 433668 89687 433669
rect 90081 433668 90147 433669
rect 91553 433668 91619 433669
rect 89621 433664 89668 433668
rect 89732 433666 89738 433668
rect 90030 433666 90036 433668
rect 89621 433608 89626 433664
rect 89621 433604 89668 433608
rect 89732 433606 89778 433666
rect 89990 433606 90036 433666
rect 90100 433664 90147 433668
rect 91502 433666 91508 433668
rect 90142 433608 90147 433664
rect 89732 433604 89738 433606
rect 90030 433604 90036 433606
rect 90100 433604 90147 433608
rect 91462 433606 91508 433666
rect 91572 433664 91619 433668
rect 91614 433608 91619 433664
rect 91502 433604 91508 433606
rect 91572 433604 91619 433608
rect 92790 433604 92796 433668
rect 92860 433666 92866 433668
rect 92933 433666 92999 433669
rect 92860 433664 92999 433666
rect 92860 433608 92938 433664
rect 92994 433608 92999 433664
rect 92860 433606 92999 433608
rect 92860 433604 92866 433606
rect 89621 433603 89687 433604
rect 90081 433603 90147 433604
rect 91553 433603 91619 433604
rect 92933 433603 92999 433606
rect 97942 433604 97948 433668
rect 98012 433666 98018 433668
rect 98453 433666 98519 433669
rect 98012 433664 98519 433666
rect 98012 433608 98458 433664
rect 98514 433608 98519 433664
rect 98012 433606 98519 433608
rect 98012 433604 98018 433606
rect 98453 433603 98519 433606
rect 99833 433666 99899 433669
rect 100937 433668 101003 433669
rect 105169 433668 105235 433669
rect 99966 433666 99972 433668
rect 99833 433664 99972 433666
rect 99833 433608 99838 433664
rect 99894 433608 99972 433664
rect 99833 433606 99972 433608
rect 99833 433603 99899 433606
rect 99966 433604 99972 433606
rect 100036 433604 100042 433668
rect 100886 433666 100892 433668
rect 100846 433606 100892 433666
rect 100956 433664 101003 433668
rect 105118 433666 105124 433668
rect 100998 433608 101003 433664
rect 100886 433604 100892 433606
rect 100956 433604 101003 433608
rect 105078 433606 105124 433666
rect 105188 433664 105235 433668
rect 105230 433608 105235 433664
rect 105118 433604 105124 433606
rect 105188 433604 105235 433608
rect 106406 433604 106412 433668
rect 106476 433666 106482 433668
rect 106733 433666 106799 433669
rect 106476 433664 106799 433666
rect 106476 433608 106738 433664
rect 106794 433608 106799 433664
rect 106476 433606 106799 433608
rect 106476 433604 106482 433606
rect 100937 433603 101003 433604
rect 105169 433603 105235 433604
rect 106733 433603 106799 433606
rect 109493 433668 109559 433669
rect 109493 433664 109540 433668
rect 109604 433666 109610 433668
rect 109493 433608 109498 433664
rect 109493 433604 109540 433608
rect 109604 433606 109650 433666
rect 109604 433604 109610 433606
rect 111006 433604 111012 433668
rect 111076 433666 111082 433668
rect 111701 433666 111767 433669
rect 111076 433664 111767 433666
rect 111076 433608 111706 433664
rect 111762 433608 111767 433664
rect 111076 433606 111767 433608
rect 111076 433604 111082 433606
rect 109493 433603 109559 433604
rect 111701 433603 111767 433606
rect 191649 433666 191715 433669
rect 255497 433666 255563 433669
rect 191649 433664 193660 433666
rect 191649 433608 191654 433664
rect 191710 433608 193660 433664
rect 191649 433606 193660 433608
rect 253460 433664 255563 433666
rect 253460 433608 255502 433664
rect 255558 433608 255563 433664
rect 253460 433606 255563 433608
rect 191649 433603 191715 433606
rect 255497 433603 255563 433606
rect 66805 433394 66871 433397
rect 115749 433394 115815 433397
rect 66805 433392 68908 433394
rect 66805 433336 66810 433392
rect 66866 433336 68908 433392
rect 66805 433334 68908 433336
rect 112700 433392 115815 433394
rect 112700 433336 115754 433392
rect 115810 433336 115815 433392
rect 112700 433334 115815 433336
rect 66805 433331 66871 433334
rect 115749 433331 115815 433334
rect 66161 432578 66227 432581
rect 66161 432576 68908 432578
rect 66161 432520 66166 432576
rect 66222 432520 68908 432576
rect 66161 432518 68908 432520
rect 66161 432515 66227 432518
rect 115841 432306 115907 432309
rect 112700 432304 115907 432306
rect 112700 432248 115846 432304
rect 115902 432248 115907 432304
rect 112700 432246 115907 432248
rect 115841 432243 115907 432246
rect 191649 432306 191715 432309
rect 191649 432304 193660 432306
rect 191649 432248 191654 432304
rect 191710 432248 193660 432304
rect 191649 432246 193660 432248
rect 191649 432243 191715 432246
rect 254209 432034 254275 432037
rect 253460 432032 254275 432034
rect 253460 431976 254214 432032
rect 254270 431976 254275 432032
rect 253460 431974 254275 431976
rect 254209 431971 254275 431974
rect 582741 431626 582807 431629
rect 583520 431626 584960 431716
rect 582741 431624 584960 431626
rect 582741 431568 582746 431624
rect 582802 431568 584960 431624
rect 582741 431566 584960 431568
rect 582741 431563 582807 431566
rect 67357 431490 67423 431493
rect 67357 431488 68908 431490
rect 67357 431432 67362 431488
rect 67418 431432 68908 431488
rect 583520 431476 584960 431566
rect 67357 431430 68908 431432
rect 67357 431427 67423 431430
rect 112670 430674 112730 431188
rect 191741 430946 191807 430949
rect 191741 430944 193660 430946
rect 191741 430888 191746 430944
rect 191802 430888 193660 430944
rect 191741 430886 193660 430888
rect 191741 430883 191807 430886
rect 180190 430674 180196 430676
rect 112670 430614 180196 430674
rect 180190 430612 180196 430614
rect 180260 430612 180266 430676
rect 255405 430674 255471 430677
rect 253460 430672 255471 430674
rect 253460 430616 255410 430672
rect 255466 430616 255471 430672
rect 253460 430614 255471 430616
rect 255405 430611 255471 430614
rect 66805 430402 66871 430405
rect 66805 430400 68908 430402
rect 66805 430344 66810 430400
rect 66866 430344 68908 430400
rect 66805 430342 68908 430344
rect 66805 430339 66871 430342
rect 114502 430130 114508 430132
rect 112700 430070 114508 430130
rect 114502 430068 114508 430070
rect 114572 430068 114578 430132
rect 191005 429586 191071 429589
rect 191005 429584 193660 429586
rect 191005 429528 191010 429584
rect 191066 429528 193660 429584
rect 191005 429526 193660 429528
rect 191005 429523 191071 429526
rect 67357 429450 67423 429453
rect 68134 429450 68140 429452
rect 67357 429448 68140 429450
rect 67357 429392 67362 429448
rect 67418 429392 68140 429448
rect 67357 429390 68140 429392
rect 67357 429387 67423 429390
rect 68134 429388 68140 429390
rect 68204 429388 68210 429452
rect 67265 429314 67331 429317
rect 114921 429314 114987 429317
rect 255405 429314 255471 429317
rect 67265 429312 68908 429314
rect 67265 429256 67270 429312
rect 67326 429256 68908 429312
rect 67265 429254 68908 429256
rect 112700 429312 114987 429314
rect 112700 429256 114926 429312
rect 114982 429256 114987 429312
rect 112700 429254 114987 429256
rect 253460 429312 255471 429314
rect 253460 429256 255410 429312
rect 255466 429256 255471 429312
rect 253460 429254 255471 429256
rect 67265 429251 67331 429254
rect 114921 429251 114987 429254
rect 255405 429251 255471 429254
rect 161054 428436 161060 428500
rect 161124 428498 161130 428500
rect 166533 428498 166599 428501
rect 161124 428496 166599 428498
rect 161124 428440 166538 428496
rect 166594 428440 166599 428496
rect 161124 428438 166599 428440
rect 161124 428436 161130 428438
rect 166533 428435 166599 428438
rect 67541 428226 67607 428229
rect 113265 428226 113331 428229
rect 115841 428226 115907 428229
rect 67541 428224 68908 428226
rect 67541 428168 67546 428224
rect 67602 428168 68908 428224
rect 67541 428166 68908 428168
rect 112700 428224 115907 428226
rect 112700 428168 113270 428224
rect 113326 428168 115846 428224
rect 115902 428168 115907 428224
rect 112700 428166 115907 428168
rect 67541 428163 67607 428166
rect 113265 428163 113331 428166
rect 115841 428163 115907 428166
rect 190821 428226 190887 428229
rect 190821 428224 193660 428226
rect 190821 428168 190826 428224
rect 190882 428168 193660 428224
rect 190821 428166 193660 428168
rect 190821 428163 190887 428166
rect 254209 427954 254275 427957
rect 253460 427952 254275 427954
rect 253460 427896 254214 427952
rect 254270 427896 254275 427952
rect 253460 427894 254275 427896
rect 254209 427891 254275 427894
rect 69422 427620 69428 427684
rect 69492 427620 69498 427684
rect 67541 427410 67607 427413
rect 69430 427410 69490 427620
rect 67541 427408 69490 427410
rect 67541 427352 67546 427408
rect 67602 427380 69490 427408
rect 67602 427352 69460 427380
rect 67541 427350 69460 427352
rect 67541 427347 67607 427350
rect 115841 427138 115907 427141
rect 112700 427136 115907 427138
rect 112700 427080 115846 427136
rect 115902 427080 115907 427136
rect 112700 427078 115907 427080
rect 115841 427075 115907 427078
rect 191741 426866 191807 426869
rect 191741 426864 193660 426866
rect 191741 426808 191746 426864
rect 191802 426808 193660 426864
rect 191741 426806 193660 426808
rect 191741 426803 191807 426806
rect 255405 426594 255471 426597
rect 253460 426592 255471 426594
rect 253460 426536 255410 426592
rect 255466 426536 255471 426592
rect 253460 426534 255471 426536
rect 255405 426531 255471 426534
rect 67357 426322 67423 426325
rect 67357 426320 68908 426322
rect 67357 426264 67362 426320
rect 67418 426264 68908 426320
rect 67357 426262 68908 426264
rect 67357 426259 67423 426262
rect 115749 426050 115815 426053
rect 112700 426048 115815 426050
rect 112700 425992 115754 426048
rect 115810 425992 115815 426048
rect 112700 425990 115815 425992
rect 115749 425987 115815 425990
rect 57605 425642 57671 425645
rect 67357 425642 67423 425645
rect 57605 425640 67423 425642
rect 57605 425584 57610 425640
rect 57666 425584 67362 425640
rect 67418 425584 67423 425640
rect 57605 425582 67423 425584
rect 57605 425579 57671 425582
rect 67357 425579 67423 425582
rect 191741 425506 191807 425509
rect 191741 425504 193660 425506
rect 191741 425448 191746 425504
rect 191802 425448 193660 425504
rect 191741 425446 193660 425448
rect 191741 425443 191807 425446
rect 66989 425234 67055 425237
rect 67398 425234 67404 425236
rect 66989 425232 67404 425234
rect 66989 425176 66994 425232
rect 67050 425176 67404 425232
rect 66989 425174 67404 425176
rect 66989 425171 67055 425174
rect 67398 425172 67404 425174
rect 67468 425234 67474 425236
rect 256601 425234 256667 425237
rect 67468 425174 68908 425234
rect 253460 425232 256667 425234
rect 253460 425176 256606 425232
rect 256662 425176 256667 425232
rect 253460 425174 256667 425176
rect 67468 425172 67474 425174
rect 256601 425171 256667 425174
rect 115105 424962 115171 424965
rect 112700 424960 115171 424962
rect 112700 424904 115110 424960
rect 115166 424904 115171 424960
rect 112700 424902 115171 424904
rect 115105 424899 115171 424902
rect 66713 424146 66779 424149
rect 115841 424146 115907 424149
rect 66713 424144 68908 424146
rect 66713 424088 66718 424144
rect 66774 424088 68908 424144
rect 66713 424086 68908 424088
rect 112700 424144 115907 424146
rect 112700 424088 115846 424144
rect 115902 424088 115907 424144
rect 112700 424086 115907 424088
rect 66713 424083 66779 424086
rect 115841 424083 115907 424086
rect 191005 423874 191071 423877
rect 191005 423872 193660 423874
rect 191005 423816 191010 423872
rect 191066 423816 193660 423872
rect 191005 423814 193660 423816
rect 191005 423811 191071 423814
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect 255497 423602 255563 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect 253460 423600 255563 423602
rect 253460 423544 255502 423600
rect 255558 423544 255563 423600
rect 253460 423542 255563 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 255497 423539 255563 423542
rect 66805 423330 66871 423333
rect 66805 423328 68908 423330
rect 66805 423272 66810 423328
rect 66866 423272 68908 423328
rect 66805 423270 68908 423272
rect 66805 423267 66871 423270
rect 114553 423058 114619 423061
rect 115841 423058 115907 423061
rect 112700 423056 115907 423058
rect 112700 423000 114558 423056
rect 114614 423000 115846 423056
rect 115902 423000 115907 423056
rect 112700 422998 115907 423000
rect 114553 422995 114619 422998
rect 115841 422995 115907 422998
rect 191741 422514 191807 422517
rect 191741 422512 193660 422514
rect 191741 422456 191746 422512
rect 191802 422456 193660 422512
rect 191741 422454 193660 422456
rect 191741 422451 191807 422454
rect 67541 422242 67607 422245
rect 255497 422242 255563 422245
rect 67541 422240 68908 422242
rect 67541 422184 67546 422240
rect 67602 422184 68908 422240
rect 67541 422182 68908 422184
rect 253460 422240 255563 422242
rect 253460 422184 255502 422240
rect 255558 422184 255563 422240
rect 253460 422182 255563 422184
rect 67541 422179 67607 422182
rect 255497 422179 255563 422182
rect 115289 421970 115355 421973
rect 112700 421968 115355 421970
rect 112700 421912 115294 421968
rect 115350 421912 115355 421968
rect 112700 421910 115355 421912
rect 115289 421907 115355 421910
rect 66805 421154 66871 421157
rect 66805 421152 68908 421154
rect 66805 421096 66810 421152
rect 66866 421096 68908 421152
rect 66805 421094 68908 421096
rect 66805 421091 66871 421094
rect 193630 421018 193690 421124
rect 190410 420958 193690 421018
rect 113173 420882 113239 420885
rect 112700 420880 113239 420882
rect 112700 420824 113178 420880
rect 113234 420824 113239 420880
rect 112700 420822 113239 420824
rect 113173 420819 113239 420822
rect 153101 420882 153167 420885
rect 190410 420882 190470 420958
rect 255497 420882 255563 420885
rect 153101 420880 190470 420882
rect 153101 420824 153106 420880
rect 153162 420824 190470 420880
rect 153101 420822 190470 420824
rect 253460 420880 255563 420882
rect 253460 420824 255502 420880
rect 255558 420824 255563 420880
rect 253460 420822 255563 420824
rect 153101 420819 153167 420822
rect 255497 420819 255563 420822
rect 66897 420066 66963 420069
rect 114645 420066 114711 420069
rect 66897 420064 68908 420066
rect 66897 420008 66902 420064
rect 66958 420008 68908 420064
rect 66897 420006 68908 420008
rect 112700 420064 114711 420066
rect 112700 420008 114650 420064
rect 114706 420008 114711 420064
rect 112700 420006 114711 420008
rect 66897 420003 66963 420006
rect 114645 420003 114711 420006
rect 192385 419794 192451 419797
rect 193121 419794 193187 419797
rect 192385 419792 193660 419794
rect 192385 419736 192390 419792
rect 192446 419736 193126 419792
rect 193182 419736 193660 419792
rect 192385 419734 193660 419736
rect 192385 419731 192451 419734
rect 193121 419731 193187 419734
rect 255405 419522 255471 419525
rect 253460 419520 255471 419522
rect 253460 419464 255410 419520
rect 255466 419464 255471 419520
rect 253460 419462 255471 419464
rect 255405 419459 255471 419462
rect 66437 418978 66503 418981
rect 113357 418978 113423 418981
rect 115841 418978 115907 418981
rect 66437 418976 68908 418978
rect 66437 418920 66442 418976
rect 66498 418920 68908 418976
rect 66437 418918 68908 418920
rect 112700 418976 115907 418978
rect 112700 418920 113362 418976
rect 113418 418920 115846 418976
rect 115902 418920 115907 418976
rect 112700 418918 115907 418920
rect 66437 418915 66503 418918
rect 113357 418915 113423 418918
rect 115841 418915 115907 418918
rect 159766 418780 159772 418844
rect 159836 418842 159842 418844
rect 166390 418842 166396 418844
rect 159836 418782 166396 418842
rect 159836 418780 159842 418782
rect 166390 418780 166396 418782
rect 166460 418780 166466 418844
rect 150934 418236 150940 418300
rect 151004 418298 151010 418300
rect 193630 418298 193690 418404
rect 151004 418238 193690 418298
rect 582373 418298 582439 418301
rect 583520 418298 584960 418388
rect 582373 418296 584960 418298
rect 582373 418240 582378 418296
rect 582434 418240 584960 418296
rect 582373 418238 584960 418240
rect 151004 418236 151010 418238
rect 582373 418235 582439 418238
rect 66437 418162 66503 418165
rect 67541 418162 67607 418165
rect 255497 418162 255563 418165
rect 66437 418160 68908 418162
rect 66437 418104 66442 418160
rect 66498 418104 67546 418160
rect 67602 418104 68908 418160
rect 66437 418102 68908 418104
rect 253460 418160 255563 418162
rect 253460 418104 255502 418160
rect 255558 418104 255563 418160
rect 583520 418148 584960 418238
rect 253460 418102 255563 418104
rect 66437 418099 66503 418102
rect 67541 418099 67607 418102
rect 255497 418099 255563 418102
rect 114553 417890 114619 417893
rect 112700 417888 114619 417890
rect 112700 417832 114558 417888
rect 114614 417832 114619 417888
rect 112700 417830 114619 417832
rect 114553 417827 114619 417830
rect 180517 417484 180583 417485
rect 180517 417482 180564 417484
rect 180472 417480 180564 417482
rect 180472 417424 180522 417480
rect 180472 417422 180564 417424
rect 180517 417420 180564 417422
rect 180628 417420 180634 417484
rect 180517 417419 180583 417420
rect 66805 417074 66871 417077
rect 191741 417074 191807 417077
rect 66805 417072 68908 417074
rect 66805 417016 66810 417072
rect 66866 417016 68908 417072
rect 66805 417014 68908 417016
rect 191741 417072 193660 417074
rect 191741 417016 191746 417072
rect 191802 417016 193660 417072
rect 191741 417014 193660 417016
rect 66805 417011 66871 417014
rect 191741 417011 191807 417014
rect 115841 416802 115907 416805
rect 255405 416802 255471 416805
rect 112700 416800 115907 416802
rect 112700 416744 115846 416800
rect 115902 416744 115907 416800
rect 112700 416742 115907 416744
rect 253460 416800 255471 416802
rect 253460 416744 255410 416800
rect 255466 416744 255471 416800
rect 253460 416742 255471 416744
rect 115841 416739 115907 416742
rect 255405 416739 255471 416742
rect 279325 416666 279391 416669
rect 281574 416666 281580 416668
rect 279325 416664 281580 416666
rect 279325 416608 279330 416664
rect 279386 416608 281580 416664
rect 279325 416606 281580 416608
rect 279325 416603 279391 416606
rect 281574 416604 281580 416606
rect 281644 416604 281650 416668
rect 66897 415986 66963 415989
rect 66897 415984 68908 415986
rect 66897 415928 66902 415984
rect 66958 415928 68908 415984
rect 66897 415926 68908 415928
rect 66897 415923 66963 415926
rect 115841 415714 115907 415717
rect 112700 415712 115907 415714
rect 112700 415656 115846 415712
rect 115902 415656 115907 415712
rect 112700 415654 115907 415656
rect 115841 415651 115907 415654
rect 191649 415442 191715 415445
rect 191649 415440 193660 415442
rect 191649 415384 191654 415440
rect 191710 415384 193660 415440
rect 191649 415382 193660 415384
rect 191649 415379 191715 415382
rect 254117 415170 254183 415173
rect 255313 415170 255379 415173
rect 253460 415168 255379 415170
rect 253460 415112 254122 415168
rect 254178 415112 255318 415168
rect 255374 415112 255379 415168
rect 253460 415110 255379 415112
rect 254117 415107 254183 415110
rect 255313 415107 255379 415110
rect 66805 414898 66871 414901
rect 114921 414898 114987 414901
rect 66805 414896 68908 414898
rect 66805 414840 66810 414896
rect 66866 414840 68908 414896
rect 66805 414838 68908 414840
rect 112700 414896 114987 414898
rect 112700 414840 114926 414896
rect 114982 414840 114987 414896
rect 112700 414838 114987 414840
rect 66805 414835 66871 414838
rect 114921 414835 114987 414838
rect 159766 414564 159772 414628
rect 159836 414626 159842 414628
rect 166349 414626 166415 414629
rect 159836 414624 166415 414626
rect 159836 414568 166354 414624
rect 166410 414568 166415 414624
rect 159836 414566 166415 414568
rect 159836 414564 159842 414566
rect 166349 414563 166415 414566
rect 67357 414082 67423 414085
rect 191189 414082 191255 414085
rect 67357 414080 68908 414082
rect 67357 414024 67362 414080
rect 67418 414024 68908 414080
rect 67357 414022 68908 414024
rect 191189 414080 193660 414082
rect 191189 414024 191194 414080
rect 191250 414024 193660 414080
rect 191189 414022 193660 414024
rect 67357 414019 67423 414022
rect 191189 414019 191255 414022
rect 114686 413810 114692 413812
rect 112700 413750 114692 413810
rect 114686 413748 114692 413750
rect 114756 413810 114762 413812
rect 115197 413810 115263 413813
rect 114756 413808 115263 413810
rect 114756 413752 115202 413808
rect 115258 413752 115263 413808
rect 114756 413750 115263 413752
rect 114756 413748 114762 413750
rect 115197 413747 115263 413750
rect 253430 413674 253490 413780
rect 253565 413674 253631 413677
rect 253430 413672 253631 413674
rect 253430 413616 253570 413672
rect 253626 413616 253631 413672
rect 253430 413614 253631 413616
rect 253565 413611 253631 413614
rect 179270 413204 179276 413268
rect 179340 413266 179346 413268
rect 192569 413266 192635 413269
rect 179340 413264 192635 413266
rect 179340 413208 192574 413264
rect 192630 413208 192635 413264
rect 179340 413206 192635 413208
rect 179340 413204 179346 413206
rect 192569 413203 192635 413206
rect 66621 412994 66687 412997
rect 66621 412992 68908 412994
rect 66621 412936 66626 412992
rect 66682 412936 68908 412992
rect 66621 412934 68908 412936
rect 66621 412931 66687 412934
rect 115841 412722 115907 412725
rect 112700 412720 115907 412722
rect 112700 412664 115846 412720
rect 115902 412664 115907 412720
rect 112700 412662 115907 412664
rect 115841 412659 115907 412662
rect 191097 412722 191163 412725
rect 191097 412720 193660 412722
rect 191097 412664 191102 412720
rect 191158 412664 193660 412720
rect 191097 412662 193660 412664
rect 191097 412659 191163 412662
rect 255497 412450 255563 412453
rect 253460 412448 255563 412450
rect 253460 412392 255502 412448
rect 255558 412392 255563 412448
rect 253460 412390 255563 412392
rect 255497 412387 255563 412390
rect 66897 411906 66963 411909
rect 66897 411904 68908 411906
rect 66897 411848 66902 411904
rect 66958 411848 68908 411904
rect 66897 411846 68908 411848
rect 66897 411843 66963 411846
rect 115749 411634 115815 411637
rect 112700 411632 115815 411634
rect 112700 411576 115754 411632
rect 115810 411576 115815 411632
rect 112700 411574 115815 411576
rect 115749 411571 115815 411574
rect 191741 411362 191807 411365
rect 191741 411360 193660 411362
rect 191741 411304 191746 411360
rect 191802 411304 193660 411360
rect 191741 411302 193660 411304
rect 191741 411299 191807 411302
rect 255497 411090 255563 411093
rect 253460 411088 255563 411090
rect 253460 411032 255502 411088
rect 255558 411032 255563 411088
rect 253460 411030 255563 411032
rect 255497 411027 255563 411030
rect 66805 410818 66871 410821
rect 66805 410816 68908 410818
rect 66805 410760 66810 410816
rect 66866 410760 68908 410816
rect 66805 410758 68908 410760
rect 66805 410755 66871 410758
rect -960 410546 480 410636
rect 3509 410546 3575 410549
rect 115841 410546 115907 410549
rect -960 410544 3575 410546
rect -960 410488 3514 410544
rect 3570 410488 3575 410544
rect -960 410486 3575 410488
rect 112700 410544 115907 410546
rect 112700 410488 115846 410544
rect 115902 410488 115907 410544
rect 112700 410486 115907 410488
rect -960 410396 480 410486
rect 3509 410483 3575 410486
rect 115841 410483 115907 410486
rect 191741 410002 191807 410005
rect 191741 410000 193660 410002
rect 191741 409944 191746 410000
rect 191802 409944 193660 410000
rect 191741 409942 193660 409944
rect 191741 409939 191807 409942
rect 67633 409730 67699 409733
rect 115841 409730 115907 409733
rect 255405 409730 255471 409733
rect 67633 409728 68908 409730
rect 67633 409672 67638 409728
rect 67694 409672 68908 409728
rect 67633 409670 68908 409672
rect 112700 409728 115907 409730
rect 112700 409672 115846 409728
rect 115902 409672 115907 409728
rect 112700 409670 115907 409672
rect 253460 409728 255471 409730
rect 253460 409672 255410 409728
rect 255466 409672 255471 409728
rect 253460 409670 255471 409672
rect 67633 409667 67699 409670
rect 115841 409667 115907 409670
rect 255405 409667 255471 409670
rect 66437 408914 66503 408917
rect 66437 408912 68908 408914
rect 66437 408856 66442 408912
rect 66498 408856 68908 408912
rect 66437 408854 68908 408856
rect 66437 408851 66503 408854
rect 115841 408642 115907 408645
rect 112700 408640 115907 408642
rect 112700 408584 115846 408640
rect 115902 408584 115907 408640
rect 112700 408582 115907 408584
rect 115841 408579 115907 408582
rect 192477 408642 192543 408645
rect 192477 408640 193660 408642
rect 192477 408584 192482 408640
rect 192538 408584 193660 408640
rect 192477 408582 193660 408584
rect 192477 408579 192543 408582
rect 255405 408370 255471 408373
rect 253460 408368 255471 408370
rect 253460 408312 255410 408368
rect 255466 408312 255471 408368
rect 253460 408310 255471 408312
rect 255405 408307 255471 408310
rect 66805 407826 66871 407829
rect 66805 407824 68908 407826
rect 66805 407768 66810 407824
rect 66866 407768 68908 407824
rect 66805 407766 68908 407768
rect 66805 407763 66871 407766
rect 112670 407146 112730 407524
rect 113081 407146 113147 407149
rect 112670 407144 113147 407146
rect 112670 407088 113086 407144
rect 113142 407088 113147 407144
rect 112670 407086 113147 407088
rect 113081 407083 113147 407086
rect 191005 407010 191071 407013
rect 255497 407010 255563 407013
rect 191005 407008 193660 407010
rect 191005 406952 191010 407008
rect 191066 406952 193660 407008
rect 191005 406950 193660 406952
rect 253460 407008 255563 407010
rect 253460 406952 255502 407008
rect 255558 406952 255563 407008
rect 253460 406950 255563 406952
rect 191005 406947 191071 406950
rect 255497 406947 255563 406950
rect 66437 406738 66503 406741
rect 66437 406736 68908 406738
rect 66437 406680 66442 406736
rect 66498 406680 68908 406736
rect 66437 406678 68908 406680
rect 66437 406675 66503 406678
rect 114461 406466 114527 406469
rect 115197 406466 115263 406469
rect 112700 406464 115263 406466
rect 112700 406408 114466 406464
rect 114522 406408 115202 406464
rect 115258 406408 115263 406464
rect 112700 406406 115263 406408
rect 114461 406403 114527 406406
rect 115197 406403 115263 406406
rect 67449 405650 67515 405653
rect 115841 405650 115907 405653
rect 67449 405648 68908 405650
rect 67449 405592 67454 405648
rect 67510 405592 68908 405648
rect 67449 405590 68908 405592
rect 112700 405648 115907 405650
rect 112700 405592 115846 405648
rect 115902 405592 115907 405648
rect 112700 405590 115907 405592
rect 67449 405587 67515 405590
rect 115841 405587 115907 405590
rect 191741 405650 191807 405653
rect 191741 405648 193660 405650
rect 191741 405592 191746 405648
rect 191802 405592 193660 405648
rect 191741 405590 193660 405592
rect 191741 405587 191807 405590
rect 252878 404836 252938 405348
rect 582465 404970 582531 404973
rect 583520 404970 584960 405060
rect 582465 404968 584960 404970
rect 582465 404912 582470 404968
rect 582526 404912 584960 404968
rect 582465 404910 584960 404912
rect 582465 404907 582531 404910
rect 252870 404772 252876 404836
rect 252940 404772 252946 404836
rect 583520 404820 584960 404910
rect 66897 404562 66963 404565
rect 115841 404562 115907 404565
rect 66897 404560 68908 404562
rect 66897 404504 66902 404560
rect 66958 404504 68908 404560
rect 66897 404502 68908 404504
rect 112700 404560 115907 404562
rect 112700 404504 115846 404560
rect 115902 404504 115907 404560
rect 112700 404502 115907 404504
rect 66897 404499 66963 404502
rect 115841 404499 115907 404502
rect 191741 404290 191807 404293
rect 191741 404288 193660 404290
rect 191741 404232 191746 404288
rect 191802 404232 193660 404288
rect 191741 404230 193660 404232
rect 191741 404227 191807 404230
rect 255405 404018 255471 404021
rect 253460 404016 255471 404018
rect 253460 403960 255410 404016
rect 255466 403960 255471 404016
rect 253460 403958 255471 403960
rect 255405 403955 255471 403958
rect 66437 403746 66503 403749
rect 66437 403744 68908 403746
rect 66437 403688 66442 403744
rect 66498 403688 68908 403744
rect 66437 403686 68908 403688
rect 66437 403683 66503 403686
rect 115841 403474 115907 403477
rect 112700 403472 115907 403474
rect 112700 403416 115846 403472
rect 115902 403416 115907 403472
rect 112700 403414 115907 403416
rect 115841 403411 115907 403414
rect 191005 402930 191071 402933
rect 191005 402928 193660 402930
rect 191005 402872 191010 402928
rect 191066 402872 193660 402928
rect 191005 402870 193660 402872
rect 191005 402867 191071 402870
rect 67633 402658 67699 402661
rect 67633 402656 68908 402658
rect 67633 402600 67638 402656
rect 67694 402600 68908 402656
rect 67633 402598 68908 402600
rect 67633 402595 67699 402598
rect 112110 402596 112116 402660
rect 112180 402596 112186 402660
rect 255405 402658 255471 402661
rect 253460 402656 255471 402658
rect 253460 402600 255410 402656
rect 255466 402600 255471 402656
rect 253460 402598 255471 402600
rect 112118 402386 112178 402596
rect 255405 402595 255471 402598
rect 113449 402386 113515 402389
rect 112118 402384 113515 402386
rect 112118 402356 113454 402384
rect 112148 402328 113454 402356
rect 113510 402328 113515 402384
rect 112148 402326 113515 402328
rect 113449 402323 113515 402326
rect 66437 401570 66503 401573
rect 191741 401570 191807 401573
rect 66437 401568 68908 401570
rect 66437 401512 66442 401568
rect 66498 401512 68908 401568
rect 66437 401510 68908 401512
rect 191741 401568 193660 401570
rect 191741 401512 191746 401568
rect 191802 401512 193660 401568
rect 191741 401510 193660 401512
rect 66437 401507 66503 401510
rect 191741 401507 191807 401510
rect 115381 401298 115447 401301
rect 255405 401298 255471 401301
rect 112700 401296 115447 401298
rect 112700 401240 115386 401296
rect 115442 401240 115447 401296
rect 112700 401238 115447 401240
rect 253460 401296 255471 401298
rect 253460 401240 255410 401296
rect 255466 401240 255471 401296
rect 253460 401238 255471 401240
rect 115381 401235 115447 401238
rect 255405 401235 255471 401238
rect 67265 400482 67331 400485
rect 114829 400482 114895 400485
rect 67265 400480 68908 400482
rect 67265 400424 67270 400480
rect 67326 400424 68908 400480
rect 67265 400422 68908 400424
rect 112700 400480 114895 400482
rect 112700 400424 114834 400480
rect 114890 400424 114895 400480
rect 112700 400422 114895 400424
rect 67265 400419 67331 400422
rect 114829 400419 114895 400422
rect 191005 400210 191071 400213
rect 191005 400208 193660 400210
rect 191005 400152 191010 400208
rect 191066 400152 193660 400208
rect 191005 400150 193660 400152
rect 191005 400147 191071 400150
rect 255405 399938 255471 399941
rect 253460 399936 255471 399938
rect 253460 399880 255410 399936
rect 255466 399880 255471 399936
rect 253460 399878 255471 399880
rect 255405 399875 255471 399878
rect 66805 399666 66871 399669
rect 66805 399664 68908 399666
rect 66805 399608 66810 399664
rect 66866 399608 68908 399664
rect 66805 399606 68908 399608
rect 66805 399603 66871 399606
rect 115841 399394 115907 399397
rect 112700 399392 115907 399394
rect 112700 399336 115846 399392
rect 115902 399336 115907 399392
rect 112700 399334 115907 399336
rect 115841 399331 115907 399334
rect 112110 398924 112116 398988
rect 112180 398986 112186 398988
rect 113030 398986 113036 398988
rect 112180 398926 113036 398986
rect 112180 398924 112186 398926
rect 113030 398924 113036 398926
rect 113100 398986 113106 398988
rect 155217 398986 155283 398989
rect 113100 398984 155283 398986
rect 113100 398928 155222 398984
rect 155278 398928 155283 398984
rect 113100 398926 155283 398928
rect 113100 398924 113106 398926
rect 155217 398923 155283 398926
rect 177798 398788 177804 398852
rect 177868 398850 177874 398852
rect 178033 398850 178099 398853
rect 177868 398848 178099 398850
rect 177868 398792 178038 398848
rect 178094 398792 178099 398848
rect 177868 398790 178099 398792
rect 177868 398788 177874 398790
rect 178033 398787 178099 398790
rect 67081 398578 67147 398581
rect 67449 398578 67515 398581
rect 190821 398578 190887 398581
rect 258993 398578 259059 398581
rect 67081 398576 68908 398578
rect 67081 398520 67086 398576
rect 67142 398520 67454 398576
rect 67510 398520 68908 398576
rect 67081 398518 68908 398520
rect 190821 398576 193660 398578
rect 190821 398520 190826 398576
rect 190882 398520 193660 398576
rect 190821 398518 193660 398520
rect 253460 398576 259059 398578
rect 253460 398520 258998 398576
rect 259054 398520 259059 398576
rect 253460 398518 259059 398520
rect 67081 398515 67147 398518
rect 67449 398515 67515 398518
rect 190821 398515 190887 398518
rect 258993 398515 259059 398518
rect 115841 398306 115907 398309
rect 112700 398304 115907 398306
rect 112700 398248 115846 398304
rect 115902 398248 115907 398304
rect 112700 398246 115907 398248
rect 115841 398243 115907 398246
rect 149053 398034 149119 398037
rect 150341 398034 150407 398037
rect 173157 398034 173223 398037
rect 149053 398032 173223 398034
rect 149053 397976 149058 398032
rect 149114 397976 150346 398032
rect 150402 397976 173162 398032
rect 173218 397976 173223 398032
rect 149053 397974 173223 397976
rect 149053 397971 149119 397974
rect 150341 397971 150407 397974
rect 173157 397971 173223 397974
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 66662 397428 66668 397492
rect 66732 397490 66738 397492
rect 66805 397490 66871 397493
rect 66732 397488 68908 397490
rect 66732 397432 66810 397488
rect 66866 397432 68908 397488
rect 66732 397430 68908 397432
rect 66732 397428 66738 397430
rect 66805 397427 66871 397430
rect 253054 397292 253060 397356
rect 253124 397292 253130 397356
rect 115841 397218 115907 397221
rect 112700 397216 115907 397218
rect 112700 397160 115846 397216
rect 115902 397160 115907 397216
rect 112700 397158 115907 397160
rect 115841 397155 115907 397158
rect 191189 397218 191255 397221
rect 191189 397216 193660 397218
rect 191189 397160 191194 397216
rect 191250 397160 193660 397216
rect 191189 397158 193660 397160
rect 191189 397155 191255 397158
rect 253062 396946 253122 397292
rect 253974 396946 253980 396948
rect 253062 396916 253980 396946
rect 253092 396886 253980 396916
rect 253974 396884 253980 396886
rect 254044 396884 254050 396948
rect 66253 396402 66319 396405
rect 113214 396402 113220 396404
rect 66253 396400 68908 396402
rect 66253 396344 66258 396400
rect 66314 396344 68908 396400
rect 66253 396342 68908 396344
rect 112700 396342 113220 396402
rect 66253 396339 66319 396342
rect 113214 396340 113220 396342
rect 113284 396402 113290 396404
rect 115749 396402 115815 396405
rect 113284 396400 115815 396402
rect 113284 396344 115754 396400
rect 115810 396344 115815 396400
rect 113284 396342 115815 396344
rect 113284 396340 113290 396342
rect 115749 396339 115815 396342
rect 191741 395858 191807 395861
rect 191741 395856 193660 395858
rect 191741 395800 191746 395856
rect 191802 395800 193660 395856
rect 191741 395798 193660 395800
rect 191741 395795 191807 395798
rect 255405 395586 255471 395589
rect 253460 395584 255471 395586
rect 253460 395528 255410 395584
rect 255466 395528 255471 395584
rect 253460 395526 255471 395528
rect 255405 395523 255471 395526
rect 66662 395252 66668 395316
rect 66732 395314 66738 395316
rect 115841 395314 115907 395317
rect 66732 395254 68908 395314
rect 112700 395312 115907 395314
rect 112700 395256 115846 395312
rect 115902 395256 115907 395312
rect 112700 395254 115907 395256
rect 66732 395252 66738 395254
rect 115841 395251 115907 395254
rect 254526 394572 254532 394636
rect 254596 394634 254602 394636
rect 256877 394634 256943 394637
rect 254596 394632 256943 394634
rect 254596 394576 256882 394632
rect 256938 394576 256943 394632
rect 254596 394574 256943 394576
rect 254596 394572 254602 394574
rect 256877 394571 256943 394574
rect 69430 393956 69490 394468
rect 115841 394226 115907 394229
rect 112700 394224 115907 394226
rect 112700 394168 115846 394224
rect 115902 394168 115907 394224
rect 112700 394166 115907 394168
rect 115841 394163 115907 394166
rect 180701 394090 180767 394093
rect 188521 394090 188587 394093
rect 180701 394088 188587 394090
rect 180701 394032 180706 394088
rect 180762 394032 188526 394088
rect 188582 394032 188587 394088
rect 180701 394030 188587 394032
rect 180701 394027 180767 394030
rect 188521 394027 188587 394030
rect 69422 393892 69428 393956
rect 69492 393892 69498 393956
rect 172421 393954 172487 393957
rect 172421 393952 180810 393954
rect 172421 393896 172426 393952
rect 172482 393896 180810 393952
rect 172421 393894 180810 393896
rect 172421 393891 172487 393894
rect 180750 393413 180810 393894
rect 67725 393410 67791 393413
rect 180750 393410 180859 393413
rect 193630 393410 193690 394468
rect 255405 394226 255471 394229
rect 253460 394224 255471 394226
rect 253460 394168 255410 394224
rect 255466 394168 255471 394224
rect 253460 394166 255471 394168
rect 255405 394163 255471 394166
rect 67725 393408 68908 393410
rect 67725 393352 67730 393408
rect 67786 393352 68908 393408
rect 67725 393350 68908 393352
rect 180750 393408 193690 393410
rect 180750 393352 180798 393408
rect 180854 393352 193690 393408
rect 180750 393350 193690 393352
rect 67725 393347 67791 393350
rect 180793 393347 180859 393350
rect 115841 393138 115907 393141
rect 112700 393136 115907 393138
rect 112700 393080 115846 393136
rect 115902 393080 115907 393136
rect 112700 393078 115907 393080
rect 115841 393075 115907 393078
rect 66621 392322 66687 392325
rect 66621 392320 68908 392322
rect 66621 392264 66626 392320
rect 66682 392264 68908 392320
rect 66621 392262 68908 392264
rect 66621 392259 66687 392262
rect 115841 392050 115907 392053
rect 112700 392048 115907 392050
rect 112700 391992 115846 392048
rect 115902 391992 115907 392048
rect 112700 391990 115907 391992
rect 115841 391987 115907 391990
rect 179413 392050 179479 392053
rect 180701 392050 180767 392053
rect 193630 392050 193690 393108
rect 254025 392866 254091 392869
rect 253460 392864 254091 392866
rect 253460 392808 254030 392864
rect 254086 392808 254091 392864
rect 253460 392806 254091 392808
rect 254025 392803 254091 392806
rect 254710 392532 254716 392596
rect 254780 392594 254786 392596
rect 268009 392594 268075 392597
rect 254780 392592 268075 392594
rect 254780 392536 268014 392592
rect 268070 392536 268075 392592
rect 254780 392534 268075 392536
rect 254780 392532 254786 392534
rect 268009 392531 268075 392534
rect 254025 392052 254091 392053
rect 179413 392048 193690 392050
rect 179413 391992 179418 392048
rect 179474 391992 180706 392048
rect 180762 391992 193690 392048
rect 179413 391990 193690 391992
rect 179413 391987 179479 391990
rect 180701 391987 180767 391990
rect 253974 391988 253980 392052
rect 254044 392050 254091 392052
rect 254044 392048 254136 392050
rect 254086 391992 254136 392048
rect 254044 391990 254136 391992
rect 254044 391988 254091 391990
rect 254025 391987 254091 391988
rect 7557 391914 7623 391917
rect 82302 391914 82308 391916
rect 7557 391912 82308 391914
rect 7557 391856 7562 391912
rect 7618 391856 82308 391912
rect 7557 391854 82308 391856
rect 7557 391851 7623 391854
rect 82302 391852 82308 391854
rect 82372 391914 82378 391916
rect 82670 391914 82676 391916
rect 82372 391854 82676 391914
rect 82372 391852 82378 391854
rect 82670 391852 82676 391854
rect 82740 391914 82746 391916
rect 128997 391914 129063 391917
rect 82740 391912 129063 391914
rect 82740 391856 129002 391912
rect 129058 391856 129063 391912
rect 82740 391854 129063 391856
rect 82740 391852 82746 391854
rect 128997 391851 129063 391854
rect 59077 391506 59143 391509
rect 114686 391506 114692 391508
rect 59077 391504 89730 391506
rect 59077 391448 59082 391504
rect 59138 391448 89730 391504
rect 59077 391446 89730 391448
rect 59077 391443 59143 391446
rect 68553 391234 68619 391237
rect 68553 391232 68908 391234
rect 68553 391176 68558 391232
rect 68614 391176 68908 391232
rect 68553 391174 68908 391176
rect 68553 391171 68619 391174
rect 82169 390962 82235 390965
rect 82302 390962 82308 390964
rect 82169 390960 82308 390962
rect 82169 390904 82174 390960
rect 82230 390904 82308 390960
rect 82169 390902 82308 390904
rect 82169 390899 82235 390902
rect 82302 390900 82308 390902
rect 82372 390900 82378 390964
rect 84510 390900 84516 390964
rect 84580 390962 84586 390964
rect 85481 390962 85547 390965
rect 84580 390960 85547 390962
rect 84580 390904 85486 390960
rect 85542 390904 85547 390960
rect 84580 390902 85547 390904
rect 89670 390962 89730 391446
rect 106046 391446 114692 391506
rect 106046 390965 106106 391446
rect 114686 391444 114692 391446
rect 114756 391444 114762 391508
rect 161197 391234 161263 391237
rect 161197 391232 171150 391234
rect 99465 390962 99531 390965
rect 89670 390960 99531 390962
rect 89670 390904 99470 390960
rect 99526 390904 99531 390960
rect 89670 390902 99531 390904
rect 84580 390900 84586 390902
rect 85481 390899 85547 390902
rect 99465 390899 99531 390902
rect 105997 390960 106106 390965
rect 105997 390904 106002 390960
rect 106058 390904 106106 390960
rect 105997 390902 106106 390904
rect 107377 390962 107443 390965
rect 107510 390962 107516 390964
rect 107377 390960 107516 390962
rect 107377 390904 107382 390960
rect 107438 390904 107516 390960
rect 107377 390902 107516 390904
rect 105997 390899 106063 390902
rect 107377 390899 107443 390902
rect 107510 390900 107516 390902
rect 107580 390900 107586 390964
rect 91318 390764 91324 390828
rect 91388 390826 91394 390828
rect 92013 390826 92079 390829
rect 96797 390828 96863 390829
rect 97073 390828 97139 390829
rect 96797 390826 96844 390828
rect 91388 390824 92079 390826
rect 91388 390768 92018 390824
rect 92074 390768 92079 390824
rect 91388 390766 92079 390768
rect 96752 390824 96844 390826
rect 96752 390768 96802 390824
rect 96752 390766 96844 390768
rect 91388 390764 91394 390766
rect 92013 390763 92079 390766
rect 96797 390764 96844 390766
rect 96908 390764 96914 390828
rect 97022 390764 97028 390828
rect 97092 390826 97139 390828
rect 97092 390824 97184 390826
rect 97134 390768 97184 390824
rect 97092 390766 97184 390768
rect 97092 390764 97139 390766
rect 96797 390763 96863 390764
rect 97073 390763 97139 390764
rect 82854 390628 82860 390692
rect 82924 390690 82930 390692
rect 83181 390690 83247 390693
rect 82924 390688 83247 390690
rect 82924 390632 83186 390688
rect 83242 390632 83247 390688
rect 82924 390630 83247 390632
rect 82924 390628 82930 390630
rect 83181 390627 83247 390630
rect 88926 390628 88932 390692
rect 88996 390690 89002 390692
rect 89713 390690 89779 390693
rect 88996 390688 89779 390690
rect 88996 390632 89718 390688
rect 89774 390632 89779 390688
rect 88996 390630 89779 390632
rect 112670 390690 112730 391204
rect 161197 391176 161202 391232
rect 161258 391176 171150 391232
rect 161197 391174 171150 391176
rect 161197 391171 161263 391174
rect 170949 390826 171015 390829
rect 171090 390826 171150 391174
rect 192661 391098 192727 391101
rect 193397 391098 193463 391101
rect 192661 391096 193463 391098
rect 192661 391040 192666 391096
rect 192722 391040 193402 391096
rect 193458 391040 193463 391096
rect 192661 391038 193463 391040
rect 192661 391035 192727 391038
rect 193397 391035 193463 391038
rect 177297 390962 177363 390965
rect 178033 390962 178099 390965
rect 177297 390960 178099 390962
rect 177297 390904 177302 390960
rect 177358 390904 178038 390960
rect 178094 390904 178099 390960
rect 177297 390902 178099 390904
rect 177297 390899 177363 390902
rect 178033 390899 178099 390902
rect 186313 390962 186379 390965
rect 193121 390962 193187 390965
rect 186313 390960 193187 390962
rect 186313 390904 186318 390960
rect 186374 390904 193126 390960
rect 193182 390904 193187 390960
rect 186313 390902 193187 390904
rect 186313 390899 186379 390902
rect 193121 390899 193187 390902
rect 193630 390826 193690 391748
rect 583520 391628 584960 391868
rect 248873 390962 248939 390965
rect 249006 390962 249012 390964
rect 248873 390960 249012 390962
rect 248873 390904 248878 390960
rect 248934 390904 249012 390960
rect 248873 390902 249012 390904
rect 248873 390899 248939 390902
rect 249006 390900 249012 390902
rect 249076 390900 249082 390964
rect 252553 390962 252619 390965
rect 252878 390962 252938 391476
rect 252553 390960 252938 390962
rect 252553 390904 252558 390960
rect 252614 390904 252938 390960
rect 252553 390902 252938 390904
rect 252553 390899 252619 390902
rect 170949 390824 193690 390826
rect 170949 390768 170954 390824
rect 171010 390768 193690 390824
rect 170949 390766 193690 390768
rect 250713 390826 250779 390829
rect 258165 390826 258231 390829
rect 250713 390824 258231 390826
rect 250713 390768 250718 390824
rect 250774 390768 258170 390824
rect 258226 390768 258231 390824
rect 250713 390766 258231 390768
rect 170949 390763 171015 390766
rect 250713 390763 250779 390766
rect 258165 390763 258231 390766
rect 183277 390690 183343 390693
rect 184933 390690 184999 390693
rect 112670 390688 184999 390690
rect 112670 390632 183282 390688
rect 183338 390632 184938 390688
rect 184994 390632 184999 390688
rect 112670 390630 184999 390632
rect 88996 390628 89002 390630
rect 89713 390627 89779 390630
rect 183277 390627 183343 390630
rect 184933 390627 184999 390630
rect 111742 390492 111748 390556
rect 111812 390554 111818 390556
rect 111977 390554 112043 390557
rect 111812 390552 112043 390554
rect 111812 390496 111982 390552
rect 112038 390496 112043 390552
rect 111812 390494 112043 390496
rect 111812 390492 111818 390494
rect 111977 390491 112043 390494
rect 147489 390554 147555 390557
rect 187601 390554 187667 390557
rect 147489 390552 187667 390554
rect 147489 390496 147494 390552
rect 147550 390496 187606 390552
rect 187662 390496 187667 390552
rect 147489 390494 187667 390496
rect 147489 390491 147555 390494
rect 187601 390491 187667 390494
rect 289905 390554 289971 390557
rect 582741 390554 582807 390557
rect 289905 390552 582807 390554
rect 289905 390496 289910 390552
rect 289966 390496 582746 390552
rect 582802 390496 582807 390552
rect 289905 390494 582807 390496
rect 289905 390491 289971 390494
rect 582741 390491 582807 390494
rect 72417 390418 72483 390421
rect 77201 390420 77267 390421
rect 72734 390418 72740 390420
rect 72417 390416 72740 390418
rect 72417 390360 72422 390416
rect 72478 390360 72740 390416
rect 72417 390358 72740 390360
rect 72417 390355 72483 390358
rect 72734 390356 72740 390358
rect 72804 390356 72810 390420
rect 77150 390418 77156 390420
rect 77110 390358 77156 390418
rect 77220 390416 77267 390420
rect 77262 390360 77267 390416
rect 77150 390356 77156 390358
rect 77220 390356 77267 390360
rect 77201 390355 77267 390356
rect 100661 390420 100727 390421
rect 104249 390420 104315 390421
rect 100661 390416 100708 390420
rect 100772 390418 100778 390420
rect 104198 390418 104204 390420
rect 100661 390360 100666 390416
rect 100661 390356 100708 390360
rect 100772 390358 100818 390418
rect 104158 390358 104204 390418
rect 104268 390416 104315 390420
rect 104310 390360 104315 390416
rect 100772 390356 100778 390358
rect 104198 390356 104204 390358
rect 104268 390356 104315 390360
rect 104934 390356 104940 390420
rect 105004 390418 105010 390420
rect 105261 390418 105327 390421
rect 105004 390416 105327 390418
rect 105004 390360 105266 390416
rect 105322 390360 105327 390416
rect 105004 390358 105327 390360
rect 105004 390356 105010 390358
rect 100661 390355 100727 390356
rect 104249 390355 104315 390356
rect 105261 390355 105327 390358
rect 160369 390418 160435 390421
rect 161565 390418 161631 390421
rect 160369 390416 161631 390418
rect 160369 390360 160374 390416
rect 160430 390360 161570 390416
rect 161626 390360 161631 390416
rect 160369 390358 161631 390360
rect 160369 390355 160435 390358
rect 161565 390355 161631 390358
rect 79910 390084 79916 390148
rect 79980 390146 79986 390148
rect 80053 390146 80119 390149
rect 81295 390146 81361 390149
rect 79980 390144 81361 390146
rect 79980 390088 80058 390144
rect 80114 390088 81300 390144
rect 81356 390088 81361 390144
rect 79980 390086 81361 390088
rect 79980 390084 79986 390086
rect 80053 390083 80119 390086
rect 81295 390083 81361 390086
rect 108297 389874 108363 389877
rect 117405 389874 117471 389877
rect 108297 389872 117471 389874
rect 108297 389816 108302 389872
rect 108358 389816 117410 389872
rect 117466 389816 117471 389872
rect 108297 389814 117471 389816
rect 108297 389811 108363 389814
rect 117405 389811 117471 389814
rect 184933 389874 184999 389877
rect 194133 389874 194199 389877
rect 184933 389872 194199 389874
rect 184933 389816 184938 389872
rect 184994 389816 194138 389872
rect 194194 389816 194199 389872
rect 184933 389814 194199 389816
rect 184933 389811 184999 389814
rect 194133 389811 194199 389814
rect 240777 389874 240843 389877
rect 269389 389874 269455 389877
rect 240777 389872 269455 389874
rect 240777 389816 240782 389872
rect 240838 389816 269394 389872
rect 269450 389816 269455 389872
rect 240777 389814 269455 389816
rect 240777 389811 240843 389814
rect 269389 389811 269455 389814
rect 193121 389466 193187 389469
rect 212533 389466 212599 389469
rect 193121 389464 212599 389466
rect 193121 389408 193126 389464
rect 193182 389408 212538 389464
rect 212594 389408 212599 389464
rect 193121 389406 212599 389408
rect 193121 389403 193187 389406
rect 212533 389403 212599 389406
rect 72417 389330 72483 389333
rect 73654 389330 73660 389332
rect 72417 389328 73660 389330
rect 72417 389272 72422 389328
rect 72478 389272 73660 389328
rect 72417 389270 73660 389272
rect 72417 389267 72483 389270
rect 73654 389268 73660 389270
rect 73724 389268 73730 389332
rect 147489 389330 147555 389333
rect 89670 389328 147555 389330
rect 89670 389272 147494 389328
rect 147550 389272 147555 389328
rect 89670 389270 147555 389272
rect 39941 389194 40007 389197
rect 87965 389194 88031 389197
rect 89670 389194 89730 389270
rect 147489 389267 147555 389270
rect 182817 389330 182883 389333
rect 229645 389330 229711 389333
rect 182817 389328 229711 389330
rect 182817 389272 182822 389328
rect 182878 389272 229650 389328
rect 229706 389272 229711 389328
rect 182817 389270 229711 389272
rect 182817 389267 182883 389270
rect 229645 389267 229711 389270
rect 39941 389192 89730 389194
rect 39941 389136 39946 389192
rect 40002 389136 87970 389192
rect 88026 389136 89730 389192
rect 39941 389134 89730 389136
rect 98913 389194 98979 389197
rect 160369 389194 160435 389197
rect 161381 389194 161447 389197
rect 98913 389192 161447 389194
rect 98913 389136 98918 389192
rect 98974 389136 160374 389192
rect 160430 389136 161386 389192
rect 161442 389136 161447 389192
rect 98913 389134 161447 389136
rect 39941 389131 40007 389134
rect 87965 389131 88031 389134
rect 98913 389131 98979 389134
rect 160369 389131 160435 389134
rect 161381 389131 161447 389134
rect 204805 389194 204871 389197
rect 289905 389194 289971 389197
rect 204805 389192 289971 389194
rect 204805 389136 204810 389192
rect 204866 389136 289910 389192
rect 289966 389136 289971 389192
rect 204805 389134 289971 389136
rect 204805 389131 204871 389134
rect 289905 389131 289971 389134
rect 96889 389058 96955 389061
rect 97625 389058 97691 389061
rect 96889 389056 97691 389058
rect 96889 389000 96894 389056
rect 96950 389000 97630 389056
rect 97686 389000 97691 389056
rect 96889 388998 97691 389000
rect 96889 388995 96955 388998
rect 97625 388995 97691 388998
rect 244222 388996 244228 389060
rect 244292 389058 244298 389060
rect 244733 389058 244799 389061
rect 244292 389056 244799 389058
rect 244292 389000 244738 389056
rect 244794 389000 244799 389056
rect 244292 388998 244799 389000
rect 244292 388996 244298 388998
rect 244733 388995 244799 388998
rect 247769 389058 247835 389061
rect 248597 389058 248663 389061
rect 247769 389056 248663 389058
rect 247769 389000 247774 389056
rect 247830 389000 248602 389056
rect 248658 389000 248663 389056
rect 247769 388998 248663 389000
rect 247769 388995 247835 388998
rect 248597 388995 248663 388998
rect 249241 389058 249307 389061
rect 249517 389058 249583 389061
rect 262213 389058 262279 389061
rect 249241 389056 262279 389058
rect 249241 389000 249246 389056
rect 249302 389000 249522 389056
rect 249578 389000 262218 389056
rect 262274 389000 262279 389056
rect 249241 388998 262279 389000
rect 249241 388995 249307 388998
rect 249517 388995 249583 388998
rect 262213 388995 262279 388998
rect 90449 388922 90515 388925
rect 221549 388922 221615 388925
rect 90449 388920 221615 388922
rect 90449 388864 90454 388920
rect 90510 388864 221554 388920
rect 221610 388864 221615 388920
rect 90449 388862 221615 388864
rect 90449 388859 90515 388862
rect 221549 388859 221615 388862
rect 77201 388786 77267 388789
rect 204805 388786 204871 388789
rect 77201 388784 204871 388786
rect 77201 388728 77206 388784
rect 77262 388728 204810 388784
rect 204866 388728 204871 388784
rect 77201 388726 204871 388728
rect 77201 388723 77267 388726
rect 204805 388723 204871 388726
rect 105169 388650 105235 388653
rect 242893 388650 242959 388653
rect 105169 388648 242959 388650
rect 105169 388592 105174 388648
rect 105230 388592 242898 388648
rect 242954 388592 242959 388648
rect 105169 388590 242959 388592
rect 105169 388587 105235 388590
rect 242893 388587 242959 388590
rect 77477 388514 77543 388517
rect 78438 388514 78444 388516
rect 77477 388512 78444 388514
rect 77477 388456 77482 388512
rect 77538 388456 78444 388512
rect 77477 388454 78444 388456
rect 77477 388451 77543 388454
rect 78438 388452 78444 388454
rect 78508 388452 78514 388516
rect 251030 388452 251036 388516
rect 251100 388514 251106 388516
rect 254209 388514 254275 388517
rect 251100 388512 254275 388514
rect 251100 388456 254214 388512
rect 254270 388456 254275 388512
rect 251100 388454 254275 388456
rect 251100 388452 251106 388454
rect 254209 388451 254275 388454
rect 254209 388106 254275 388109
rect 254710 388106 254716 388108
rect 254209 388104 254716 388106
rect 254209 388048 254214 388104
rect 254270 388048 254716 388104
rect 254209 388046 254716 388048
rect 254209 388043 254275 388046
rect 254710 388044 254716 388046
rect 254780 388044 254786 388108
rect 99465 387970 99531 387973
rect 100150 387970 100156 387972
rect 99465 387968 100156 387970
rect 99465 387912 99470 387968
rect 99526 387912 100156 387968
rect 99465 387910 100156 387912
rect 99465 387907 99531 387910
rect 100150 387908 100156 387910
rect 100220 387908 100226 387972
rect 50797 387698 50863 387701
rect 50981 387698 51047 387701
rect 155677 387698 155743 387701
rect 50797 387696 155743 387698
rect 50797 387640 50802 387696
rect 50858 387640 50986 387696
rect 51042 387640 155682 387696
rect 155738 387640 155743 387696
rect 50797 387638 155743 387640
rect 50797 387635 50863 387638
rect 50981 387635 51047 387638
rect 155677 387635 155743 387638
rect 173617 387698 173683 387701
rect 198181 387698 198247 387701
rect 265157 387698 265223 387701
rect 265709 387698 265775 387701
rect 173617 387696 265775 387698
rect 173617 387640 173622 387696
rect 173678 387640 198186 387696
rect 198242 387640 265162 387696
rect 265218 387640 265714 387696
rect 265770 387640 265775 387696
rect 173617 387638 265775 387640
rect 173617 387635 173683 387638
rect 198181 387635 198247 387638
rect 265157 387635 265223 387638
rect 265709 387635 265775 387638
rect 82721 387562 82787 387565
rect 84694 387562 84700 387564
rect 82721 387560 84700 387562
rect 82721 387504 82726 387560
rect 82782 387504 84700 387560
rect 82721 387502 84700 387504
rect 82721 387499 82787 387502
rect 84694 387500 84700 387502
rect 84764 387500 84770 387564
rect 93393 387562 93459 387565
rect 122833 387562 122899 387565
rect 123477 387562 123543 387565
rect 93393 387560 123543 387562
rect 93393 387504 93398 387560
rect 93454 387504 122838 387560
rect 122894 387504 123482 387560
rect 123538 387504 123543 387560
rect 93393 387502 123543 387504
rect 93393 387499 93459 387502
rect 122833 387499 122899 387502
rect 123477 387499 123543 387502
rect 179137 387562 179203 387565
rect 232589 387562 232655 387565
rect 179137 387560 232655 387562
rect 179137 387504 179142 387560
rect 179198 387504 232594 387560
rect 232650 387504 232655 387560
rect 179137 387502 232655 387504
rect 179137 387499 179203 387502
rect 232589 387499 232655 387502
rect 190177 387426 190243 387429
rect 191097 387426 191163 387429
rect 190177 387424 191163 387426
rect 190177 387368 190182 387424
rect 190238 387368 191102 387424
rect 191158 387368 191163 387424
rect 190177 387366 191163 387368
rect 190177 387363 190243 387366
rect 191097 387363 191163 387366
rect 73061 387018 73127 387021
rect 78254 387018 78260 387020
rect 73061 387016 78260 387018
rect 73061 386960 73066 387016
rect 73122 386960 78260 387016
rect 73061 386958 78260 386960
rect 73061 386955 73127 386958
rect 78254 386956 78260 386958
rect 78324 386956 78330 387020
rect 155677 387018 155743 387021
rect 187049 387018 187115 387021
rect 155677 387016 187115 387018
rect 155677 386960 155682 387016
rect 155738 386960 187054 387016
rect 187110 386960 187115 387016
rect 155677 386958 187115 386960
rect 155677 386955 155743 386958
rect 187049 386955 187115 386958
rect 78765 386882 78831 386885
rect 87454 386882 87460 386884
rect 78765 386880 87460 386882
rect 78765 386824 78770 386880
rect 78826 386824 87460 386880
rect 78765 386822 87460 386824
rect 78765 386819 78831 386822
rect 87454 386820 87460 386822
rect 87524 386820 87530 386884
rect 167729 386338 167795 386341
rect 201125 386338 201191 386341
rect 167729 386336 201191 386338
rect 167729 386280 167734 386336
rect 167790 386280 201130 386336
rect 201186 386280 201191 386336
rect 167729 386278 201191 386280
rect 167729 386275 167795 386278
rect 201125 386275 201191 386278
rect 224953 386338 225019 386341
rect 225781 386338 225847 386341
rect 277853 386338 277919 386341
rect 224953 386336 277919 386338
rect 224953 386280 224958 386336
rect 225014 386280 225786 386336
rect 225842 386280 277858 386336
rect 277914 386280 277919 386336
rect 224953 386278 277919 386280
rect 224953 386275 225019 386278
rect 225781 386275 225847 386278
rect 277853 386275 277919 386278
rect 170489 386202 170555 386205
rect 170990 386202 170996 386204
rect 170489 386200 170996 386202
rect 170489 386144 170494 386200
rect 170550 386144 170996 386200
rect 170489 386142 170996 386144
rect 170489 386139 170555 386142
rect 170990 386140 170996 386142
rect 171060 386140 171066 386204
rect 171869 386202 171935 386205
rect 172237 386202 172303 386205
rect 187693 386202 187759 386205
rect 220077 386202 220143 386205
rect 171869 386200 180810 386202
rect 171869 386144 171874 386200
rect 171930 386144 172242 386200
rect 172298 386144 180810 386200
rect 171869 386142 180810 386144
rect 171869 386139 171935 386142
rect 172237 386139 172303 386142
rect 180750 386066 180810 386142
rect 187693 386200 220143 386202
rect 187693 386144 187698 386200
rect 187754 386144 220082 386200
rect 220138 386144 220143 386200
rect 187693 386142 220143 386144
rect 187693 386139 187759 386142
rect 220077 386139 220143 386142
rect 242893 386202 242959 386205
rect 266537 386202 266603 386205
rect 266997 386202 267063 386205
rect 242893 386200 267063 386202
rect 242893 386144 242898 386200
rect 242954 386144 266542 386200
rect 266598 386144 267002 386200
rect 267058 386144 267063 386200
rect 242893 386142 267063 386144
rect 242893 386139 242959 386142
rect 266537 386139 266603 386142
rect 266997 386139 267063 386142
rect 200205 386066 200271 386069
rect 180750 386064 200271 386066
rect 180750 386008 200210 386064
rect 200266 386008 200271 386064
rect 180750 386006 200271 386008
rect 200205 386003 200271 386006
rect 89621 385930 89687 385933
rect 100886 385930 100892 385932
rect 89621 385928 100892 385930
rect 89621 385872 89626 385928
rect 89682 385872 100892 385928
rect 89621 385870 100892 385872
rect 89621 385867 89687 385870
rect 100886 385868 100892 385870
rect 100956 385868 100962 385932
rect 80881 385794 80947 385797
rect 110505 385794 110571 385797
rect 116209 385794 116275 385797
rect 80881 385792 116275 385794
rect 80881 385736 80886 385792
rect 80942 385736 110510 385792
rect 110566 385736 116214 385792
rect 116270 385736 116275 385792
rect 80881 385734 116275 385736
rect 80881 385731 80947 385734
rect 110505 385731 110571 385734
rect 116209 385731 116275 385734
rect 66662 385596 66668 385660
rect 66732 385658 66738 385660
rect 188981 385658 189047 385661
rect 66732 385656 189047 385658
rect 66732 385600 188986 385656
rect 189042 385600 189047 385656
rect 66732 385598 189047 385600
rect 66732 385596 66738 385598
rect 188981 385595 189047 385598
rect 213177 385658 213243 385661
rect 224953 385658 225019 385661
rect 213177 385656 225019 385658
rect 213177 385600 213182 385656
rect 213238 385600 224958 385656
rect 225014 385600 225019 385656
rect 213177 385598 225019 385600
rect 213177 385595 213243 385598
rect 224953 385595 225019 385598
rect 271086 385596 271092 385660
rect 271156 385658 271162 385660
rect 283005 385658 283071 385661
rect 271156 385656 283071 385658
rect 271156 385600 283010 385656
rect 283066 385600 283071 385656
rect 271156 385598 283071 385600
rect 271156 385596 271162 385598
rect 283005 385595 283071 385598
rect 78581 385114 78647 385117
rect 85798 385114 85804 385116
rect 78581 385112 85804 385114
rect 78581 385056 78586 385112
rect 78642 385056 85804 385112
rect 78581 385054 85804 385056
rect 78581 385051 78647 385054
rect 85798 385052 85804 385054
rect 85868 385052 85874 385116
rect 79409 384978 79475 384981
rect 129733 384978 129799 384981
rect 79409 384976 129799 384978
rect 79409 384920 79414 384976
rect 79470 384920 129738 384976
rect 129794 384920 129799 384976
rect 79409 384918 129799 384920
rect 79409 384915 79475 384918
rect 129733 384915 129799 384918
rect 163865 384978 163931 384981
rect 164877 384978 164943 384981
rect 163865 384976 164943 384978
rect 163865 384920 163870 384976
rect 163926 384920 164882 384976
rect 164938 384920 164943 384976
rect 163865 384918 164943 384920
rect 163865 384915 163931 384918
rect 164877 384915 164943 384918
rect 247677 384978 247743 384981
rect 291193 384978 291259 384981
rect 247677 384976 291259 384978
rect 247677 384920 247682 384976
rect 247738 384920 291198 384976
rect 291254 384920 291259 384976
rect 247677 384918 291259 384920
rect 247677 384915 247743 384918
rect 291193 384915 291259 384918
rect 259269 384842 259335 384845
rect 248370 384840 259335 384842
rect 248370 384784 259274 384840
rect 259330 384784 259335 384840
rect 248370 384782 259335 384784
rect -960 384284 480 384524
rect 154297 384434 154363 384437
rect 187550 384434 187556 384436
rect 154297 384432 187556 384434
rect 154297 384376 154302 384432
rect 154358 384376 187556 384432
rect 154297 384374 187556 384376
rect 154297 384371 154363 384374
rect 187550 384372 187556 384374
rect 187620 384372 187626 384436
rect 190269 384434 190335 384437
rect 198825 384434 198891 384437
rect 190269 384432 198891 384434
rect 190269 384376 190274 384432
rect 190330 384376 198830 384432
rect 198886 384376 198891 384432
rect 190269 384374 198891 384376
rect 190269 384371 190335 384374
rect 198825 384371 198891 384374
rect 235349 384434 235415 384437
rect 244365 384434 244431 384437
rect 235349 384432 244431 384434
rect 235349 384376 235354 384432
rect 235410 384376 244370 384432
rect 244426 384376 244431 384432
rect 235349 384374 244431 384376
rect 235349 384371 235415 384374
rect 244365 384371 244431 384374
rect 91093 384298 91159 384301
rect 163865 384298 163931 384301
rect 91093 384296 163931 384298
rect 91093 384240 91098 384296
rect 91154 384240 163870 384296
rect 163926 384240 163931 384296
rect 91093 384238 163931 384240
rect 91093 384235 91159 384238
rect 163865 384235 163931 384238
rect 180149 384298 180215 384301
rect 213453 384298 213519 384301
rect 180149 384296 213519 384298
rect 180149 384240 180154 384296
rect 180210 384240 213458 384296
rect 213514 384240 213519 384296
rect 180149 384238 213519 384240
rect 180149 384235 180215 384238
rect 213453 384235 213519 384238
rect 218789 384298 218855 384301
rect 239029 384298 239095 384301
rect 248370 384298 248430 384782
rect 259269 384779 259335 384782
rect 218789 384296 248430 384298
rect 218789 384240 218794 384296
rect 218850 384240 239034 384296
rect 239090 384240 248430 384296
rect 218789 384238 248430 384240
rect 218789 384235 218855 384238
rect 239029 384235 239095 384238
rect 71681 383618 71747 383621
rect 171041 383618 171107 383621
rect 198733 383618 198799 383621
rect 71681 383616 198799 383618
rect 71681 383560 71686 383616
rect 71742 383560 171046 383616
rect 171102 383560 198738 383616
rect 198794 383560 198799 383616
rect 71681 383558 198799 383560
rect 71681 383555 71747 383558
rect 171041 383555 171107 383558
rect 198733 383555 198799 383558
rect 70485 383482 70551 383485
rect 119337 383482 119403 383485
rect 70485 383480 119403 383482
rect 70485 383424 70490 383480
rect 70546 383424 119342 383480
rect 119398 383424 119403 383480
rect 70485 383422 119403 383424
rect 70485 383419 70551 383422
rect 119337 383419 119403 383422
rect 186957 383074 187023 383077
rect 244273 383074 244339 383077
rect 259545 383074 259611 383077
rect 186957 383072 259611 383074
rect 186957 383016 186962 383072
rect 187018 383016 244278 383072
rect 244334 383016 259550 383072
rect 259606 383016 259611 383072
rect 186957 383014 259611 383016
rect 186957 383011 187023 383014
rect 244273 383011 244339 383014
rect 259545 383011 259611 383014
rect 73797 382938 73863 382941
rect 80094 382938 80100 382940
rect 73797 382936 80100 382938
rect 73797 382880 73802 382936
rect 73858 382880 80100 382936
rect 73797 382878 80100 382880
rect 73797 382875 73863 382878
rect 80094 382876 80100 382878
rect 80164 382876 80170 382940
rect 86861 382938 86927 382941
rect 94446 382938 94452 382940
rect 86861 382936 94452 382938
rect 86861 382880 86866 382936
rect 86922 382880 94452 382936
rect 86861 382878 94452 382880
rect 86861 382875 86927 382878
rect 94446 382876 94452 382878
rect 94516 382876 94522 382940
rect 103329 382938 103395 382941
rect 114502 382938 114508 382940
rect 103329 382936 114508 382938
rect 103329 382880 103334 382936
rect 103390 382880 114508 382936
rect 103329 382878 114508 382880
rect 103329 382875 103395 382878
rect 114502 382876 114508 382878
rect 114572 382876 114578 382940
rect 198733 382938 198799 382941
rect 276105 382938 276171 382941
rect 198733 382936 276171 382938
rect 198733 382880 198738 382936
rect 198794 382880 276110 382936
rect 276166 382880 276171 382936
rect 198733 382878 276171 382880
rect 198733 382875 198799 382878
rect 276105 382875 276171 382878
rect 95141 382394 95207 382397
rect 102726 382394 102732 382396
rect 95141 382392 102732 382394
rect 95141 382336 95146 382392
rect 95202 382336 102732 382392
rect 95141 382334 102732 382336
rect 95141 382331 95207 382334
rect 102726 382332 102732 382334
rect 102796 382332 102802 382396
rect 177665 382394 177731 382397
rect 180006 382394 180012 382396
rect 177665 382392 180012 382394
rect 177665 382336 177670 382392
rect 177726 382336 180012 382392
rect 177665 382334 180012 382336
rect 177665 382331 177731 382334
rect 180006 382332 180012 382334
rect 180076 382332 180082 382396
rect 85573 382258 85639 382261
rect 139301 382258 139367 382261
rect 85573 382256 139367 382258
rect 85573 382200 85578 382256
rect 85634 382200 139306 382256
rect 139362 382200 139367 382256
rect 85573 382198 139367 382200
rect 85573 382195 85639 382198
rect 139301 382195 139367 382198
rect 187550 382196 187556 382260
rect 187620 382258 187626 382260
rect 291377 382258 291443 382261
rect 187620 382256 291443 382258
rect 187620 382200 291382 382256
rect 291438 382200 291443 382256
rect 187620 382198 291443 382200
rect 187620 382196 187626 382198
rect 291377 382195 291443 382198
rect 139301 381714 139367 381717
rect 173617 381714 173683 381717
rect 139301 381712 173683 381714
rect 139301 381656 139306 381712
rect 139362 381656 173622 381712
rect 173678 381656 173683 381712
rect 139301 381654 173683 381656
rect 139301 381651 139367 381654
rect 173617 381651 173683 381654
rect 218329 381714 218395 381717
rect 248454 381714 248460 381716
rect 218329 381712 248460 381714
rect 218329 381656 218334 381712
rect 218390 381656 248460 381712
rect 218329 381654 248460 381656
rect 218329 381651 218395 381654
rect 248454 381652 248460 381654
rect 248524 381652 248530 381716
rect 148317 381578 148383 381581
rect 227805 381578 227871 381581
rect 148317 381576 227871 381578
rect 148317 381520 148322 381576
rect 148378 381520 227810 381576
rect 227866 381520 227871 381576
rect 148317 381518 227871 381520
rect 148317 381515 148383 381518
rect 227805 381515 227871 381518
rect 107745 380898 107811 380901
rect 247677 380898 247743 380901
rect 107745 380896 247743 380898
rect 107745 380840 107750 380896
rect 107806 380840 247682 380896
rect 247738 380840 247743 380896
rect 107745 380838 247743 380840
rect 107745 380835 107811 380838
rect 247677 380835 247743 380838
rect 180241 380762 180307 380765
rect 280286 380762 280292 380764
rect 180241 380760 280292 380762
rect 180241 380704 180246 380760
rect 180302 380704 280292 380760
rect 180241 380702 280292 380704
rect 180241 380699 180307 380702
rect 280286 380700 280292 380702
rect 280356 380762 280362 380764
rect 280429 380762 280495 380765
rect 280356 380760 280495 380762
rect 280356 380704 280434 380760
rect 280490 380704 280495 380760
rect 280356 380702 280495 380704
rect 280356 380700 280362 380702
rect 280429 380699 280495 380702
rect 105997 379402 106063 379405
rect 243077 379402 243143 379405
rect 105997 379400 243143 379402
rect 105997 379344 106002 379400
rect 106058 379344 243082 379400
rect 243138 379344 243143 379400
rect 105997 379342 243143 379344
rect 105997 379339 106063 379342
rect 243077 379339 243143 379342
rect 173157 379266 173223 379269
rect 273437 379266 273503 379269
rect 173157 379264 273503 379266
rect 173157 379208 173162 379264
rect 173218 379208 273442 379264
rect 273498 379208 273503 379264
rect 173157 379206 273503 379208
rect 173157 379203 173223 379206
rect 273437 379203 273503 379206
rect 273294 378932 273300 378996
rect 273364 378994 273370 378996
rect 273437 378994 273503 378997
rect 273364 378992 273503 378994
rect 273364 378936 273442 378992
rect 273498 378936 273503 378992
rect 273364 378934 273503 378936
rect 273364 378932 273370 378934
rect 273437 378931 273503 378934
rect 80697 378722 80763 378725
rect 122925 378722 122991 378725
rect 80697 378720 122991 378722
rect 80697 378664 80702 378720
rect 80758 378664 122930 378720
rect 122986 378664 122991 378720
rect 80697 378662 122991 378664
rect 80697 378659 80763 378662
rect 122925 378659 122991 378662
rect 192702 378660 192708 378724
rect 192772 378722 192778 378724
rect 212625 378722 212691 378725
rect 192772 378720 212691 378722
rect 192772 378664 212630 378720
rect 212686 378664 212691 378720
rect 192772 378662 212691 378664
rect 192772 378660 192778 378662
rect 212625 378659 212691 378662
rect 582373 378450 582439 378453
rect 583520 378450 584960 378540
rect 582373 378448 584960 378450
rect 582373 378392 582378 378448
rect 582434 378392 584960 378448
rect 582373 378390 584960 378392
rect 582373 378387 582439 378390
rect 583520 378300 584960 378390
rect 188981 378178 189047 378181
rect 188981 378176 189090 378178
rect 188981 378120 188986 378176
rect 189042 378120 189090 378176
rect 188981 378115 189090 378120
rect 144269 378042 144335 378045
rect 144729 378042 144795 378045
rect 189030 378042 189090 378115
rect 288382 378042 288388 378044
rect 144269 378040 151830 378042
rect 144269 377984 144274 378040
rect 144330 377984 144734 378040
rect 144790 377984 151830 378040
rect 144269 377982 151830 377984
rect 189030 377982 288388 378042
rect 144269 377979 144335 377982
rect 144729 377979 144795 377982
rect 151770 377906 151830 377982
rect 288382 377980 288388 377982
rect 288452 378042 288458 378044
rect 288617 378042 288683 378045
rect 288452 378040 288683 378042
rect 288452 377984 288622 378040
rect 288678 377984 288683 378040
rect 288452 377982 288683 377984
rect 288452 377980 288458 377982
rect 288617 377979 288683 377982
rect 220721 377906 220787 377909
rect 151770 377904 220787 377906
rect 151770 377848 220726 377904
rect 220782 377848 220787 377904
rect 151770 377846 220787 377848
rect 220721 377843 220787 377846
rect 69606 377436 69612 377500
rect 69676 377498 69682 377500
rect 97257 377498 97323 377501
rect 69676 377496 97323 377498
rect 69676 377440 97262 377496
rect 97318 377440 97323 377496
rect 69676 377438 97323 377440
rect 69676 377436 69682 377438
rect 97257 377435 97323 377438
rect 3417 377362 3483 377365
rect 119981 377362 120047 377365
rect 3417 377360 120047 377362
rect 3417 377304 3422 377360
rect 3478 377304 119986 377360
rect 120042 377304 120047 377360
rect 3417 377302 120047 377304
rect 3417 377299 3483 377302
rect 119981 377299 120047 377302
rect 228449 377362 228515 377365
rect 241646 377362 241652 377364
rect 228449 377360 241652 377362
rect 228449 377304 228454 377360
rect 228510 377304 241652 377360
rect 228449 377302 241652 377304
rect 228449 377299 228515 377302
rect 241646 377300 241652 377302
rect 241716 377300 241722 377364
rect 124949 376682 125015 376685
rect 276013 376682 276079 376685
rect 276422 376682 276428 376684
rect 124949 376680 276428 376682
rect 124949 376624 124954 376680
rect 125010 376624 276018 376680
rect 276074 376624 276428 376680
rect 124949 376622 276428 376624
rect 124949 376619 125015 376622
rect 276013 376619 276079 376622
rect 276422 376620 276428 376622
rect 276492 376620 276498 376684
rect 67633 376546 67699 376549
rect 161473 376546 161539 376549
rect 162117 376546 162183 376549
rect 67633 376544 162183 376546
rect 67633 376488 67638 376544
rect 67694 376488 161478 376544
rect 161534 376488 162122 376544
rect 162178 376488 162183 376544
rect 67633 376486 162183 376488
rect 67633 376483 67699 376486
rect 161473 376483 161539 376486
rect 162117 376483 162183 376486
rect 189717 376546 189783 376549
rect 190177 376546 190243 376549
rect 291469 376546 291535 376549
rect 189717 376544 291535 376546
rect 189717 376488 189722 376544
rect 189778 376488 190182 376544
rect 190238 376488 291474 376544
rect 291530 376488 291535 376544
rect 189717 376486 291535 376488
rect 189717 376483 189783 376486
rect 190177 376483 190243 376486
rect 291469 376483 291535 376486
rect 81985 376410 82051 376413
rect 149697 376410 149763 376413
rect 81985 376408 149763 376410
rect 81985 376352 81990 376408
rect 82046 376352 149702 376408
rect 149758 376352 149763 376408
rect 81985 376350 149763 376352
rect 81985 376347 82051 376350
rect 149697 376347 149763 376350
rect 64597 375322 64663 375325
rect 188337 375322 188403 375325
rect 253933 375322 253999 375325
rect 254117 375322 254183 375325
rect 64597 375320 188403 375322
rect 64597 375264 64602 375320
rect 64658 375264 188342 375320
rect 188398 375264 188403 375320
rect 64597 375262 188403 375264
rect 64597 375259 64663 375262
rect 188337 375259 188403 375262
rect 238710 375320 254183 375322
rect 238710 375264 253938 375320
rect 253994 375264 254122 375320
rect 254178 375264 254183 375320
rect 238710 375262 254183 375264
rect 141417 375186 141483 375189
rect 238710 375186 238770 375262
rect 253933 375259 253999 375262
rect 254117 375259 254183 375262
rect 141417 375184 238770 375186
rect 141417 375128 141422 375184
rect 141478 375128 238770 375184
rect 141417 375126 238770 375128
rect 141417 375123 141483 375126
rect 184289 373962 184355 373965
rect 245653 373962 245719 373965
rect 184289 373960 245719 373962
rect 184289 373904 184294 373960
rect 184350 373904 245658 373960
rect 245714 373904 245719 373960
rect 184289 373902 245719 373904
rect 184289 373899 184355 373902
rect 245653 373899 245719 373902
rect 88333 373282 88399 373285
rect 137369 373282 137435 373285
rect 144269 373282 144335 373285
rect 88333 373280 144335 373282
rect 88333 373224 88338 373280
rect 88394 373224 137374 373280
rect 137430 373224 144274 373280
rect 144330 373224 144335 373280
rect 88333 373222 144335 373224
rect 88333 373219 88399 373222
rect 137369 373219 137435 373222
rect 144269 373219 144335 373222
rect 146937 373282 147003 373285
rect 188429 373282 188495 373285
rect 146937 373280 188495 373282
rect 146937 373224 146942 373280
rect 146998 373224 188434 373280
rect 188490 373224 188495 373280
rect 146937 373222 188495 373224
rect 146937 373219 147003 373222
rect 188429 373219 188495 373222
rect 208393 373282 208459 373285
rect 284293 373282 284359 373285
rect 208393 373280 284359 373282
rect 208393 373224 208398 373280
rect 208454 373224 284298 373280
rect 284354 373224 284359 373280
rect 208393 373222 284359 373224
rect 208393 373219 208459 373222
rect 284293 373219 284359 373222
rect 245653 372738 245719 372741
rect 246297 372738 246363 372741
rect 245653 372736 246363 372738
rect 245653 372680 245658 372736
rect 245714 372680 246302 372736
rect 246358 372680 246363 372736
rect 245653 372678 246363 372680
rect 245653 372675 245719 372678
rect 246297 372675 246363 372678
rect 109677 371922 109743 371925
rect 249241 371922 249307 371925
rect 249609 371922 249675 371925
rect 109677 371920 249675 371922
rect 109677 371864 109682 371920
rect 109738 371864 249246 371920
rect 249302 371864 249614 371920
rect 249670 371864 249675 371920
rect 109677 371862 249675 371864
rect 109677 371859 109743 371862
rect 249241 371859 249307 371862
rect 249609 371859 249675 371862
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 109033 371378 109099 371381
rect 109677 371378 109743 371381
rect 109033 371376 109743 371378
rect 109033 371320 109038 371376
rect 109094 371320 109682 371376
rect 109738 371320 109743 371376
rect 109033 371318 109743 371320
rect 109033 371315 109099 371318
rect 109677 371315 109743 371318
rect 73153 371242 73219 371245
rect 167729 371242 167795 371245
rect 73153 371240 167795 371242
rect 73153 371184 73158 371240
rect 73214 371184 167734 371240
rect 167790 371184 167795 371240
rect 73153 371182 167795 371184
rect 73153 371179 73219 371182
rect 167729 371179 167795 371182
rect 99281 370562 99347 370565
rect 111006 370562 111012 370564
rect 99281 370560 111012 370562
rect 99281 370504 99286 370560
rect 99342 370504 111012 370560
rect 99281 370502 111012 370504
rect 99281 370499 99347 370502
rect 111006 370500 111012 370502
rect 111076 370500 111082 370564
rect 181478 370500 181484 370564
rect 181548 370562 181554 370564
rect 190453 370562 190519 370565
rect 181548 370560 190519 370562
rect 181548 370504 190458 370560
rect 190514 370504 190519 370560
rect 181548 370502 190519 370504
rect 181548 370500 181554 370502
rect 190453 370499 190519 370502
rect 166993 369882 167059 369885
rect 167729 369882 167795 369885
rect 166993 369880 167795 369882
rect 166993 369824 166998 369880
rect 167054 369824 167734 369880
rect 167790 369824 167795 369880
rect 166993 369822 167795 369824
rect 166993 369819 167059 369822
rect 167729 369819 167795 369822
rect 168189 369746 168255 369749
rect 171777 369746 171843 369749
rect 168189 369744 171843 369746
rect 168189 369688 168194 369744
rect 168250 369688 171782 369744
rect 171838 369688 171843 369744
rect 168189 369686 171843 369688
rect 168189 369683 168255 369686
rect 171777 369683 171843 369686
rect 77201 369204 77267 369205
rect 77150 369140 77156 369204
rect 77220 369202 77267 369204
rect 229737 369202 229803 369205
rect 267733 369202 267799 369205
rect 77220 369200 84210 369202
rect 77262 369144 84210 369200
rect 77220 369142 84210 369144
rect 77220 369140 77267 369142
rect 77201 369139 77267 369140
rect 84150 369066 84210 369142
rect 229737 369200 267799 369202
rect 229737 369144 229742 369200
rect 229798 369144 267738 369200
rect 267794 369144 267799 369200
rect 229737 369142 267799 369144
rect 229737 369139 229803 369142
rect 267733 369139 267799 369142
rect 137277 369066 137343 369069
rect 84150 369064 137343 369066
rect 84150 369008 137282 369064
rect 137338 369008 137343 369064
rect 84150 369006 137343 369008
rect 137277 369003 137343 369006
rect 209773 369066 209839 369069
rect 277485 369066 277551 369069
rect 209773 369064 277551 369066
rect 209773 369008 209778 369064
rect 209834 369008 277490 369064
rect 277546 369008 277551 369064
rect 209773 369006 277551 369008
rect 209773 369003 209839 369006
rect 277485 369003 277551 369006
rect 154389 368386 154455 368389
rect 267825 368386 267891 368389
rect 154389 368384 267891 368386
rect 154389 368328 154394 368384
rect 154450 368328 267830 368384
rect 267886 368328 267891 368384
rect 154389 368326 267891 368328
rect 154389 368323 154455 368326
rect 267825 368323 267891 368326
rect 156597 367026 156663 367029
rect 157241 367026 157307 367029
rect 252686 367026 252692 367028
rect 156597 367024 252692 367026
rect 156597 366968 156602 367024
rect 156658 366968 157246 367024
rect 157302 366968 252692 367024
rect 156597 366966 252692 366968
rect 156597 366963 156663 366966
rect 157241 366963 157307 366966
rect 252686 366964 252692 366966
rect 252756 366964 252762 367028
rect 170489 366890 170555 366893
rect 244365 366890 244431 366893
rect 170489 366888 248430 366890
rect 170489 366832 170494 366888
rect 170550 366832 244370 366888
rect 244426 366832 248430 366888
rect 170489 366830 248430 366832
rect 170489 366827 170555 366830
rect 244365 366827 244431 366830
rect 248370 366346 248430 366830
rect 258390 366346 258396 366348
rect 248370 366286 258396 366346
rect 258390 366284 258396 366286
rect 258460 366284 258466 366348
rect 67449 365666 67515 365669
rect 169017 365666 169083 365669
rect 67449 365664 169083 365666
rect 67449 365608 67454 365664
rect 67510 365608 169022 365664
rect 169078 365608 169083 365664
rect 67449 365606 169083 365608
rect 67449 365603 67515 365606
rect 169017 365603 169083 365606
rect 582465 365122 582531 365125
rect 583520 365122 584960 365212
rect 582465 365120 584960 365122
rect 582465 365064 582470 365120
rect 582526 365064 584960 365120
rect 582465 365062 584960 365064
rect 582465 365059 582531 365062
rect 222929 364986 222995 364989
rect 247718 364986 247724 364988
rect 222929 364984 247724 364986
rect 222929 364928 222934 364984
rect 222990 364928 247724 364984
rect 222929 364926 247724 364928
rect 222929 364923 222995 364926
rect 247718 364924 247724 364926
rect 247788 364924 247794 364988
rect 249609 364986 249675 364989
rect 270718 364986 270724 364988
rect 249609 364984 270724 364986
rect 249609 364928 249614 364984
rect 249670 364928 270724 364984
rect 249609 364926 270724 364928
rect 249609 364923 249675 364926
rect 270718 364924 270724 364926
rect 270788 364924 270794 364988
rect 583520 364972 584960 365062
rect 225597 363626 225663 363629
rect 262254 363626 262260 363628
rect 225597 363624 262260 363626
rect 225597 363568 225602 363624
rect 225658 363568 262260 363624
rect 225597 363566 262260 363568
rect 225597 363563 225663 363566
rect 262254 363564 262260 363566
rect 262324 363564 262330 363628
rect 188429 362946 188495 362949
rect 270769 362946 270835 362949
rect 188429 362944 270835 362946
rect 188429 362888 188434 362944
rect 188490 362888 270774 362944
rect 270830 362888 270835 362944
rect 188429 362886 270835 362888
rect 188429 362883 188495 362886
rect 270769 362883 270835 362886
rect 70393 362266 70459 362269
rect 71630 362266 71636 362268
rect 70393 362264 71636 362266
rect 70393 362208 70398 362264
rect 70454 362208 71636 362264
rect 70393 362206 71636 362208
rect 70393 362203 70459 362206
rect 71630 362204 71636 362206
rect 71700 362266 71706 362268
rect 195973 362266 196039 362269
rect 71700 362264 196039 362266
rect 71700 362208 195978 362264
rect 196034 362208 196039 362264
rect 71700 362206 196039 362208
rect 71700 362204 71706 362206
rect 195973 362203 196039 362206
rect 228541 362266 228607 362269
rect 242249 362266 242315 362269
rect 228541 362264 242315 362266
rect 228541 362208 228546 362264
rect 228602 362208 242254 362264
rect 242310 362208 242315 362264
rect 228541 362206 242315 362208
rect 228541 362203 228607 362206
rect 242249 362203 242315 362206
rect 246389 362266 246455 362269
rect 256734 362266 256740 362268
rect 246389 362264 256740 362266
rect 246389 362208 246394 362264
rect 246450 362208 256740 362264
rect 246389 362206 256740 362208
rect 246389 362203 246455 362206
rect 256734 362204 256740 362206
rect 256804 362204 256810 362268
rect 144177 361586 144243 361589
rect 251817 361586 251883 361589
rect 144177 361584 251883 361586
rect 144177 361528 144182 361584
rect 144238 361528 251822 361584
rect 251878 361528 251883 361584
rect 144177 361526 251883 361528
rect 144177 361523 144243 361526
rect 251817 361523 251883 361526
rect 211797 359410 211863 359413
rect 265065 359410 265131 359413
rect 211797 359408 265131 359410
rect 211797 359352 211802 359408
rect 211858 359352 265070 359408
rect 265126 359352 265131 359408
rect 211797 359350 265131 359352
rect 211797 359347 211863 359350
rect 265065 359347 265131 359350
rect 240041 359138 240107 359141
rect 245878 359138 245884 359140
rect 240041 359136 245884 359138
rect 240041 359080 240046 359136
rect 240102 359080 245884 359136
rect 240041 359078 245884 359080
rect 240041 359075 240107 359078
rect 245878 359076 245884 359078
rect 245948 359076 245954 359140
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 195237 358050 195303 358053
rect 271873 358050 271939 358053
rect 195237 358048 271939 358050
rect 195237 357992 195242 358048
rect 195298 357992 271878 358048
rect 271934 357992 271939 358048
rect 195237 357990 271939 357992
rect 195237 357987 195303 357990
rect 271873 357987 271939 357990
rect 238017 356826 238083 356829
rect 273478 356826 273484 356828
rect 238017 356824 273484 356826
rect 238017 356768 238022 356824
rect 238078 356768 273484 356824
rect 238017 356766 273484 356768
rect 238017 356763 238083 356766
rect 273478 356764 273484 356766
rect 273548 356764 273554 356828
rect 206369 356690 206435 356693
rect 259494 356690 259500 356692
rect 206369 356688 259500 356690
rect 206369 356632 206374 356688
rect 206430 356632 259500 356688
rect 206369 356630 259500 356632
rect 206369 356627 206435 356630
rect 259494 356628 259500 356630
rect 259564 356628 259570 356692
rect 217409 355330 217475 355333
rect 280102 355330 280108 355332
rect 217409 355328 280108 355330
rect 217409 355272 217414 355328
rect 217470 355272 280108 355328
rect 217409 355270 280108 355272
rect 217409 355267 217475 355270
rect 280102 355268 280108 355270
rect 280172 355268 280178 355332
rect 214557 353970 214623 353973
rect 257061 353970 257127 353973
rect 214557 353968 257127 353970
rect 214557 353912 214562 353968
rect 214618 353912 257066 353968
rect 257122 353912 257127 353968
rect 214557 353910 257127 353912
rect 214557 353907 214623 353910
rect 257061 353907 257127 353910
rect 162526 351868 162532 351932
rect 162596 351930 162602 351932
rect 169702 351930 169708 351932
rect 162596 351870 169708 351930
rect 162596 351868 162602 351870
rect 169702 351868 169708 351870
rect 169772 351868 169778 351932
rect 582557 351930 582623 351933
rect 583520 351930 584960 352020
rect 582557 351928 584960 351930
rect 582557 351872 582562 351928
rect 582618 351872 584960 351928
rect 582557 351870 584960 351872
rect 582557 351867 582623 351870
rect 226977 351794 227043 351797
rect 259453 351794 259519 351797
rect 263726 351794 263732 351796
rect 226977 351792 263732 351794
rect 226977 351736 226982 351792
rect 227038 351736 259458 351792
rect 259514 351736 263732 351792
rect 226977 351734 263732 351736
rect 226977 351731 227043 351734
rect 259453 351731 259519 351734
rect 263726 351732 263732 351734
rect 263796 351732 263802 351796
rect 583520 351780 584960 351870
rect 179086 351188 179092 351252
rect 179156 351250 179162 351252
rect 189809 351250 189875 351253
rect 179156 351248 189875 351250
rect 179156 351192 189814 351248
rect 189870 351192 189875 351248
rect 179156 351190 189875 351192
rect 179156 351188 179162 351190
rect 189809 351187 189875 351190
rect 183369 351114 183435 351117
rect 244222 351114 244228 351116
rect 183369 351112 244228 351114
rect 183369 351056 183374 351112
rect 183430 351056 244228 351112
rect 183369 351054 244228 351056
rect 183369 351051 183435 351054
rect 244222 351052 244228 351054
rect 244292 351052 244298 351116
rect 206277 349754 206343 349757
rect 262438 349754 262444 349756
rect 206277 349752 262444 349754
rect 206277 349696 206282 349752
rect 206338 349696 262444 349752
rect 206277 349694 262444 349696
rect 206277 349691 206343 349694
rect 262438 349692 262444 349694
rect 262508 349692 262514 349756
rect 151261 347850 151327 347853
rect 262305 347850 262371 347853
rect 151261 347848 262371 347850
rect 151261 347792 151266 347848
rect 151322 347792 262310 347848
rect 262366 347792 262371 347848
rect 151261 347790 262371 347792
rect 151261 347787 151327 347790
rect 262305 347787 262371 347790
rect 246297 347034 246363 347037
rect 260281 347034 260347 347037
rect 246297 347032 260347 347034
rect 246297 346976 246302 347032
rect 246358 346976 260286 347032
rect 260342 346976 260347 347032
rect 246297 346974 260347 346976
rect 246297 346971 246363 346974
rect 260281 346971 260347 346974
rect 82905 346490 82971 346493
rect 272057 346490 272123 346493
rect 82905 346488 272123 346490
rect 82905 346432 82910 346488
rect 82966 346432 272062 346488
rect 272118 346432 272123 346488
rect 82905 346430 272123 346432
rect 82905 346427 82971 346430
rect 272057 346427 272123 346430
rect 214373 345810 214439 345813
rect 267958 345810 267964 345812
rect 214373 345808 267964 345810
rect 214373 345752 214378 345808
rect 214434 345752 267964 345808
rect 214373 345750 267964 345752
rect 214373 345747 214439 345750
rect 267958 345748 267964 345750
rect 268028 345748 268034 345812
rect 184841 345674 184907 345677
rect 254526 345674 254532 345676
rect 184841 345672 254532 345674
rect 184841 345616 184846 345672
rect 184902 345616 254532 345672
rect 184841 345614 254532 345616
rect 184841 345611 184907 345614
rect 254526 345612 254532 345614
rect 254596 345612 254602 345676
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 217317 344314 217383 344317
rect 269062 344314 269068 344316
rect 217317 344312 269068 344314
rect 217317 344256 217322 344312
rect 217378 344256 269068 344312
rect 217317 344254 269068 344256
rect 217317 344251 217383 344254
rect 269062 344252 269068 344254
rect 269132 344252 269138 344316
rect 154481 343634 154547 343637
rect 175549 343634 175615 343637
rect 154481 343632 175615 343634
rect 154481 343576 154486 343632
rect 154542 343576 175554 343632
rect 175610 343576 175615 343632
rect 154481 343574 175615 343576
rect 154481 343571 154547 343574
rect 175549 343571 175615 343574
rect 224217 343090 224283 343093
rect 246389 343090 246455 343093
rect 224217 343088 246455 343090
rect 224217 343032 224222 343088
rect 224278 343032 246394 343088
rect 246450 343032 246455 343088
rect 224217 343030 246455 343032
rect 224217 343027 224283 343030
rect 246389 343027 246455 343030
rect 19333 342954 19399 342957
rect 154481 342954 154547 342957
rect 19333 342952 154547 342954
rect 19333 342896 19338 342952
rect 19394 342896 154486 342952
rect 154542 342896 154547 342952
rect 19333 342894 154547 342896
rect 19333 342891 19399 342894
rect 154481 342891 154547 342894
rect 177757 342954 177823 342957
rect 225597 342954 225663 342957
rect 177757 342952 225663 342954
rect 177757 342896 177762 342952
rect 177818 342896 225602 342952
rect 225658 342896 225663 342952
rect 177757 342894 225663 342896
rect 177757 342891 177823 342894
rect 225597 342891 225663 342894
rect 173566 341532 173572 341596
rect 173636 341594 173642 341596
rect 214373 341594 214439 341597
rect 173636 341592 214439 341594
rect 173636 341536 214378 341592
rect 214434 341536 214439 341592
rect 173636 341534 214439 341536
rect 173636 341532 173642 341534
rect 214373 341531 214439 341534
rect 163630 341396 163636 341460
rect 163700 341458 163706 341460
rect 171777 341458 171843 341461
rect 163700 341456 171843 341458
rect 163700 341400 171782 341456
rect 171838 341400 171843 341456
rect 163700 341398 171843 341400
rect 163700 341396 163706 341398
rect 171777 341395 171843 341398
rect 196617 341458 196683 341461
rect 260925 341458 260991 341461
rect 196617 341456 260991 341458
rect 196617 341400 196622 341456
rect 196678 341400 260930 341456
rect 260986 341400 260991 341456
rect 196617 341398 260991 341400
rect 196617 341395 196683 341398
rect 260925 341395 260991 341398
rect 268009 341458 268075 341461
rect 268326 341458 268332 341460
rect 268009 341456 268332 341458
rect 268009 341400 268014 341456
rect 268070 341400 268332 341456
rect 268009 341398 268332 341400
rect 268009 341395 268075 341398
rect 268326 341396 268332 341398
rect 268396 341396 268402 341460
rect 160686 339492 160692 339556
rect 160756 339554 160762 339556
rect 161238 339554 161244 339556
rect 160756 339494 161244 339554
rect 160756 339492 160762 339494
rect 161238 339492 161244 339494
rect 161308 339554 161314 339556
rect 226977 339554 227043 339557
rect 161308 339552 227043 339554
rect 161308 339496 226982 339552
rect 227038 339496 227043 339552
rect 161308 339494 227043 339496
rect 161308 339492 161314 339494
rect 226977 339491 227043 339494
rect 154021 338738 154087 338741
rect 190545 338738 190611 338741
rect 191741 338738 191807 338741
rect 154021 338736 191807 338738
rect 154021 338680 154026 338736
rect 154082 338680 190550 338736
rect 190606 338680 191746 338736
rect 191802 338680 191807 338736
rect 154021 338678 191807 338680
rect 154021 338675 154087 338678
rect 190545 338675 190611 338678
rect 191741 338675 191807 338678
rect 200757 338738 200823 338741
rect 293953 338738 294019 338741
rect 200757 338736 294019 338738
rect 200757 338680 200762 338736
rect 200818 338680 293958 338736
rect 294014 338680 294019 338736
rect 200757 338678 294019 338680
rect 200757 338675 200823 338678
rect 293953 338675 294019 338678
rect 583520 338452 584960 338692
rect 41321 337378 41387 337381
rect 173750 337378 173756 337380
rect 41321 337376 173756 337378
rect 41321 337320 41326 337376
rect 41382 337320 173756 337376
rect 41321 337318 173756 337320
rect 41321 337315 41387 337318
rect 173750 337316 173756 337318
rect 173820 337378 173826 337380
rect 224953 337378 225019 337381
rect 173820 337376 225019 337378
rect 173820 337320 224958 337376
rect 225014 337320 225019 337376
rect 173820 337318 225019 337320
rect 173820 337316 173826 337318
rect 224953 337315 225019 337318
rect 225137 337378 225203 337381
rect 245694 337378 245700 337380
rect 225137 337376 245700 337378
rect 225137 337320 225142 337376
rect 225198 337320 245700 337376
rect 225137 337318 245700 337320
rect 225137 337315 225203 337318
rect 245694 337316 245700 337318
rect 245764 337316 245770 337380
rect 156638 336228 156644 336292
rect 156708 336290 156714 336292
rect 201677 336290 201743 336293
rect 156708 336288 201743 336290
rect 156708 336232 201682 336288
rect 201738 336232 201743 336288
rect 156708 336230 201743 336232
rect 156708 336228 156714 336230
rect 201677 336227 201743 336230
rect 141366 336092 141372 336156
rect 141436 336154 141442 336156
rect 165521 336154 165587 336157
rect 141436 336152 165587 336154
rect 141436 336096 165526 336152
rect 165582 336096 165587 336152
rect 141436 336094 165587 336096
rect 141436 336092 141442 336094
rect 165521 336091 165587 336094
rect 8293 336018 8359 336021
rect 156638 336018 156644 336020
rect 8293 336016 156644 336018
rect 8293 335960 8298 336016
rect 8354 335960 156644 336016
rect 8293 335958 156644 335960
rect 8293 335955 8359 335958
rect 156638 335956 156644 335958
rect 156708 335956 156714 336020
rect 191741 336018 191807 336021
rect 266445 336018 266511 336021
rect 191741 336016 266511 336018
rect 191741 335960 191746 336016
rect 191802 335960 266450 336016
rect 266506 335960 266511 336016
rect 191741 335958 266511 335960
rect 191741 335955 191807 335958
rect 266445 335955 266511 335958
rect 153193 335474 153259 335477
rect 225137 335474 225203 335477
rect 153193 335472 225203 335474
rect 153193 335416 153198 335472
rect 153254 335416 225142 335472
rect 225198 335416 225203 335472
rect 153193 335414 225203 335416
rect 153193 335411 153259 335414
rect 225137 335411 225203 335414
rect 130469 334794 130535 334797
rect 190453 334794 190519 334797
rect 213913 334794 213979 334797
rect 130469 334792 213979 334794
rect 130469 334736 130474 334792
rect 130530 334736 190458 334792
rect 190514 334736 213918 334792
rect 213974 334736 213979 334792
rect 130469 334734 213979 334736
rect 130469 334731 130535 334734
rect 190453 334731 190519 334734
rect 213913 334731 213979 334734
rect 12433 334658 12499 334661
rect 158478 334658 158484 334660
rect 12433 334656 158484 334658
rect 12433 334600 12438 334656
rect 12494 334600 158484 334656
rect 12433 334598 158484 334600
rect 12433 334595 12499 334598
rect 158478 334596 158484 334598
rect 158548 334658 158554 334660
rect 219433 334658 219499 334661
rect 158548 334656 219499 334658
rect 158548 334600 219438 334656
rect 219494 334600 219499 334656
rect 158548 334598 219499 334600
rect 158548 334596 158554 334598
rect 219433 334595 219499 334598
rect 222101 334658 222167 334661
rect 242934 334658 242940 334660
rect 222101 334656 242940 334658
rect 222101 334600 222106 334656
rect 222162 334600 242940 334656
rect 222101 334598 242940 334600
rect 222101 334595 222167 334598
rect 242934 334596 242940 334598
rect 243004 334596 243010 334660
rect 253197 334658 253263 334661
rect 267958 334658 267964 334660
rect 253197 334656 267964 334658
rect 253197 334600 253202 334656
rect 253258 334600 267964 334656
rect 253197 334598 267964 334600
rect 253197 334595 253263 334598
rect 267958 334596 267964 334598
rect 268028 334596 268034 334660
rect 267733 334116 267799 334117
rect 267733 334112 267780 334116
rect 267844 334114 267850 334116
rect 267733 334056 267738 334112
rect 267733 334052 267780 334056
rect 267844 334054 267890 334114
rect 267844 334052 267850 334054
rect 267733 334051 267799 334052
rect 149697 333434 149763 333437
rect 159766 333434 159772 333436
rect 149697 333432 159772 333434
rect 149697 333376 149702 333432
rect 149758 333376 159772 333432
rect 149697 333374 159772 333376
rect 149697 333371 149763 333374
rect 159766 333372 159772 333374
rect 159836 333434 159842 333436
rect 207289 333434 207355 333437
rect 159836 333432 207355 333434
rect 159836 333376 207294 333432
rect 207350 333376 207355 333432
rect 159836 333374 207355 333376
rect 159836 333372 159842 333374
rect 207289 333371 207355 333374
rect 137461 333298 137527 333301
rect 146201 333298 146267 333301
rect 212533 333298 212599 333301
rect 137461 333296 212599 333298
rect 137461 333240 137466 333296
rect 137522 333240 146206 333296
rect 146262 333240 212538 333296
rect 212594 333240 212599 333296
rect 137461 333238 212599 333240
rect 137461 333235 137527 333238
rect 146201 333235 146267 333238
rect 212533 333235 212599 333238
rect 230381 333298 230447 333301
rect 258574 333298 258580 333300
rect 230381 333296 258580 333298
rect 230381 333240 230386 333296
rect 230442 333240 258580 333296
rect 230381 333238 258580 333240
rect 230381 333235 230447 333238
rect 258574 333236 258580 333238
rect 258644 333236 258650 333300
rect 124857 332618 124923 332621
rect 229277 332618 229343 332621
rect 230381 332618 230447 332621
rect 124857 332616 230447 332618
rect 124857 332560 124862 332616
rect 124918 332560 229282 332616
rect 229338 332560 230386 332616
rect 230442 332560 230447 332616
rect 124857 332558 230447 332560
rect 124857 332555 124923 332558
rect 229277 332555 229343 332558
rect 230381 332555 230447 332558
rect -960 332196 480 332436
rect 20713 331802 20779 331805
rect 158437 331802 158503 331805
rect 201493 331802 201559 331805
rect 274909 331802 274975 331805
rect 20713 331800 201559 331802
rect 20713 331744 20718 331800
rect 20774 331744 158442 331800
rect 158498 331744 201498 331800
rect 201554 331744 201559 331800
rect 20713 331742 201559 331744
rect 20713 331739 20779 331742
rect 158437 331739 158503 331742
rect 201493 331739 201559 331742
rect 209730 331800 274975 331802
rect 209730 331744 274914 331800
rect 274970 331744 274975 331800
rect 209730 331742 274975 331744
rect 133137 331258 133203 331261
rect 208393 331258 208459 331261
rect 209730 331258 209790 331742
rect 274909 331739 274975 331742
rect 133137 331256 209790 331258
rect 133137 331200 133142 331256
rect 133198 331200 208398 331256
rect 208454 331200 209790 331256
rect 133137 331198 209790 331200
rect 133137 331195 133203 331198
rect 208393 331195 208459 331198
rect 140681 331122 140747 331125
rect 144085 331122 144151 331125
rect 140681 331120 144151 331122
rect 140681 331064 140686 331120
rect 140742 331064 144090 331120
rect 144146 331064 144151 331120
rect 140681 331062 144151 331064
rect 140681 331059 140747 331062
rect 144085 331059 144151 331062
rect 251909 330714 251975 330717
rect 263910 330714 263916 330716
rect 251909 330712 263916 330714
rect 251909 330656 251914 330712
rect 251970 330656 263916 330712
rect 251909 330654 263916 330656
rect 251909 330651 251975 330654
rect 263910 330652 263916 330654
rect 263980 330652 263986 330716
rect 154481 330578 154547 330581
rect 166257 330580 166323 330581
rect 166206 330578 166212 330580
rect 154481 330576 166212 330578
rect 166276 330576 166323 330580
rect 154481 330520 154486 330576
rect 154542 330520 166212 330576
rect 166318 330520 166323 330576
rect 154481 330518 166212 330520
rect 154481 330515 154547 330518
rect 166206 330516 166212 330518
rect 166276 330516 166323 330520
rect 166257 330515 166323 330516
rect 238109 330578 238175 330581
rect 252502 330578 252508 330580
rect 238109 330576 252508 330578
rect 238109 330520 238114 330576
rect 238170 330520 252508 330576
rect 238109 330518 252508 330520
rect 238109 330515 238175 330518
rect 252502 330516 252508 330518
rect 252572 330516 252578 330580
rect 16573 330442 16639 330445
rect 172094 330442 172100 330444
rect 16573 330440 172100 330442
rect 16573 330384 16578 330440
rect 16634 330384 172100 330440
rect 16573 330382 172100 330384
rect 16573 330379 16639 330382
rect 172094 330380 172100 330382
rect 172164 330442 172170 330444
rect 172237 330442 172303 330445
rect 172164 330440 172303 330442
rect 172164 330384 172242 330440
rect 172298 330384 172303 330440
rect 172164 330382 172303 330384
rect 172164 330380 172170 330382
rect 172237 330379 172303 330382
rect 191557 330442 191623 330445
rect 263542 330442 263548 330444
rect 191557 330440 263548 330442
rect 191557 330384 191562 330440
rect 191618 330384 263548 330440
rect 191557 330382 263548 330384
rect 191557 330379 191623 330382
rect 263542 330380 263548 330382
rect 263612 330380 263618 330444
rect 143533 329898 143599 329901
rect 144085 329898 144151 329901
rect 207105 329898 207171 329901
rect 143533 329896 207171 329898
rect 143533 329840 143538 329896
rect 143594 329840 144090 329896
rect 144146 329840 207110 329896
rect 207166 329840 207171 329896
rect 143533 329838 207171 329840
rect 143533 329835 143599 329838
rect 144085 329835 144151 329838
rect 207105 329835 207171 329838
rect 216673 329762 216739 329765
rect 217409 329762 217475 329765
rect 216673 329760 217475 329762
rect 216673 329704 216678 329760
rect 216734 329704 217414 329760
rect 217470 329704 217475 329760
rect 216673 329702 217475 329704
rect 216673 329699 216739 329702
rect 217409 329699 217475 329702
rect 201677 329218 201743 329221
rect 219525 329218 219591 329221
rect 201677 329216 219591 329218
rect 201677 329160 201682 329216
rect 201738 329160 219530 329216
rect 219586 329160 219591 329216
rect 201677 329158 219591 329160
rect 201677 329155 201743 329158
rect 219525 329155 219591 329158
rect 253289 329218 253355 329221
rect 260966 329218 260972 329220
rect 253289 329216 260972 329218
rect 253289 329160 253294 329216
rect 253350 329160 260972 329216
rect 253289 329158 260972 329160
rect 253289 329155 253355 329158
rect 260966 329156 260972 329158
rect 261036 329156 261042 329220
rect 219341 329082 219407 329085
rect 299473 329082 299539 329085
rect 219341 329080 299539 329082
rect 219341 329024 219346 329080
rect 219402 329024 299478 329080
rect 299534 329024 299539 329080
rect 219341 329022 299539 329024
rect 219341 329019 219407 329022
rect 299473 329019 299539 329022
rect 131849 328674 131915 328677
rect 216673 328674 216739 328677
rect 131849 328672 216739 328674
rect 131849 328616 131854 328672
rect 131910 328616 216678 328672
rect 216734 328616 216739 328672
rect 131849 328614 216739 328616
rect 131849 328611 131915 328614
rect 216673 328611 216739 328614
rect 34513 328538 34579 328541
rect 222285 328538 222351 328541
rect 34513 328536 222351 328538
rect 34513 328480 34518 328536
rect 34574 328480 222290 328536
rect 222346 328480 222351 328536
rect 34513 328478 222351 328480
rect 34513 328475 34579 328478
rect 222285 328475 222351 328478
rect 205633 328402 205699 328405
rect 206369 328402 206435 328405
rect 205633 328400 206435 328402
rect 205633 328344 205638 328400
rect 205694 328344 206374 328400
rect 206430 328344 206435 328400
rect 205633 328342 206435 328344
rect 205633 328339 205699 328342
rect 206369 328339 206435 328342
rect 135897 327450 135963 327453
rect 205633 327450 205699 327453
rect 135897 327448 205699 327450
rect 135897 327392 135902 327448
rect 135958 327392 205638 327448
rect 205694 327392 205699 327448
rect 135897 327390 205699 327392
rect 135897 327387 135963 327390
rect 205633 327387 205699 327390
rect 162117 327314 162183 327317
rect 259494 327314 259500 327316
rect 162117 327312 259500 327314
rect 162117 327256 162122 327312
rect 162178 327256 259500 327312
rect 162117 327254 259500 327256
rect 162117 327251 162183 327254
rect 259494 327252 259500 327254
rect 259564 327252 259570 327316
rect 22093 327178 22159 327181
rect 220997 327178 221063 327181
rect 222101 327178 222167 327181
rect 22093 327176 222167 327178
rect 22093 327120 22098 327176
rect 22154 327120 221002 327176
rect 221058 327120 222106 327176
rect 222162 327120 222167 327176
rect 22093 327118 222167 327120
rect 22093 327115 22159 327118
rect 220997 327115 221063 327118
rect 222101 327115 222167 327118
rect 223573 327042 223639 327045
rect 224217 327042 224283 327045
rect 223573 327040 224283 327042
rect 223573 326984 223578 327040
rect 223634 326984 224222 327040
rect 224278 326984 224283 327040
rect 223573 326982 224283 326984
rect 223573 326979 223639 326982
rect 224217 326979 224283 326982
rect 153285 326362 153351 326365
rect 161289 326362 161355 326365
rect 204253 326362 204319 326365
rect 153285 326360 204319 326362
rect 153285 326304 153290 326360
rect 153346 326304 161294 326360
rect 161350 326304 204258 326360
rect 204314 326304 204319 326360
rect 153285 326302 204319 326304
rect 153285 326299 153351 326302
rect 161289 326299 161355 326302
rect 204253 326299 204319 326302
rect 41413 325818 41479 325821
rect 223573 325818 223639 325821
rect 41413 325816 223639 325818
rect 41413 325760 41418 325816
rect 41474 325760 223578 325816
rect 223634 325760 223639 325816
rect 41413 325758 223639 325760
rect 41413 325755 41479 325758
rect 223573 325755 223639 325758
rect 247125 325818 247191 325821
rect 265750 325818 265756 325820
rect 247125 325816 265756 325818
rect 247125 325760 247130 325816
rect 247186 325760 265756 325816
rect 247125 325758 265756 325760
rect 247125 325755 247191 325758
rect 265750 325756 265756 325758
rect 265820 325818 265826 325820
rect 265820 325758 579630 325818
rect 265820 325756 265826 325758
rect 579570 325682 579630 325758
rect 579570 325622 583586 325682
rect 583526 325410 583586 325622
rect 583342 325364 583586 325410
rect 583342 325350 584960 325364
rect 583342 325274 583402 325350
rect 583520 325274 584960 325350
rect 583342 325214 584960 325274
rect 155166 325076 155172 325140
rect 155236 325138 155242 325140
rect 234521 325138 234587 325141
rect 155236 325136 234587 325138
rect 155236 325080 234526 325136
rect 234582 325080 234587 325136
rect 583520 325124 584960 325214
rect 155236 325078 234587 325080
rect 155236 325076 155242 325078
rect 234521 325075 234587 325078
rect 67357 325002 67423 325005
rect 135989 325002 136055 325005
rect 258574 325002 258580 325004
rect 67357 325000 258580 325002
rect 67357 324944 67362 325000
rect 67418 324944 135994 325000
rect 136050 324944 258580 325000
rect 67357 324942 258580 324944
rect 67357 324939 67423 324942
rect 135989 324939 136055 324942
rect 258574 324940 258580 324942
rect 258644 324940 258650 325004
rect 123477 323778 123543 323781
rect 162117 323778 162183 323781
rect 123477 323776 162183 323778
rect 123477 323720 123482 323776
rect 123538 323720 162122 323776
rect 162178 323720 162183 323776
rect 123477 323718 162183 323720
rect 123477 323715 123543 323718
rect 162117 323715 162183 323718
rect 26233 323642 26299 323645
rect 162710 323642 162716 323644
rect 26233 323640 162716 323642
rect 26233 323584 26238 323640
rect 26294 323584 162716 323640
rect 26233 323582 162716 323584
rect 26233 323579 26299 323582
rect 162710 323580 162716 323582
rect 162780 323642 162786 323644
rect 202045 323642 202111 323645
rect 162780 323640 202111 323642
rect 162780 323584 202050 323640
rect 202106 323584 202111 323640
rect 162780 323582 202111 323584
rect 162780 323580 162786 323582
rect 202045 323579 202111 323582
rect 209037 323642 209103 323645
rect 267917 323642 267983 323645
rect 209037 323640 267983 323642
rect 209037 323584 209042 323640
rect 209098 323584 267922 323640
rect 267978 323584 267983 323640
rect 209037 323582 267983 323584
rect 209037 323579 209103 323582
rect 267917 323579 267983 323582
rect 173709 322962 173775 322965
rect 177297 322962 177363 322965
rect 173709 322960 177363 322962
rect 173709 322904 173714 322960
rect 173770 322904 177302 322960
rect 177358 322904 177363 322960
rect 173709 322902 177363 322904
rect 173709 322899 173775 322902
rect 177297 322899 177363 322902
rect 191649 322146 191715 322149
rect 267733 322146 267799 322149
rect 191649 322144 267799 322146
rect 191649 322088 191654 322144
rect 191710 322088 267738 322144
rect 267794 322088 267799 322144
rect 191649 322086 267799 322088
rect 191649 322083 191715 322086
rect 267733 322083 267799 322086
rect 152733 321602 152799 321605
rect 208485 321602 208551 321605
rect 209129 321602 209195 321605
rect 152733 321600 209195 321602
rect 152733 321544 152738 321600
rect 152794 321544 208490 321600
rect 208546 321544 209134 321600
rect 209190 321544 209195 321600
rect 152733 321542 209195 321544
rect 152733 321539 152799 321542
rect 208485 321539 208551 321542
rect 209129 321539 209195 321542
rect 181989 320922 182055 320925
rect 193305 320922 193371 320925
rect 181989 320920 193371 320922
rect 181989 320864 181994 320920
rect 182050 320864 193310 320920
rect 193366 320864 193371 320920
rect 181989 320862 193371 320864
rect 181989 320859 182055 320862
rect 193305 320859 193371 320862
rect 15193 320786 15259 320789
rect 155718 320786 155724 320788
rect 15193 320784 155724 320786
rect 15193 320728 15198 320784
rect 15254 320728 155724 320784
rect 15193 320726 155724 320728
rect 15193 320723 15259 320726
rect 155718 320724 155724 320726
rect 155788 320786 155794 320788
rect 197353 320786 197419 320789
rect 155788 320784 197419 320786
rect 155788 320728 197358 320784
rect 197414 320728 197419 320784
rect 155788 320726 197419 320728
rect 155788 320724 155794 320726
rect 197353 320723 197419 320726
rect 97758 320180 97764 320244
rect 97828 320242 97834 320244
rect 284477 320242 284543 320245
rect 97828 320240 284543 320242
rect 97828 320184 284482 320240
rect 284538 320184 284543 320240
rect 97828 320182 284543 320184
rect 97828 320180 97834 320182
rect 284477 320179 284543 320182
rect 154113 319426 154179 319429
rect 170806 319426 170812 319428
rect 154113 319424 170812 319426
rect -960 319290 480 319380
rect 154113 319368 154118 319424
rect 154174 319368 170812 319424
rect 154113 319366 170812 319368
rect 154113 319363 154179 319366
rect 170806 319364 170812 319366
rect 170876 319426 170882 319428
rect 204713 319426 204779 319429
rect 170876 319424 204779 319426
rect 170876 319368 204718 319424
rect 204774 319368 204779 319424
rect 170876 319366 204779 319368
rect 170876 319364 170882 319366
rect 204713 319363 204779 319366
rect 204897 319426 204963 319429
rect 254025 319426 254091 319429
rect 204897 319424 254091 319426
rect 204897 319368 204902 319424
rect 204958 319368 254030 319424
rect 254086 319368 254091 319424
rect 204897 319366 254091 319368
rect 204897 319363 204963 319366
rect 254025 319363 254091 319366
rect 260189 319426 260255 319429
rect 269062 319426 269068 319428
rect 260189 319424 269068 319426
rect 260189 319368 260194 319424
rect 260250 319368 269068 319424
rect 260189 319366 269068 319368
rect 260189 319363 260255 319366
rect 269062 319364 269068 319366
rect 269132 319364 269138 319428
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 169518 318820 169524 318884
rect 169588 318882 169594 318884
rect 203057 318882 203123 318885
rect 169588 318880 203123 318882
rect 169588 318824 203062 318880
rect 203118 318824 203123 318880
rect 169588 318822 203123 318824
rect 169588 318820 169594 318822
rect 203057 318819 203123 318822
rect 214005 318746 214071 318749
rect 214557 318746 214623 318749
rect 214005 318744 214623 318746
rect 214005 318688 214010 318744
rect 214066 318688 214562 318744
rect 214618 318688 214623 318744
rect 214005 318686 214623 318688
rect 214005 318683 214071 318686
rect 214557 318683 214623 318686
rect 152549 318202 152615 318205
rect 152917 318202 152983 318205
rect 208577 318202 208643 318205
rect 152549 318200 208643 318202
rect 152549 318144 152554 318200
rect 152610 318144 152922 318200
rect 152978 318144 208582 318200
rect 208638 318144 208643 318200
rect 152549 318142 208643 318144
rect 152549 318139 152615 318142
rect 152917 318139 152983 318142
rect 208577 318139 208643 318142
rect 109534 318004 109540 318068
rect 109604 318066 109610 318068
rect 167637 318066 167703 318069
rect 109604 318064 167703 318066
rect 109604 318008 167642 318064
rect 167698 318008 167703 318064
rect 109604 318006 167703 318008
rect 109604 318004 109610 318006
rect 167637 318003 167703 318006
rect 233969 318066 234035 318069
rect 264973 318066 265039 318069
rect 233969 318064 265039 318066
rect 233969 318008 233974 318064
rect 234030 318008 264978 318064
rect 265034 318008 265039 318064
rect 233969 318006 265039 318008
rect 233969 318003 234035 318006
rect 264973 318003 265039 318006
rect 79726 317460 79732 317524
rect 79796 317522 79802 317524
rect 106917 317522 106983 317525
rect 79796 317520 106983 317522
rect 79796 317464 106922 317520
rect 106978 317464 106983 317520
rect 79796 317462 106983 317464
rect 79796 317460 79802 317462
rect 106917 317459 106983 317462
rect 147121 317522 147187 317525
rect 152549 317522 152615 317525
rect 147121 317520 152615 317522
rect 147121 317464 147126 317520
rect 147182 317464 152554 317520
rect 152610 317464 152615 317520
rect 147121 317462 152615 317464
rect 147121 317459 147187 317462
rect 152549 317459 152615 317462
rect 162117 317522 162183 317525
rect 214005 317522 214071 317525
rect 162117 317520 214071 317522
rect 162117 317464 162122 317520
rect 162178 317464 214010 317520
rect 214066 317464 214071 317520
rect 162117 317462 214071 317464
rect 162117 317459 162183 317462
rect 214005 317459 214071 317462
rect 254577 317386 254643 317389
rect 256734 317386 256740 317388
rect 254577 317384 256740 317386
rect 254577 317328 254582 317384
rect 254638 317328 256740 317384
rect 254577 317326 256740 317328
rect 254577 317323 254643 317326
rect 256734 317324 256740 317326
rect 256804 317324 256810 317388
rect 230565 316842 230631 316845
rect 161430 316840 230631 316842
rect 161430 316784 230570 316840
rect 230626 316784 230631 316840
rect 161430 316782 230631 316784
rect 89437 316706 89503 316709
rect 99465 316706 99531 316709
rect 89437 316704 99531 316706
rect 89437 316648 89442 316704
rect 89498 316648 99470 316704
rect 99526 316648 99531 316704
rect 89437 316646 99531 316648
rect 89437 316643 89503 316646
rect 99465 316643 99531 316646
rect 137277 316706 137343 316709
rect 159909 316706 159975 316709
rect 161430 316706 161490 316782
rect 230565 316779 230631 316782
rect 137277 316704 161490 316706
rect 137277 316648 137282 316704
rect 137338 316648 159914 316704
rect 159970 316648 161490 316704
rect 137277 316646 161490 316648
rect 195973 316706 196039 316709
rect 276238 316706 276244 316708
rect 195973 316704 276244 316706
rect 195973 316648 195978 316704
rect 196034 316648 276244 316704
rect 195973 316646 276244 316648
rect 137277 316643 137343 316646
rect 159909 316643 159975 316646
rect 195973 316643 196039 316646
rect 276238 316644 276244 316646
rect 276308 316644 276314 316708
rect 175181 316162 175247 316165
rect 195421 316162 195487 316165
rect 175181 316160 195487 316162
rect 175181 316104 175186 316160
rect 175242 316104 195426 316160
rect 195482 316104 195487 316160
rect 175181 316102 195487 316104
rect 175181 316099 175247 316102
rect 195421 316099 195487 316102
rect 86718 315964 86724 316028
rect 86788 316026 86794 316028
rect 148869 316026 148935 316029
rect 86788 316024 148935 316026
rect 86788 315968 148874 316024
rect 148930 315968 148935 316024
rect 86788 315966 148935 315968
rect 86788 315964 86794 315966
rect 148869 315963 148935 315966
rect 93761 315346 93827 315349
rect 105118 315346 105124 315348
rect 93761 315344 105124 315346
rect 93761 315288 93766 315344
rect 93822 315288 105124 315344
rect 93761 315286 105124 315288
rect 93761 315283 93827 315286
rect 105118 315284 105124 315286
rect 105188 315284 105194 315348
rect 195329 315346 195395 315349
rect 204989 315346 205055 315349
rect 195329 315344 205055 315346
rect 195329 315288 195334 315344
rect 195390 315288 204994 315344
rect 205050 315288 205055 315344
rect 195329 315286 205055 315288
rect 195329 315283 195395 315286
rect 204989 315283 205055 315286
rect 220077 315346 220143 315349
rect 254117 315346 254183 315349
rect 220077 315344 254183 315346
rect 220077 315288 220082 315344
rect 220138 315288 254122 315344
rect 254178 315288 254183 315344
rect 220077 315286 254183 315288
rect 220077 315283 220143 315286
rect 254117 315283 254183 315286
rect 155217 314802 155283 314805
rect 213085 314802 213151 314805
rect 155217 314800 213151 314802
rect 155217 314744 155222 314800
rect 155278 314744 213090 314800
rect 213146 314744 213151 314800
rect 155217 314742 213151 314744
rect 155217 314739 155283 314742
rect 213085 314739 213151 314742
rect 237281 314122 237347 314125
rect 269113 314122 269179 314125
rect 237281 314120 269179 314122
rect 237281 314064 237286 314120
rect 237342 314064 269118 314120
rect 269174 314064 269179 314120
rect 237281 314062 269179 314064
rect 237281 314059 237347 314062
rect 269113 314059 269179 314062
rect 86769 313986 86835 313989
rect 95182 313986 95188 313988
rect 86769 313984 95188 313986
rect 86769 313928 86774 313984
rect 86830 313928 95188 313984
rect 86769 313926 95188 313928
rect 86769 313923 86835 313926
rect 95182 313924 95188 313926
rect 95252 313924 95258 313988
rect 208577 313986 208643 313989
rect 235993 313986 236059 313989
rect 208577 313984 236059 313986
rect 208577 313928 208582 313984
rect 208638 313928 235998 313984
rect 236054 313928 236059 313984
rect 208577 313926 236059 313928
rect 208577 313923 208643 313926
rect 235993 313923 236059 313926
rect 238661 313986 238727 313989
rect 270534 313986 270540 313988
rect 238661 313984 270540 313986
rect 238661 313928 238666 313984
rect 238722 313928 270540 313984
rect 238661 313926 270540 313928
rect 238661 313923 238727 313926
rect 270534 313924 270540 313926
rect 270604 313924 270610 313988
rect 166758 313380 166764 313444
rect 166828 313442 166834 313444
rect 213177 313442 213243 313445
rect 166828 313440 213243 313442
rect 166828 313384 213182 313440
rect 213238 313384 213243 313440
rect 166828 313382 213243 313384
rect 166828 313380 166834 313382
rect 213177 313379 213243 313382
rect 148685 313306 148751 313309
rect 200205 313306 200271 313309
rect 200757 313306 200823 313309
rect 148685 313304 200823 313306
rect 148685 313248 148690 313304
rect 148746 313248 200210 313304
rect 200266 313248 200762 313304
rect 200818 313248 200823 313304
rect 148685 313246 200823 313248
rect 148685 313243 148751 313246
rect 200205 313243 200271 313246
rect 200757 313243 200823 313246
rect 84101 312490 84167 312493
rect 92790 312490 92796 312492
rect 84101 312488 92796 312490
rect 84101 312432 84106 312488
rect 84162 312432 92796 312488
rect 84101 312430 92796 312432
rect 84101 312427 84167 312430
rect 92790 312428 92796 312430
rect 92860 312428 92866 312492
rect 95325 312490 95391 312493
rect 109534 312490 109540 312492
rect 95325 312488 109540 312490
rect 95325 312432 95330 312488
rect 95386 312432 109540 312488
rect 95325 312430 109540 312432
rect 95325 312427 95391 312430
rect 109534 312428 109540 312430
rect 109604 312428 109610 312492
rect 159357 312082 159423 312085
rect 160686 312082 160692 312084
rect 159357 312080 160692 312082
rect 159357 312024 159362 312080
rect 159418 312024 160692 312080
rect 159357 312022 160692 312024
rect 159357 312019 159423 312022
rect 160686 312020 160692 312022
rect 160756 312020 160762 312084
rect 176653 312082 176719 312085
rect 177665 312082 177731 312085
rect 211337 312082 211403 312085
rect 176653 312080 211403 312082
rect 176653 312024 176658 312080
rect 176714 312024 177670 312080
rect 177726 312024 211342 312080
rect 211398 312024 211403 312080
rect 176653 312022 211403 312024
rect 176653 312019 176719 312022
rect 177665 312019 177731 312022
rect 211337 312019 211403 312022
rect 233141 312082 233207 312085
rect 266302 312082 266308 312084
rect 233141 312080 266308 312082
rect 233141 312024 233146 312080
rect 233202 312024 266308 312080
rect 233141 312022 266308 312024
rect 233141 312019 233207 312022
rect 266302 312020 266308 312022
rect 266372 312020 266378 312084
rect 582649 312082 582715 312085
rect 583520 312082 584960 312172
rect 582649 312080 584960 312082
rect 582649 312024 582654 312080
rect 582710 312024 584960 312080
rect 582649 312022 584960 312024
rect 582649 312019 582715 312022
rect 140037 311946 140103 311949
rect 228265 311946 228331 311949
rect 140037 311944 228331 311946
rect 140037 311888 140042 311944
rect 140098 311888 228270 311944
rect 228326 311888 228331 311944
rect 140037 311886 228331 311888
rect 140037 311883 140103 311886
rect 228265 311883 228331 311886
rect 244825 311946 244891 311949
rect 245009 311946 245075 311949
rect 291193 311946 291259 311949
rect 244825 311944 291259 311946
rect 244825 311888 244830 311944
rect 244886 311888 245014 311944
rect 245070 311888 291198 311944
rect 291254 311888 291259 311944
rect 583520 311932 584960 312022
rect 244825 311886 291259 311888
rect 244825 311883 244891 311886
rect 245009 311883 245075 311886
rect 291193 311883 291259 311886
rect 169109 311402 169175 311405
rect 176653 311402 176719 311405
rect 169109 311400 176719 311402
rect 169109 311344 169114 311400
rect 169170 311344 176658 311400
rect 176714 311344 176719 311400
rect 169109 311342 176719 311344
rect 169109 311339 169175 311342
rect 176653 311339 176719 311342
rect 260281 311402 260347 311405
rect 266486 311402 266492 311404
rect 260281 311400 266492 311402
rect 260281 311344 260286 311400
rect 260342 311344 266492 311400
rect 260281 311342 266492 311344
rect 260281 311339 260347 311342
rect 266486 311340 266492 311342
rect 266556 311340 266562 311404
rect 173801 311266 173867 311269
rect 225873 311266 225939 311269
rect 161430 311264 225939 311266
rect 161430 311208 173806 311264
rect 173862 311208 225878 311264
rect 225934 311208 225939 311264
rect 161430 311206 225939 311208
rect 80789 311130 80855 311133
rect 90030 311130 90036 311132
rect 80789 311128 90036 311130
rect 80789 311072 80794 311128
rect 80850 311072 90036 311128
rect 80789 311070 90036 311072
rect 80789 311067 80855 311070
rect 90030 311068 90036 311070
rect 90100 311068 90106 311132
rect 91001 311130 91067 311133
rect 98494 311130 98500 311132
rect 91001 311128 98500 311130
rect 91001 311072 91006 311128
rect 91062 311072 98500 311128
rect 91001 311070 98500 311072
rect 91001 311067 91067 311070
rect 98494 311068 98500 311070
rect 98564 311068 98570 311132
rect 145557 311130 145623 311133
rect 161430 311130 161490 311206
rect 173801 311203 173867 311206
rect 225873 311203 225939 311206
rect 249609 311266 249675 311269
rect 252461 311266 252527 311269
rect 269757 311266 269823 311269
rect 249609 311264 269823 311266
rect 249609 311208 249614 311264
rect 249670 311208 252466 311264
rect 252522 311208 269762 311264
rect 269818 311208 269823 311264
rect 249609 311206 269823 311208
rect 249609 311203 249675 311206
rect 252461 311203 252527 311206
rect 269757 311203 269823 311206
rect 211245 311130 211311 311133
rect 282913 311130 282979 311133
rect 145557 311128 161490 311130
rect 145557 311072 145562 311128
rect 145618 311072 161490 311128
rect 145557 311070 161490 311072
rect 200070 311128 282979 311130
rect 200070 311072 211250 311128
rect 211306 311072 282918 311128
rect 282974 311072 282979 311128
rect 200070 311070 282979 311072
rect 145557 311067 145623 311070
rect 177481 310586 177547 310589
rect 200070 310586 200130 311070
rect 211245 311067 211311 311070
rect 282913 311067 282979 311070
rect 177481 310584 200130 310586
rect 177481 310528 177486 310584
rect 177542 310528 200130 310584
rect 177481 310526 200130 310528
rect 177481 310523 177547 310526
rect 57697 310450 57763 310453
rect 144729 310450 144795 310453
rect 57697 310448 144795 310450
rect 57697 310392 57702 310448
rect 57758 310392 144734 310448
rect 144790 310392 144795 310448
rect 57697 310390 144795 310392
rect 57697 310387 57763 310390
rect 144729 310387 144795 310390
rect 94497 309770 94563 309773
rect 106406 309770 106412 309772
rect 94497 309768 106412 309770
rect 94497 309712 94502 309768
rect 94558 309712 106412 309768
rect 94497 309710 106412 309712
rect 94497 309707 94563 309710
rect 106406 309708 106412 309710
rect 106476 309708 106482 309772
rect 144729 309770 144795 309773
rect 176653 309770 176719 309773
rect 144729 309768 176719 309770
rect 144729 309712 144734 309768
rect 144790 309712 176658 309768
rect 176714 309712 176719 309768
rect 144729 309710 176719 309712
rect 144729 309707 144795 309710
rect 176653 309707 176719 309710
rect 185669 309498 185735 309501
rect 226425 309498 226491 309501
rect 185669 309496 226491 309498
rect 185669 309440 185674 309496
rect 185730 309440 226430 309496
rect 226486 309440 226491 309496
rect 185669 309438 226491 309440
rect 185669 309435 185735 309438
rect 226425 309435 226491 309438
rect 146937 309362 147003 309365
rect 195973 309362 196039 309365
rect 146937 309360 196039 309362
rect 146937 309304 146942 309360
rect 146998 309304 195978 309360
rect 196034 309304 196039 309360
rect 146937 309302 196039 309304
rect 146937 309299 147003 309302
rect 195973 309299 196039 309302
rect 251817 309362 251883 309365
rect 295517 309362 295583 309365
rect 251817 309360 295583 309362
rect 251817 309304 251822 309360
rect 251878 309304 295522 309360
rect 295578 309304 295583 309360
rect 251817 309302 295583 309304
rect 251817 309299 251883 309302
rect 295517 309299 295583 309302
rect 187693 309226 187759 309229
rect 278773 309226 278839 309229
rect 278957 309226 279023 309229
rect 187693 309224 279023 309226
rect 187693 309168 187698 309224
rect 187754 309168 278778 309224
rect 278834 309168 278962 309224
rect 279018 309168 279023 309224
rect 187693 309166 279023 309168
rect 187693 309163 187759 309166
rect 278773 309163 278839 309166
rect 278957 309163 279023 309166
rect 76649 309090 76715 309093
rect 83038 309090 83044 309092
rect 76649 309088 83044 309090
rect 76649 309032 76654 309088
rect 76710 309032 83044 309088
rect 76649 309030 83044 309032
rect 76649 309027 76715 309030
rect 83038 309028 83044 309030
rect 83108 309028 83114 309092
rect 233417 309090 233483 309093
rect 233969 309090 234035 309093
rect 233417 309088 234035 309090
rect 233417 309032 233422 309088
rect 233478 309032 233974 309088
rect 234030 309032 234035 309088
rect 233417 309030 234035 309032
rect 233417 309027 233483 309030
rect 233969 309027 234035 309030
rect 276013 309090 276079 309093
rect 276289 309090 276355 309093
rect 276013 309088 276355 309090
rect 276013 309032 276018 309088
rect 276074 309032 276294 309088
rect 276350 309032 276355 309088
rect 276013 309030 276355 309032
rect 276013 309027 276079 309030
rect 276289 309027 276355 309030
rect 84009 308410 84075 308413
rect 92606 308410 92612 308412
rect 84009 308408 92612 308410
rect 84009 308352 84014 308408
rect 84070 308352 92612 308408
rect 84009 308350 92612 308352
rect 84009 308347 84075 308350
rect 92606 308348 92612 308350
rect 92676 308348 92682 308412
rect 194726 308076 194732 308140
rect 194796 308138 194802 308140
rect 229737 308138 229803 308141
rect 194796 308136 229803 308138
rect 194796 308080 229742 308136
rect 229798 308080 229803 308136
rect 194796 308078 229803 308080
rect 194796 308076 194802 308078
rect 229737 308075 229803 308078
rect 187049 308002 187115 308005
rect 233417 308002 233483 308005
rect 187049 308000 233483 308002
rect 187049 307944 187054 308000
rect 187110 307944 233422 308000
rect 233478 307944 233483 308000
rect 187049 307942 233483 307944
rect 187049 307939 187115 307942
rect 233417 307939 233483 307942
rect 247677 308002 247743 308005
rect 291285 308002 291351 308005
rect 247677 308000 291351 308002
rect 247677 307944 247682 308000
rect 247738 307944 291290 308000
rect 291346 307944 291351 308000
rect 247677 307942 291351 307944
rect 247677 307939 247743 307942
rect 291285 307939 291351 307942
rect 70301 307866 70367 307869
rect 76046 307866 76052 307868
rect 70301 307864 76052 307866
rect 70301 307808 70306 307864
rect 70362 307808 76052 307864
rect 70301 307806 76052 307808
rect 70301 307803 70367 307806
rect 76046 307804 76052 307806
rect 76116 307804 76122 307868
rect 120717 307866 120783 307869
rect 276013 307866 276079 307869
rect 120717 307864 276079 307866
rect 120717 307808 120722 307864
rect 120778 307808 276018 307864
rect 276074 307808 276079 307864
rect 120717 307806 276079 307808
rect 120717 307803 120783 307806
rect 276013 307803 276079 307806
rect 84510 307668 84516 307732
rect 84580 307730 84586 307732
rect 86953 307730 87019 307733
rect 84580 307728 87019 307730
rect 84580 307672 86958 307728
rect 87014 307672 87019 307728
rect 84580 307670 87019 307672
rect 84580 307668 84586 307670
rect 86953 307667 87019 307670
rect 246389 307186 246455 307189
rect 259678 307186 259684 307188
rect 246389 307184 259684 307186
rect 246389 307128 246394 307184
rect 246450 307128 259684 307184
rect 246389 307126 259684 307128
rect 246389 307123 246455 307126
rect 259678 307124 259684 307126
rect 259748 307124 259754 307188
rect 88241 307050 88307 307053
rect 97942 307050 97948 307052
rect 88241 307048 97948 307050
rect 88241 306992 88246 307048
rect 88302 306992 97948 307048
rect 88241 306990 97948 306992
rect 88241 306987 88307 306990
rect 97942 306988 97948 306990
rect 98012 306988 98018 307052
rect 122097 307050 122163 307053
rect 142061 307050 142127 307053
rect 156597 307050 156663 307053
rect 122097 307048 156663 307050
rect 122097 306992 122102 307048
rect 122158 306992 142066 307048
rect 142122 306992 156602 307048
rect 156658 306992 156663 307048
rect 122097 306990 156663 306992
rect 122097 306987 122163 306990
rect 142061 306987 142127 306990
rect 156597 306987 156663 306990
rect 251909 307050 251975 307053
rect 267733 307050 267799 307053
rect 251909 307048 267799 307050
rect 251909 306992 251914 307048
rect 251970 306992 267738 307048
rect 267794 306992 267799 307048
rect 251909 306990 267799 306992
rect 251909 306987 251975 306990
rect 267733 306987 267799 306990
rect 160185 306914 160251 306917
rect 252277 306914 252343 306917
rect 160185 306912 252343 306914
rect 160185 306856 160190 306912
rect 160246 306856 252282 306912
rect 252338 306856 252343 306912
rect 160185 306854 252343 306856
rect 160185 306851 160251 306854
rect 252277 306851 252343 306854
rect 176101 306778 176167 306781
rect 213821 306778 213887 306781
rect 176101 306776 213887 306778
rect 176101 306720 176106 306776
rect 176162 306720 213826 306776
rect 213882 306720 213887 306776
rect 176101 306718 213887 306720
rect 176101 306715 176167 306718
rect 213821 306715 213887 306718
rect 182817 306642 182883 306645
rect 226885 306642 226951 306645
rect 182817 306640 226951 306642
rect 182817 306584 182822 306640
rect 182878 306584 226890 306640
rect 226946 306584 226951 306640
rect 182817 306582 226951 306584
rect 182817 306579 182883 306582
rect 226885 306579 226951 306582
rect 77293 306506 77359 306509
rect 86718 306506 86724 306508
rect 77293 306504 86724 306506
rect 77293 306448 77298 306504
rect 77354 306448 86724 306504
rect 77293 306446 86724 306448
rect 77293 306443 77359 306446
rect 86718 306444 86724 306446
rect 86788 306444 86794 306508
rect 251357 306506 251423 306509
rect 296713 306506 296779 306509
rect 251357 306504 296779 306506
rect 251357 306448 251362 306504
rect 251418 306448 296718 306504
rect 296774 306448 296779 306504
rect 251357 306446 296779 306448
rect 251357 306443 251423 306446
rect 296713 306443 296779 306446
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 83457 305826 83523 305829
rect 91502 305826 91508 305828
rect 83457 305824 91508 305826
rect 83457 305768 83462 305824
rect 83518 305768 91508 305824
rect 83457 305766 91508 305768
rect 83457 305763 83523 305766
rect 91502 305764 91508 305766
rect 91572 305764 91578 305828
rect 240777 305826 240843 305829
rect 256969 305826 257035 305829
rect 240777 305824 257035 305826
rect 240777 305768 240782 305824
rect 240838 305768 256974 305824
rect 257030 305768 257035 305824
rect 240777 305766 257035 305768
rect 240777 305763 240843 305766
rect 256969 305763 257035 305766
rect 90357 305690 90423 305693
rect 188061 305690 188127 305693
rect 90357 305688 188127 305690
rect 90357 305632 90362 305688
rect 90418 305632 188066 305688
rect 188122 305632 188127 305688
rect 90357 305630 188127 305632
rect 90357 305627 90423 305630
rect 188061 305627 188127 305630
rect 198733 305690 198799 305693
rect 242157 305690 242223 305693
rect 198733 305688 242223 305690
rect 198733 305632 198738 305688
rect 198794 305632 242162 305688
rect 242218 305632 242223 305688
rect 198733 305630 242223 305632
rect 198733 305627 198799 305630
rect 242157 305627 242223 305630
rect 187785 305282 187851 305285
rect 217133 305282 217199 305285
rect 217317 305282 217383 305285
rect 187785 305280 217383 305282
rect 187785 305224 187790 305280
rect 187846 305224 217138 305280
rect 217194 305224 217322 305280
rect 217378 305224 217383 305280
rect 187785 305222 217383 305224
rect 187785 305219 187851 305222
rect 217133 305219 217199 305222
rect 217317 305219 217383 305222
rect 186405 305146 186471 305149
rect 205817 305146 205883 305149
rect 206277 305146 206343 305149
rect 186405 305144 206343 305146
rect 186405 305088 186410 305144
rect 186466 305088 205822 305144
rect 205878 305088 206282 305144
rect 206338 305088 206343 305144
rect 186405 305086 206343 305088
rect 186405 305083 186471 305086
rect 205817 305083 205883 305086
rect 206277 305083 206343 305086
rect 185342 304948 185348 305012
rect 185412 305010 185418 305012
rect 186814 305010 186820 305012
rect 185412 304950 186820 305010
rect 185412 304948 185418 304950
rect 186814 304948 186820 304950
rect 186884 305010 186890 305012
rect 187509 305010 187575 305013
rect 186884 305008 187575 305010
rect 186884 304952 187514 305008
rect 187570 304952 187575 305008
rect 186884 304950 187575 304952
rect 186884 304948 186890 304950
rect 187509 304947 187575 304950
rect 246941 305010 247007 305013
rect 302325 305010 302391 305013
rect 246941 305008 302391 305010
rect 246941 304952 246946 305008
rect 247002 304952 302330 305008
rect 302386 304952 302391 305008
rect 246941 304950 302391 304952
rect 246941 304947 247007 304950
rect 302325 304947 302391 304950
rect 159214 304268 159220 304332
rect 159284 304330 159290 304332
rect 198733 304330 198799 304333
rect 159284 304328 198799 304330
rect 159284 304272 198738 304328
rect 198794 304272 198799 304328
rect 159284 304270 198799 304272
rect 159284 304268 159290 304270
rect 198733 304267 198799 304270
rect 223849 304330 223915 304333
rect 238017 304330 238083 304333
rect 223849 304328 238083 304330
rect 223849 304272 223854 304328
rect 223910 304272 238022 304328
rect 238078 304272 238083 304328
rect 223849 304270 238083 304272
rect 223849 304267 223915 304270
rect 238017 304267 238083 304270
rect 82629 304194 82695 304197
rect 89662 304194 89668 304196
rect 82629 304192 89668 304194
rect 82629 304136 82634 304192
rect 82690 304136 89668 304192
rect 82629 304134 89668 304136
rect 82629 304131 82695 304134
rect 89662 304132 89668 304134
rect 89732 304132 89738 304196
rect 101254 304132 101260 304196
rect 101324 304194 101330 304196
rect 113265 304194 113331 304197
rect 101324 304192 113331 304194
rect 101324 304136 113270 304192
rect 113326 304136 113331 304192
rect 101324 304134 113331 304136
rect 101324 304132 101330 304134
rect 113265 304131 113331 304134
rect 182766 304132 182772 304196
rect 182836 304194 182842 304196
rect 227621 304194 227687 304197
rect 182836 304192 227687 304194
rect 182836 304136 227626 304192
rect 227682 304136 227687 304192
rect 182836 304134 227687 304136
rect 182836 304132 182842 304134
rect 227621 304131 227687 304134
rect 249057 304194 249123 304197
rect 262438 304194 262444 304196
rect 249057 304192 262444 304194
rect 249057 304136 249062 304192
rect 249118 304136 262444 304192
rect 249057 304134 262444 304136
rect 249057 304131 249123 304134
rect 262438 304132 262444 304134
rect 262508 304132 262514 304196
rect 273437 303922 273503 303925
rect 248370 303920 273503 303922
rect 248370 303864 273442 303920
rect 273498 303864 273503 303920
rect 248370 303862 273503 303864
rect 242985 303786 243051 303789
rect 243537 303786 243603 303789
rect 248370 303786 248430 303862
rect 273437 303859 273503 303862
rect 242985 303784 248430 303786
rect 242985 303728 242990 303784
rect 243046 303728 243542 303784
rect 243598 303728 248430 303784
rect 242985 303726 248430 303728
rect 242985 303723 243051 303726
rect 243537 303723 243603 303726
rect 249742 303724 249748 303788
rect 249812 303786 249818 303788
rect 250805 303786 250871 303789
rect 249812 303784 250871 303786
rect 249812 303728 250810 303784
rect 250866 303728 250871 303784
rect 249812 303726 250871 303728
rect 249812 303724 249818 303726
rect 250805 303723 250871 303726
rect 226977 303650 227043 303653
rect 227989 303650 228055 303653
rect 226977 303648 228055 303650
rect 226977 303592 226982 303648
rect 227038 303592 227994 303648
rect 228050 303592 228055 303648
rect 226977 303590 228055 303592
rect 226977 303587 227043 303590
rect 227989 303587 228055 303590
rect 244917 303650 244983 303653
rect 253197 303650 253263 303653
rect 244917 303648 253263 303650
rect 244917 303592 244922 303648
rect 244978 303592 253202 303648
rect 253258 303592 253263 303648
rect 244917 303590 253263 303592
rect 244917 303587 244983 303590
rect 253197 303587 253263 303590
rect 262254 303588 262260 303652
rect 262324 303650 262330 303652
rect 262489 303650 262555 303653
rect 262324 303648 262555 303650
rect 262324 303592 262494 303648
rect 262550 303592 262555 303648
rect 262324 303590 262555 303592
rect 262324 303588 262330 303590
rect 262489 303587 262555 303590
rect 151670 302772 151676 302836
rect 151740 302834 151746 302836
rect 166257 302834 166323 302837
rect 151740 302832 166323 302834
rect 151740 302776 166262 302832
rect 166318 302776 166323 302832
rect 151740 302774 166323 302776
rect 151740 302772 151746 302774
rect 166257 302771 166323 302774
rect 239121 302834 239187 302837
rect 582373 302834 582439 302837
rect 239121 302832 582439 302834
rect 239121 302776 239126 302832
rect 239182 302776 582378 302832
rect 582434 302776 582439 302832
rect 239121 302774 582439 302776
rect 239121 302771 239187 302774
rect 582373 302771 582439 302774
rect 175181 302562 175247 302565
rect 186221 302564 186287 302565
rect 178534 302562 178540 302564
rect 175181 302560 178540 302562
rect 175181 302504 175186 302560
rect 175242 302504 178540 302560
rect 175181 302502 178540 302504
rect 175181 302499 175247 302502
rect 178534 302500 178540 302502
rect 178604 302500 178610 302564
rect 186221 302562 186268 302564
rect 186140 302560 186268 302562
rect 186332 302562 186338 302564
rect 208209 302562 208275 302565
rect 186332 302560 208275 302562
rect 186140 302504 186226 302560
rect 186332 302504 208214 302560
rect 208270 302504 208275 302560
rect 186140 302502 186268 302504
rect 186221 302500 186268 302502
rect 186332 302502 208275 302504
rect 186332 302500 186338 302502
rect 186221 302499 186287 302500
rect 208209 302499 208275 302502
rect 166942 302364 166948 302428
rect 167012 302426 167018 302428
rect 168230 302426 168236 302428
rect 167012 302366 168236 302426
rect 167012 302364 167018 302366
rect 168230 302364 168236 302366
rect 168300 302426 168306 302428
rect 238201 302426 238267 302429
rect 168300 302424 238267 302426
rect 168300 302368 238206 302424
rect 238262 302368 238267 302424
rect 168300 302366 238267 302368
rect 168300 302364 168306 302366
rect 238201 302363 238267 302366
rect 248965 302426 249031 302429
rect 249701 302426 249767 302429
rect 259269 302426 259335 302429
rect 248965 302424 259335 302426
rect 248965 302368 248970 302424
rect 249026 302368 249706 302424
rect 249762 302368 259274 302424
rect 259330 302368 259335 302424
rect 248965 302366 259335 302368
rect 248965 302363 249031 302366
rect 249701 302363 249767 302366
rect 259269 302363 259335 302366
rect 17953 302290 18019 302293
rect 220813 302290 220879 302293
rect 17953 302288 220879 302290
rect 17953 302232 17958 302288
rect 18014 302232 220818 302288
rect 220874 302232 220879 302288
rect 17953 302230 220879 302232
rect 17953 302227 18019 302230
rect 220813 302227 220879 302230
rect 252277 302290 252343 302293
rect 254209 302290 254275 302293
rect 252277 302288 254275 302290
rect 252277 302232 252282 302288
rect 252338 302232 254214 302288
rect 254270 302232 254275 302288
rect 252277 302230 254275 302232
rect 252277 302227 252343 302230
rect 254209 302227 254275 302230
rect 258717 302290 258783 302293
rect 259453 302290 259519 302293
rect 258717 302288 259519 302290
rect 258717 302232 258722 302288
rect 258778 302232 259458 302288
rect 259514 302232 259519 302288
rect 258717 302230 259519 302232
rect 258717 302227 258783 302230
rect 259453 302227 259519 302230
rect 192937 301882 193003 301885
rect 195329 301882 195395 301885
rect 192937 301880 195395 301882
rect 192937 301824 192942 301880
rect 192998 301824 195334 301880
rect 195390 301824 195395 301880
rect 192937 301822 195395 301824
rect 192937 301819 193003 301822
rect 195329 301819 195395 301822
rect 193765 301746 193831 301749
rect 195053 301746 195119 301749
rect 193765 301744 195119 301746
rect 193765 301688 193770 301744
rect 193826 301688 195058 301744
rect 195114 301688 195119 301744
rect 193765 301686 195119 301688
rect 193765 301683 193831 301686
rect 195053 301683 195119 301686
rect 226885 301744 226951 301749
rect 226885 301688 226890 301744
rect 226946 301688 226951 301744
rect 226885 301683 226951 301688
rect 86534 301548 86540 301612
rect 86604 301610 86610 301612
rect 91093 301610 91159 301613
rect 86604 301608 91159 301610
rect 86604 301552 91098 301608
rect 91154 301552 91159 301608
rect 86604 301550 91159 301552
rect 86604 301548 86610 301550
rect 91093 301547 91159 301550
rect 122833 301610 122899 301613
rect 166942 301610 166948 301612
rect 122833 301608 166948 301610
rect 122833 301552 122838 301608
rect 122894 301552 166948 301608
rect 122833 301550 166948 301552
rect 122833 301547 122899 301550
rect 166942 301548 166948 301550
rect 167012 301548 167018 301612
rect 28993 301474 29059 301477
rect 169150 301474 169156 301476
rect 28993 301472 169156 301474
rect 28993 301416 28998 301472
rect 29054 301416 169156 301472
rect 28993 301414 169156 301416
rect 28993 301411 29059 301414
rect 169150 301412 169156 301414
rect 169220 301412 169226 301476
rect 226888 301474 226948 301683
rect 252686 301548 252692 301612
rect 252756 301610 252762 301612
rect 252921 301610 252987 301613
rect 252756 301608 252987 301610
rect 252756 301552 252926 301608
rect 252982 301552 252987 301608
rect 252756 301550 252987 301552
rect 252756 301548 252762 301550
rect 252921 301547 252987 301550
rect 259637 301474 259703 301477
rect 226888 301472 259703 301474
rect 226888 301416 259642 301472
rect 259698 301416 259703 301472
rect 226888 301414 259703 301416
rect 259637 301411 259703 301414
rect 152641 301202 152707 301205
rect 223757 301202 223823 301205
rect 152641 301200 223823 301202
rect 152641 301144 152646 301200
rect 152702 301144 223762 301200
rect 223818 301144 223823 301200
rect 152641 301142 223823 301144
rect 152641 301139 152707 301142
rect 223757 301139 223823 301142
rect 244774 301004 244780 301068
rect 244844 301066 244850 301068
rect 253430 301066 253490 301172
rect 287145 301066 287211 301069
rect 244844 301064 287211 301066
rect 244844 301008 287150 301064
rect 287206 301008 287211 301064
rect 244844 301006 287211 301008
rect 244844 301004 244850 301006
rect 287145 301003 287211 301006
rect 191465 300930 191531 300933
rect 195973 300930 196039 300933
rect 236729 300930 236795 300933
rect 191465 300928 193660 300930
rect 191465 300872 191470 300928
rect 191526 300872 193660 300928
rect 191465 300870 193660 300872
rect 195838 300928 196039 300930
rect 195838 300872 195978 300928
rect 196034 300872 196039 300928
rect 195838 300870 196039 300872
rect 191465 300867 191531 300870
rect 193489 300794 193555 300797
rect 195838 300794 195898 300870
rect 195973 300867 196039 300870
rect 236686 300928 236795 300930
rect 236686 300872 236734 300928
rect 236790 300872 236795 300928
rect 236686 300867 236795 300872
rect 249701 300930 249767 300933
rect 249701 300928 249810 300930
rect 249701 300872 249706 300928
rect 249762 300872 249810 300928
rect 249701 300867 249810 300872
rect 236686 300794 236746 300867
rect 193489 300792 195898 300794
rect 193489 300736 193494 300792
rect 193550 300736 195898 300792
rect 193489 300734 195898 300736
rect 219390 300734 236746 300794
rect 193489 300731 193555 300734
rect 115933 300250 115999 300253
rect 219390 300250 219450 300734
rect 248454 300732 248460 300796
rect 248524 300794 248530 300796
rect 249750 300794 249810 300867
rect 255497 300794 255563 300797
rect 248524 300734 249810 300794
rect 253460 300792 255563 300794
rect 253460 300736 255502 300792
rect 255558 300736 255563 300792
rect 253460 300734 255563 300736
rect 248524 300732 248530 300734
rect 249750 300658 249810 300734
rect 255497 300731 255563 300734
rect 261017 300658 261083 300661
rect 249750 300656 261083 300658
rect 249750 300600 261022 300656
rect 261078 300600 261083 300656
rect 249750 300598 261083 300600
rect 261017 300595 261083 300598
rect 255589 300386 255655 300389
rect 253460 300384 255655 300386
rect 253460 300328 255594 300384
rect 255650 300328 255655 300384
rect 253460 300326 255655 300328
rect 255589 300323 255655 300326
rect 115933 300248 219450 300250
rect 115933 300192 115938 300248
rect 115994 300192 219450 300248
rect 115933 300190 219450 300192
rect 115933 300187 115999 300190
rect 5533 300114 5599 300117
rect 193489 300114 193555 300117
rect 5533 300112 193555 300114
rect 5533 300056 5538 300112
rect 5594 300056 193494 300112
rect 193550 300056 193555 300112
rect 5533 300054 193555 300056
rect 5533 300051 5599 300054
rect 193489 300051 193555 300054
rect 193673 300114 193739 300117
rect 194726 300114 194732 300116
rect 193673 300112 194732 300114
rect 193673 300056 193678 300112
rect 193734 300056 194732 300112
rect 193673 300054 194732 300056
rect 193673 300051 193739 300054
rect 194726 300052 194732 300054
rect 194796 300052 194802 300116
rect 253062 299845 253122 299948
rect 253013 299840 253122 299845
rect 253289 299842 253355 299845
rect 189993 299570 190059 299573
rect 193630 299570 193690 299812
rect 253013 299784 253018 299840
rect 253074 299784 253122 299840
rect 253013 299782 253122 299784
rect 253246 299840 253355 299842
rect 253246 299784 253294 299840
rect 253350 299784 253355 299840
rect 253013 299779 253079 299782
rect 253246 299779 253355 299784
rect 189993 299568 193690 299570
rect 189993 299512 189998 299568
rect 190054 299512 193690 299568
rect 253246 299570 253306 299779
rect 262857 299570 262923 299573
rect 253246 299568 262923 299570
rect 253246 299540 262862 299568
rect 189993 299510 193690 299512
rect 253276 299512 262862 299540
rect 262918 299512 262923 299568
rect 253276 299510 262923 299512
rect 189993 299507 190059 299510
rect 262857 299507 262923 299510
rect 255497 299162 255563 299165
rect 253460 299160 255563 299162
rect 253460 299104 255502 299160
rect 255558 299104 255563 299160
rect 253460 299102 255563 299104
rect 255497 299099 255563 299102
rect 252829 299026 252895 299029
rect 252829 299024 252938 299026
rect 252829 298968 252834 299024
rect 252890 298968 252938 299024
rect 252829 298963 252938 298968
rect 193121 298890 193187 298893
rect 180750 298888 193187 298890
rect 180750 298832 193126 298888
rect 193182 298832 193187 298888
rect 180750 298830 193187 298832
rect 11053 298754 11119 298757
rect 180750 298754 180810 298830
rect 193121 298827 193187 298830
rect 11053 298752 180810 298754
rect 11053 298696 11058 298752
rect 11114 298696 180810 298752
rect 11053 298694 180810 298696
rect 191465 298754 191531 298757
rect 191465 298752 193660 298754
rect 191465 298696 191470 298752
rect 191526 298696 193660 298752
rect 191465 298694 193660 298696
rect 11053 298691 11119 298694
rect 191465 298691 191531 298694
rect 252878 298618 252938 298963
rect 255865 298754 255931 298757
rect 256734 298754 256740 298756
rect 255865 298752 256740 298754
rect 255865 298696 255870 298752
rect 255926 298696 256740 298752
rect 255865 298694 256740 298696
rect 255865 298691 255931 298694
rect 256734 298692 256740 298694
rect 256804 298754 256810 298756
rect 278773 298754 278839 298757
rect 583520 298754 584960 298844
rect 256804 298752 278839 298754
rect 256804 298696 278778 298752
rect 278834 298696 278839 298752
rect 256804 298694 278839 298696
rect 256804 298692 256810 298694
rect 278773 298691 278839 298694
rect 583342 298694 584960 298754
rect 255589 298618 255655 298621
rect 252878 298616 255655 298618
rect 252878 298588 255594 298616
rect 252908 298560 255594 298588
rect 255650 298560 255655 298616
rect 252908 298558 255655 298560
rect 583342 298618 583402 298694
rect 583520 298618 584960 298694
rect 583342 298604 584960 298618
rect 583342 298558 583586 298604
rect 255589 298555 255655 298558
rect 255497 298210 255563 298213
rect 253460 298208 255563 298210
rect 253460 298152 255502 298208
rect 255558 298152 255563 298208
rect 253460 298150 255563 298152
rect 255497 298147 255563 298150
rect 273110 298148 273116 298212
rect 273180 298210 273186 298212
rect 583526 298210 583586 298558
rect 273180 298150 583586 298210
rect 273180 298148 273186 298150
rect 127801 298074 127867 298077
rect 128261 298074 128327 298077
rect 176101 298074 176167 298077
rect 127801 298072 176167 298074
rect 127801 298016 127806 298072
rect 127862 298016 128266 298072
rect 128322 298016 176106 298072
rect 176162 298016 176167 298072
rect 127801 298014 176167 298016
rect 127801 298011 127867 298014
rect 128261 298011 128327 298014
rect 176101 298011 176167 298014
rect 252829 298074 252895 298077
rect 259269 298074 259335 298077
rect 265617 298074 265683 298077
rect 252829 298072 252938 298074
rect 252829 298016 252834 298072
rect 252890 298016 252938 298072
rect 252829 298011 252938 298016
rect 259269 298072 265683 298074
rect 259269 298016 259274 298072
rect 259330 298016 265622 298072
rect 265678 298016 265683 298072
rect 259269 298014 265683 298016
rect 259269 298011 259335 298014
rect 265617 298011 265683 298014
rect 252878 297802 252938 298011
rect 256049 297802 256115 297805
rect 252878 297800 256115 297802
rect 252878 297772 256054 297800
rect 252908 297744 256054 297772
rect 256110 297744 256115 297800
rect 252908 297742 256115 297744
rect 256049 297739 256115 297742
rect 191465 297666 191531 297669
rect 191465 297664 193660 297666
rect 191465 297608 191470 297664
rect 191526 297608 193660 297664
rect 191465 297606 193660 297608
rect 191465 297603 191531 297606
rect 27613 297394 27679 297397
rect 127801 297394 127867 297397
rect 27613 297392 127867 297394
rect 27613 297336 27618 297392
rect 27674 297336 127806 297392
rect 127862 297336 127867 297392
rect 27613 297334 127867 297336
rect 27613 297331 27679 297334
rect 127801 297331 127867 297334
rect 134701 297394 134767 297397
rect 186405 297394 186471 297397
rect 255865 297394 255931 297397
rect 134701 297392 186471 297394
rect 134701 297336 134706 297392
rect 134762 297336 186410 297392
rect 186466 297336 186471 297392
rect 134701 297334 186471 297336
rect 253460 297392 255931 297394
rect 253460 297336 255870 297392
rect 255926 297336 255931 297392
rect 253460 297334 255931 297336
rect 134701 297331 134767 297334
rect 186405 297331 186471 297334
rect 255865 297331 255931 297334
rect 186814 296924 186820 296988
rect 186884 296986 186890 296988
rect 192937 296986 193003 296989
rect 255497 296986 255563 296989
rect 186884 296984 193003 296986
rect 186884 296928 192942 296984
rect 192998 296928 193003 296984
rect 186884 296926 193003 296928
rect 253460 296984 255563 296986
rect 253460 296928 255502 296984
rect 255558 296928 255563 296984
rect 253460 296926 255563 296928
rect 186884 296924 186890 296926
rect 192937 296923 193003 296926
rect 255497 296923 255563 296926
rect 259678 296652 259684 296716
rect 259748 296714 259754 296716
rect 259821 296714 259887 296717
rect 259748 296712 259887 296714
rect 259748 296656 259826 296712
rect 259882 296656 259887 296712
rect 259748 296654 259887 296656
rect 259748 296652 259754 296654
rect 259821 296651 259887 296654
rect 255497 296578 255563 296581
rect 253460 296576 255563 296578
rect 192017 296034 192083 296037
rect 193630 296034 193690 296548
rect 253460 296520 255502 296576
rect 255558 296520 255563 296576
rect 253460 296518 255563 296520
rect 255497 296515 255563 296518
rect 255313 296170 255379 296173
rect 253460 296168 255379 296170
rect 253460 296112 255318 296168
rect 255374 296112 255379 296168
rect 253460 296110 255379 296112
rect 255313 296107 255379 296110
rect 192017 296032 193690 296034
rect 192017 295976 192022 296032
rect 192078 295976 193690 296032
rect 192017 295974 193690 295976
rect 192017 295971 192083 295974
rect 253933 295626 253999 295629
rect 253460 295624 253999 295626
rect 253460 295568 253938 295624
rect 253994 295568 253999 295624
rect 253460 295566 253999 295568
rect 253933 295563 253999 295566
rect 189901 295490 189967 295493
rect 255313 295490 255379 295493
rect 255681 295490 255747 295493
rect 189901 295488 193660 295490
rect 189901 295432 189906 295488
rect 189962 295432 193660 295488
rect 189901 295430 193660 295432
rect 255313 295488 255747 295490
rect 255313 295432 255318 295488
rect 255374 295432 255686 295488
rect 255742 295432 255747 295488
rect 255313 295430 255747 295432
rect 189901 295427 189967 295430
rect 255313 295427 255379 295430
rect 255681 295427 255747 295430
rect 141693 295354 141759 295357
rect 142061 295354 142127 295357
rect 192017 295354 192083 295357
rect 141693 295352 192083 295354
rect 141693 295296 141698 295352
rect 141754 295296 142066 295352
rect 142122 295296 192022 295352
rect 192078 295296 192083 295352
rect 141693 295294 192083 295296
rect 141693 295291 141759 295294
rect 142061 295291 142127 295294
rect 192017 295291 192083 295294
rect 148910 295156 148916 295220
rect 148980 295218 148986 295220
rect 193673 295218 193739 295221
rect 148980 295216 193739 295218
rect 148980 295160 193678 295216
rect 193734 295160 193739 295216
rect 148980 295158 193739 295160
rect 148980 295156 148986 295158
rect 193673 295155 193739 295158
rect 253430 295082 253490 295188
rect 256693 295082 256759 295085
rect 266445 295082 266511 295085
rect 253430 295080 266511 295082
rect 253430 295024 256698 295080
rect 256754 295024 266450 295080
rect 266506 295024 266511 295080
rect 253430 295022 266511 295024
rect 256693 295019 256759 295022
rect 266445 295019 266511 295022
rect 256693 294810 256759 294813
rect 253460 294808 256759 294810
rect 253460 294752 256698 294808
rect 256754 294752 256759 294808
rect 253460 294750 256759 294752
rect 256693 294747 256759 294750
rect 81934 294612 81940 294676
rect 82004 294674 82010 294676
rect 88425 294674 88491 294677
rect 82004 294672 88491 294674
rect 82004 294616 88430 294672
rect 88486 294616 88491 294672
rect 82004 294614 88491 294616
rect 82004 294612 82010 294614
rect 88425 294611 88491 294614
rect 4153 294538 4219 294541
rect 148910 294538 148916 294540
rect 4153 294536 148916 294538
rect 4153 294480 4158 294536
rect 4214 294480 148916 294536
rect 4153 294478 148916 294480
rect 4153 294475 4219 294478
rect 148910 294476 148916 294478
rect 148980 294476 148986 294540
rect 191465 294402 191531 294405
rect 255313 294402 255379 294405
rect 191465 294400 193660 294402
rect 191465 294344 191470 294400
rect 191526 294344 193660 294400
rect 191465 294342 193660 294344
rect 253460 294400 255379 294402
rect 253460 294344 255318 294400
rect 255374 294344 255379 294400
rect 253460 294342 255379 294344
rect 191465 294339 191531 294342
rect 255313 294339 255379 294342
rect 255405 293994 255471 293997
rect 253460 293992 255471 293994
rect 253460 293936 255410 293992
rect 255466 293936 255471 293992
rect 253460 293934 255471 293936
rect 255405 293931 255471 293934
rect 256785 293586 256851 293589
rect 253460 293584 256851 293586
rect 253460 293556 256790 293584
rect 253430 293528 256790 293556
rect 256846 293528 256851 293584
rect 253430 293526 256851 293528
rect 252829 293450 252895 293453
rect 253430 293450 253490 293526
rect 256785 293523 256851 293526
rect 252829 293448 253490 293450
rect 252829 293392 252834 293448
rect 252890 293392 253490 293448
rect 252829 293390 253490 293392
rect 252829 293387 252895 293390
rect 191465 293314 191531 293317
rect 191465 293312 193660 293314
rect -960 293178 480 293268
rect 191465 293256 191470 293312
rect 191526 293256 193660 293312
rect 191465 293254 193660 293256
rect 191465 293251 191531 293254
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 79961 293178 80027 293181
rect 87086 293178 87092 293180
rect 79961 293176 87092 293178
rect 79961 293120 79966 293176
rect 80022 293120 87092 293176
rect 79961 293118 87092 293120
rect 79961 293115 80027 293118
rect 87086 293116 87092 293118
rect 87156 293116 87162 293180
rect 255313 293178 255379 293181
rect 253460 293176 255379 293178
rect 253460 293148 255318 293176
rect 253430 293120 255318 293148
rect 255374 293120 255379 293176
rect 253430 293118 255379 293120
rect 253197 292906 253263 292909
rect 253430 292906 253490 293118
rect 255313 293115 255379 293118
rect 253197 292904 253490 292906
rect 253197 292848 253202 292904
rect 253258 292848 253490 292904
rect 253197 292846 253490 292848
rect 253197 292843 253263 292846
rect 255405 292634 255471 292637
rect 253460 292632 255471 292634
rect 253460 292576 255410 292632
rect 255466 292576 255471 292632
rect 253460 292574 255471 292576
rect 255405 292571 255471 292574
rect 191465 292226 191531 292229
rect 256601 292226 256667 292229
rect 191465 292224 193660 292226
rect 191465 292168 191470 292224
rect 191526 292168 193660 292224
rect 191465 292166 193660 292168
rect 253460 292224 256667 292226
rect 253460 292168 256606 292224
rect 256662 292168 256667 292224
rect 253460 292166 256667 292168
rect 191465 292163 191531 292166
rect 256601 292163 256667 292166
rect 182909 291954 182975 291957
rect 185342 291954 185348 291956
rect 182909 291952 185348 291954
rect 182909 291896 182914 291952
rect 182970 291896 185348 291952
rect 182909 291894 185348 291896
rect 182909 291891 182975 291894
rect 185342 291892 185348 291894
rect 185412 291892 185418 291956
rect 24853 291818 24919 291821
rect 192477 291818 192543 291821
rect 256601 291818 256667 291821
rect 24853 291816 192543 291818
rect 24853 291760 24858 291816
rect 24914 291760 192482 291816
rect 192538 291760 192543 291816
rect 24853 291758 192543 291760
rect 253460 291816 256667 291818
rect 253460 291760 256606 291816
rect 256662 291760 256667 291816
rect 253460 291758 256667 291760
rect 24853 291755 24919 291758
rect 192477 291755 192543 291758
rect 256601 291755 256667 291758
rect 260966 291682 260972 291684
rect 253430 291622 260972 291682
rect 253430 291380 253490 291622
rect 260966 291620 260972 291622
rect 261036 291620 261042 291684
rect 260966 291212 260972 291276
rect 261036 291274 261042 291276
rect 261201 291274 261267 291277
rect 261036 291272 261267 291274
rect 261036 291216 261206 291272
rect 261262 291216 261267 291272
rect 261036 291214 261267 291216
rect 261036 291212 261042 291214
rect 261201 291211 261267 291214
rect 68870 291076 68876 291140
rect 68940 291138 68946 291140
rect 69657 291138 69723 291141
rect 68940 291136 69723 291138
rect 68940 291080 69662 291136
rect 69718 291080 69723 291136
rect 68940 291078 69723 291080
rect 68940 291076 68946 291078
rect 69657 291075 69723 291078
rect 78438 291076 78444 291140
rect 78508 291138 78514 291140
rect 80053 291138 80119 291141
rect 78508 291136 80119 291138
rect 78508 291080 80058 291136
rect 80114 291080 80119 291136
rect 78508 291078 80119 291080
rect 78508 291076 78514 291078
rect 80053 291075 80119 291078
rect 80646 291076 80652 291140
rect 80716 291138 80722 291140
rect 82077 291138 82143 291141
rect 80716 291136 82143 291138
rect 80716 291080 82082 291136
rect 82138 291080 82143 291136
rect 80716 291078 82143 291080
rect 80716 291076 80722 291078
rect 82077 291075 82143 291078
rect 87321 291138 87387 291141
rect 88241 291138 88307 291141
rect 87321 291136 88307 291138
rect 87321 291080 87326 291136
rect 87382 291080 88246 291136
rect 88302 291080 88307 291136
rect 87321 291078 88307 291080
rect 87321 291075 87387 291078
rect 88241 291075 88307 291078
rect 191465 291138 191531 291141
rect 191465 291136 193660 291138
rect 191465 291080 191470 291136
rect 191526 291080 193660 291136
rect 191465 291078 193660 291080
rect 191465 291075 191531 291078
rect 256509 291002 256575 291005
rect 253460 291000 256575 291002
rect 253460 290944 256514 291000
rect 256570 290944 256575 291000
rect 253460 290942 256575 290944
rect 256509 290939 256575 290942
rect 256509 290594 256575 290597
rect 253460 290592 256575 290594
rect 253460 290536 256514 290592
rect 256570 290536 256575 290592
rect 253460 290534 256575 290536
rect 256509 290531 256575 290534
rect 3417 290458 3483 290461
rect 87597 290458 87663 290461
rect 3417 290456 87663 290458
rect 3417 290400 3422 290456
rect 3478 290400 87602 290456
rect 87658 290400 87663 290456
rect 3417 290398 87663 290400
rect 3417 290395 3483 290398
rect 87597 290395 87663 290398
rect 163957 290458 164023 290461
rect 186037 290458 186103 290461
rect 163957 290456 186103 290458
rect 163957 290400 163962 290456
rect 164018 290400 186042 290456
rect 186098 290400 186103 290456
rect 163957 290398 186103 290400
rect 163957 290395 164023 290398
rect 186037 290395 186103 290398
rect 91502 289988 91508 290052
rect 91572 290050 91578 290052
rect 95233 290050 95299 290053
rect 91572 290048 95299 290050
rect 91572 289992 95238 290048
rect 95294 289992 95299 290048
rect 91572 289990 95299 289992
rect 91572 289988 91578 289990
rect 95233 289987 95299 289990
rect 190821 290050 190887 290053
rect 258574 290050 258580 290052
rect 190821 290048 193660 290050
rect 190821 289992 190826 290048
rect 190882 289992 193660 290048
rect 190821 289990 193660 289992
rect 253460 289990 258580 290050
rect 190821 289987 190887 289990
rect 258574 289988 258580 289990
rect 258644 289988 258650 290052
rect 87321 289914 87387 289917
rect 100109 289914 100175 289917
rect 87321 289912 100175 289914
rect 87321 289856 87326 289912
rect 87382 289856 100114 289912
rect 100170 289856 100175 289912
rect 87321 289854 100175 289856
rect 87321 289851 87387 289854
rect 100109 289851 100175 289854
rect 63309 289778 63375 289781
rect 153101 289778 153167 289781
rect 63309 289776 153167 289778
rect 63309 289720 63314 289776
rect 63370 289720 153106 289776
rect 153162 289720 153167 289776
rect 63309 289718 153167 289720
rect 63309 289715 63375 289718
rect 153101 289715 153167 289718
rect 88006 289580 88012 289644
rect 88076 289642 88082 289644
rect 89713 289642 89779 289645
rect 256509 289642 256575 289645
rect 88076 289640 89779 289642
rect 88076 289584 89718 289640
rect 89774 289584 89779 289640
rect 88076 289582 89779 289584
rect 253460 289640 256575 289642
rect 253460 289584 256514 289640
rect 256570 289584 256575 289640
rect 253460 289582 256575 289584
rect 88076 289580 88082 289582
rect 89713 289579 89779 289582
rect 256509 289579 256575 289582
rect 256601 289234 256667 289237
rect 253460 289232 256667 289234
rect 253460 289176 256606 289232
rect 256662 289176 256667 289232
rect 253460 289174 256667 289176
rect 256601 289171 256667 289174
rect 153101 289098 153167 289101
rect 180241 289098 180307 289101
rect 153101 289096 180307 289098
rect 153101 289040 153106 289096
rect 153162 289040 180246 289096
rect 180302 289040 180307 289096
rect 153101 289038 180307 289040
rect 153101 289035 153167 289038
rect 180241 289035 180307 289038
rect 191465 288962 191531 288965
rect 191465 288960 193660 288962
rect 191465 288904 191470 288960
rect 191526 288904 193660 288960
rect 191465 288902 193660 288904
rect 191465 288899 191531 288902
rect 259494 288826 259500 288828
rect 253460 288766 259500 288826
rect 259494 288764 259500 288766
rect 259564 288764 259570 288828
rect 74625 288690 74691 288693
rect 79174 288690 79180 288692
rect 74625 288688 79180 288690
rect 74625 288632 74630 288688
rect 74686 288632 79180 288688
rect 74625 288630 79180 288632
rect 74625 288627 74691 288630
rect 79174 288628 79180 288630
rect 79244 288628 79250 288692
rect 69013 288554 69079 288557
rect 74758 288554 74764 288556
rect 69013 288552 74764 288554
rect 69013 288496 69018 288552
rect 69074 288496 74764 288552
rect 69013 288494 74764 288496
rect 69013 288491 69079 288494
rect 74758 288492 74764 288494
rect 74828 288492 74834 288556
rect 173893 288418 173959 288421
rect 174629 288418 174695 288421
rect 256969 288418 257035 288421
rect 257981 288418 258047 288421
rect 173893 288416 174695 288418
rect 173893 288360 173898 288416
rect 173954 288360 174634 288416
rect 174690 288360 174695 288416
rect 173893 288358 174695 288360
rect 253460 288416 258047 288418
rect 253460 288360 256974 288416
rect 257030 288360 257986 288416
rect 258042 288360 258047 288416
rect 253460 288358 258047 288360
rect 173893 288355 173959 288358
rect 174629 288355 174695 288358
rect 256969 288355 257035 288358
rect 257981 288355 258047 288358
rect 255865 288010 255931 288013
rect 253460 288008 255931 288010
rect 253460 287952 255870 288008
rect 255926 287952 255931 288008
rect 253460 287950 255931 287952
rect 255865 287947 255931 287950
rect 88609 287874 88675 287877
rect 99966 287874 99972 287876
rect 88609 287872 99972 287874
rect 88609 287816 88614 287872
rect 88670 287816 99972 287872
rect 88609 287814 99972 287816
rect 88609 287811 88675 287814
rect 99966 287812 99972 287814
rect 100036 287812 100042 287876
rect 191465 287874 191531 287877
rect 191465 287872 193660 287874
rect 191465 287816 191470 287872
rect 191526 287816 193660 287872
rect 191465 287814 193660 287816
rect 191465 287811 191531 287814
rect 64597 287738 64663 287741
rect 64781 287738 64847 287741
rect 173893 287738 173959 287741
rect 64597 287736 173959 287738
rect 64597 287680 64602 287736
rect 64658 287680 64786 287736
rect 64842 287680 173898 287736
rect 173954 287680 173959 287736
rect 64597 287678 173959 287680
rect 64597 287675 64663 287678
rect 64781 287675 64847 287678
rect 173893 287675 173959 287678
rect 257981 287738 258047 287741
rect 267733 287738 267799 287741
rect 257981 287736 267799 287738
rect 257981 287680 257986 287736
rect 258042 287680 267738 287736
rect 267794 287680 267799 287736
rect 257981 287678 267799 287680
rect 257981 287675 258047 287678
rect 267733 287675 267799 287678
rect 255957 287602 256023 287605
rect 253460 287600 256023 287602
rect 253460 287544 255962 287600
rect 256018 287544 256023 287600
rect 253460 287542 256023 287544
rect 255957 287539 256023 287542
rect 69841 287194 69907 287197
rect 74942 287194 74948 287196
rect 69841 287192 74948 287194
rect 69841 287136 69846 287192
rect 69902 287136 74948 287192
rect 69841 287134 74948 287136
rect 69841 287131 69907 287134
rect 74942 287132 74948 287134
rect 75012 287132 75018 287196
rect 253430 286922 253490 287028
rect 253430 286862 263610 286922
rect 191373 286786 191439 286789
rect 191373 286784 193660 286786
rect 191373 286728 191378 286784
rect 191434 286728 193660 286784
rect 191373 286726 193660 286728
rect 191373 286723 191439 286726
rect 255865 286650 255931 286653
rect 253460 286648 255931 286650
rect 253460 286592 255870 286648
rect 255926 286592 255931 286648
rect 253460 286590 255931 286592
rect 255865 286587 255931 286590
rect 142981 286378 143047 286381
rect 187049 286378 187115 286381
rect 142981 286376 187115 286378
rect 142981 286320 142986 286376
rect 143042 286320 187054 286376
rect 187110 286320 187115 286376
rect 142981 286318 187115 286320
rect 142981 286315 143047 286318
rect 187049 286315 187115 286318
rect 256509 286242 256575 286245
rect 253460 286240 256575 286242
rect 253460 286184 256514 286240
rect 256570 286184 256575 286240
rect 253460 286182 256575 286184
rect 256509 286179 256575 286182
rect 90265 286106 90331 286109
rect 91001 286106 91067 286109
rect 90265 286104 91067 286106
rect 90265 286048 90270 286104
rect 90326 286048 91006 286104
rect 91062 286048 91067 286104
rect 90265 286046 91067 286048
rect 263550 286106 263610 286862
rect 268326 286106 268332 286108
rect 263550 286046 268332 286106
rect 90265 286043 90331 286046
rect 91001 286043 91067 286046
rect 268326 286044 268332 286046
rect 268396 286044 268402 286108
rect 89161 285970 89227 285973
rect 148593 285970 148659 285973
rect 89161 285968 148659 285970
rect 89161 285912 89166 285968
rect 89222 285912 148598 285968
rect 148654 285912 148659 285968
rect 89161 285910 148659 285912
rect 89161 285907 89227 285910
rect 148593 285907 148659 285910
rect 46841 285834 46907 285837
rect 73797 285834 73863 285837
rect 46841 285832 73863 285834
rect 46841 285776 46846 285832
rect 46902 285776 73802 285832
rect 73858 285776 73863 285832
rect 46841 285774 73863 285776
rect 46841 285771 46907 285774
rect 73797 285771 73863 285774
rect 83089 285834 83155 285837
rect 84009 285834 84075 285837
rect 116669 285834 116735 285837
rect 266629 285834 266695 285837
rect 83089 285832 116735 285834
rect 83089 285776 83094 285832
rect 83150 285776 84014 285832
rect 84070 285776 116674 285832
rect 116730 285776 116735 285832
rect 83089 285774 116735 285776
rect 253460 285832 267750 285834
rect 253460 285776 266634 285832
rect 266690 285776 267750 285832
rect 253460 285774 267750 285776
rect 83089 285771 83155 285774
rect 84009 285771 84075 285774
rect 116669 285771 116735 285774
rect 266629 285771 266695 285774
rect 83406 285636 83412 285700
rect 83476 285698 83482 285700
rect 84101 285698 84167 285701
rect 83476 285696 84167 285698
rect 83476 285640 84106 285696
rect 84162 285640 84167 285696
rect 83476 285638 84167 285640
rect 83476 285636 83482 285638
rect 84101 285635 84167 285638
rect 86718 285636 86724 285700
rect 86788 285698 86794 285700
rect 86861 285698 86927 285701
rect 86788 285696 86927 285698
rect 86788 285640 86866 285696
rect 86922 285640 86927 285696
rect 86788 285638 86927 285640
rect 86788 285636 86794 285638
rect 86861 285635 86927 285638
rect 166758 285636 166764 285700
rect 166828 285698 166834 285700
rect 167085 285698 167151 285701
rect 166828 285696 167151 285698
rect 166828 285640 167090 285696
rect 167146 285640 167151 285696
rect 166828 285638 167151 285640
rect 166828 285636 166834 285638
rect 167085 285635 167151 285638
rect 191465 285698 191531 285701
rect 267690 285698 267750 285774
rect 268326 285772 268332 285836
rect 268396 285834 268402 285836
rect 276238 285834 276244 285836
rect 268396 285774 276244 285834
rect 268396 285772 268402 285774
rect 276238 285772 276244 285774
rect 276308 285772 276314 285836
rect 269113 285698 269179 285701
rect 191465 285696 193660 285698
rect 191465 285640 191470 285696
rect 191526 285640 193660 285696
rect 191465 285638 193660 285640
rect 267690 285696 269179 285698
rect 267690 285640 269118 285696
rect 269174 285640 269179 285696
rect 267690 285638 269179 285640
rect 191465 285635 191531 285638
rect 269113 285635 269179 285638
rect 256601 285426 256667 285429
rect 253460 285424 256667 285426
rect 253460 285368 256606 285424
rect 256662 285368 256667 285424
rect 253460 285366 256667 285368
rect 256601 285363 256667 285366
rect 262213 285290 262279 285293
rect 263133 285290 263199 285293
rect 253430 285288 263199 285290
rect 253430 285232 262218 285288
rect 262274 285232 263138 285288
rect 263194 285232 263199 285288
rect 583520 285276 584960 285516
rect 253430 285230 263199 285232
rect 148409 285018 148475 285021
rect 186262 285018 186268 285020
rect 148409 285016 186268 285018
rect 148409 284960 148414 285016
rect 148470 284960 186268 285016
rect 148409 284958 186268 284960
rect 148409 284955 148475 284958
rect 186262 284956 186268 284958
rect 186332 284956 186338 285020
rect 253430 284988 253490 285230
rect 262213 285227 262279 285230
rect 263133 285227 263199 285230
rect 61745 284882 61811 284885
rect 165613 284882 165679 284885
rect 61745 284880 165679 284882
rect 61745 284824 61750 284880
rect 61806 284824 165618 284880
rect 165674 284824 165679 284880
rect 61745 284822 165679 284824
rect 61745 284819 61811 284822
rect 165613 284819 165679 284822
rect 191465 284610 191531 284613
rect 191465 284608 193660 284610
rect 191465 284552 191470 284608
rect 191526 284552 193660 284608
rect 191465 284550 193660 284552
rect 253460 284550 263978 284610
rect 191465 284547 191531 284550
rect 93945 284338 94011 284341
rect 137553 284338 137619 284341
rect 93945 284336 137619 284338
rect 93945 284280 93950 284336
rect 94006 284280 137558 284336
rect 137614 284280 137619 284336
rect 93945 284278 137619 284280
rect 93945 284275 94011 284278
rect 137553 284275 137619 284278
rect 165613 284338 165679 284341
rect 166441 284338 166507 284341
rect 165613 284336 166507 284338
rect 165613 284280 165618 284336
rect 165674 284280 166446 284336
rect 166502 284280 166507 284336
rect 165613 284278 166507 284280
rect 165613 284275 165679 284278
rect 166441 284275 166507 284278
rect 263133 284338 263199 284341
rect 263685 284338 263751 284341
rect 263133 284336 263751 284338
rect 263133 284280 263138 284336
rect 263194 284280 263690 284336
rect 263746 284280 263751 284336
rect 263133 284278 263751 284280
rect 263918 284338 263978 284550
rect 266353 284338 266419 284341
rect 266721 284338 266787 284341
rect 263918 284336 266787 284338
rect 263918 284280 266358 284336
rect 266414 284280 266726 284336
rect 266782 284280 266787 284336
rect 263918 284278 266787 284280
rect 263133 284275 263199 284278
rect 263685 284275 263751 284278
rect 266353 284275 266419 284278
rect 266721 284275 266787 284278
rect 73470 284140 73476 284204
rect 73540 284202 73546 284204
rect 73889 284202 73955 284205
rect 73540 284200 73955 284202
rect 73540 284144 73894 284200
rect 73950 284144 73955 284200
rect 73540 284142 73955 284144
rect 73540 284140 73546 284142
rect 73889 284139 73955 284142
rect 75678 284140 75684 284204
rect 75748 284202 75754 284204
rect 76557 284202 76623 284205
rect 75748 284200 76623 284202
rect 75748 284144 76562 284200
rect 76618 284144 76623 284200
rect 75748 284142 76623 284144
rect 75748 284140 75754 284142
rect 76557 284139 76623 284142
rect 78254 284140 78260 284204
rect 78324 284202 78330 284204
rect 78673 284202 78739 284205
rect 78324 284200 78739 284202
rect 78324 284144 78678 284200
rect 78734 284144 78739 284200
rect 78324 284142 78739 284144
rect 78324 284140 78330 284142
rect 78673 284139 78739 284142
rect 91134 284140 91140 284204
rect 91204 284202 91210 284204
rect 92289 284202 92355 284205
rect 91204 284200 92355 284202
rect 91204 284144 92294 284200
rect 92350 284144 92355 284200
rect 91204 284142 92355 284144
rect 91204 284140 91210 284142
rect 92289 284139 92355 284142
rect 253430 283930 253490 284036
rect 262213 283930 262279 283933
rect 253430 283928 262279 283930
rect 253430 283872 262218 283928
rect 262274 283872 262279 283928
rect 253430 283870 262279 283872
rect 262213 283867 262279 283870
rect 71865 283658 71931 283661
rect 72417 283658 72483 283661
rect 71865 283656 72483 283658
rect 71865 283600 71870 283656
rect 71926 283600 72422 283656
rect 72478 283600 72483 283656
rect 71865 283598 72483 283600
rect 71865 283595 71931 283598
rect 72417 283595 72483 283598
rect 92381 283658 92447 283661
rect 255773 283658 255839 283661
rect 92381 283656 99390 283658
rect 92381 283600 92386 283656
rect 92442 283600 99390 283656
rect 92381 283598 99390 283600
rect 253460 283656 255839 283658
rect 253460 283600 255778 283656
rect 255834 283600 255839 283656
rect 253460 283598 255839 283600
rect 92381 283595 92447 283598
rect 71589 283522 71655 283525
rect 64830 283520 71655 283522
rect 64830 283464 71594 283520
rect 71650 283464 71655 283520
rect 64830 283462 71655 283464
rect 64830 283389 64890 283462
rect 71589 283459 71655 283462
rect 71814 283460 71820 283524
rect 71884 283522 71890 283524
rect 71957 283522 72023 283525
rect 73245 283524 73311 283525
rect 73245 283522 73292 283524
rect 71884 283520 72023 283522
rect 71884 283464 71962 283520
rect 72018 283464 72023 283520
rect 71884 283462 72023 283464
rect 73200 283520 73292 283522
rect 73200 283464 73250 283520
rect 73200 283462 73292 283464
rect 71884 283460 71890 283462
rect 71957 283459 72023 283462
rect 73245 283460 73292 283462
rect 73356 283460 73362 283524
rect 75310 283460 75316 283524
rect 75380 283522 75386 283524
rect 75821 283522 75887 283525
rect 75380 283520 75887 283522
rect 75380 283464 75826 283520
rect 75882 283464 75887 283520
rect 75380 283462 75887 283464
rect 75380 283460 75386 283462
rect 73245 283459 73311 283460
rect 75821 283459 75887 283462
rect 76966 283460 76972 283524
rect 77036 283522 77042 283524
rect 79041 283522 79107 283525
rect 77036 283520 79107 283522
rect 77036 283464 79046 283520
rect 79102 283464 79107 283520
rect 77036 283462 79107 283464
rect 77036 283460 77042 283462
rect 79041 283459 79107 283462
rect 89805 283524 89871 283525
rect 89805 283520 89852 283524
rect 89916 283522 89922 283524
rect 89805 283464 89810 283520
rect 89805 283460 89852 283464
rect 89916 283462 89962 283522
rect 89916 283460 89922 283462
rect 93342 283460 93348 283524
rect 93412 283522 93418 283524
rect 94037 283522 94103 283525
rect 93412 283520 94103 283522
rect 93412 283464 94042 283520
rect 94098 283464 94103 283520
rect 93412 283462 94103 283464
rect 93412 283460 93418 283462
rect 89805 283459 89871 283460
rect 94037 283459 94103 283462
rect 64781 283384 64890 283389
rect 64781 283328 64786 283384
rect 64842 283328 64890 283384
rect 64781 283326 64890 283328
rect 64781 283323 64847 283326
rect 67582 283324 67588 283388
rect 67652 283386 67658 283388
rect 67652 283326 80070 283386
rect 67652 283324 67658 283326
rect 67817 283250 67883 283253
rect 69054 283250 69060 283252
rect 67817 283248 69060 283250
rect 67817 283192 67822 283248
rect 67878 283192 69060 283248
rect 67817 283190 69060 283192
rect 67817 283187 67883 283190
rect 69054 283188 69060 283190
rect 69124 283188 69130 283252
rect 71865 283250 71931 283253
rect 69430 283248 71931 283250
rect 69430 283192 71870 283248
rect 71926 283192 71931 283248
rect 69430 283190 71931 283192
rect 80010 283250 80070 283326
rect 94078 283324 94084 283388
rect 94148 283386 94154 283388
rect 94681 283386 94747 283389
rect 94148 283384 94747 283386
rect 94148 283328 94686 283384
rect 94742 283328 94747 283384
rect 94148 283326 94747 283328
rect 94148 283324 94154 283326
rect 94681 283323 94747 283326
rect 96889 283386 96955 283389
rect 97758 283386 97764 283388
rect 96889 283384 97764 283386
rect 96889 283328 96894 283384
rect 96950 283328 97764 283384
rect 96889 283326 97764 283328
rect 96889 283323 96955 283326
rect 97758 283324 97764 283326
rect 97828 283324 97834 283388
rect 99330 283386 99390 283598
rect 255773 283595 255839 283598
rect 269757 283658 269823 283661
rect 281758 283658 281764 283660
rect 269757 283656 281764 283658
rect 269757 283600 269762 283656
rect 269818 283600 281764 283656
rect 269757 283598 281764 283600
rect 269757 283595 269823 283598
rect 281758 283596 281764 283598
rect 281828 283596 281834 283660
rect 145649 283522 145715 283525
rect 182909 283522 182975 283525
rect 145649 283520 182975 283522
rect 145649 283464 145654 283520
rect 145710 283464 182914 283520
rect 182970 283464 182975 283520
rect 145649 283462 182975 283464
rect 145649 283459 145715 283462
rect 182909 283459 182975 283462
rect 193121 283522 193187 283525
rect 259361 283522 259427 283525
rect 274909 283522 274975 283525
rect 193121 283520 193660 283522
rect 193121 283464 193126 283520
rect 193182 283464 193660 283520
rect 193121 283462 193660 283464
rect 259361 283520 274975 283522
rect 259361 283464 259366 283520
rect 259422 283464 274914 283520
rect 274970 283464 274975 283520
rect 259361 283462 274975 283464
rect 193121 283459 193187 283462
rect 259361 283459 259427 283462
rect 274909 283459 274975 283462
rect 100201 283386 100267 283389
rect 99330 283384 100267 283386
rect 99330 283328 100206 283384
rect 100262 283328 100267 283384
rect 99330 283326 100267 283328
rect 100201 283323 100267 283326
rect 112529 283250 112595 283253
rect 256417 283250 256483 283253
rect 80010 283248 112595 283250
rect 80010 283192 112534 283248
rect 112590 283192 112595 283248
rect 80010 283190 112595 283192
rect 253460 283248 256483 283250
rect 253460 283192 256422 283248
rect 256478 283192 256483 283248
rect 253460 283190 256483 283192
rect 57697 283114 57763 283117
rect 69430 283114 69490 283190
rect 71865 283187 71931 283190
rect 112529 283187 112595 283190
rect 256417 283187 256483 283190
rect 57697 283112 69490 283114
rect 57697 283056 57702 283112
rect 57758 283056 69490 283112
rect 57697 283054 69490 283056
rect 57697 283051 57763 283054
rect 69430 282948 69490 283054
rect 79910 283052 79916 283116
rect 79980 283114 79986 283116
rect 81985 283114 82051 283117
rect 79980 283112 82051 283114
rect 79980 283056 81990 283112
rect 82046 283056 82051 283112
rect 79980 283054 82051 283056
rect 79980 283052 79986 283054
rect 81985 283051 82051 283054
rect 84694 283052 84700 283116
rect 84764 283114 84770 283116
rect 88425 283114 88491 283117
rect 84764 283112 88491 283114
rect 84764 283056 88430 283112
rect 88486 283056 88491 283112
rect 84764 283054 88491 283056
rect 84764 283052 84770 283054
rect 88425 283051 88491 283054
rect 70158 282916 70164 282980
rect 70228 282978 70234 282980
rect 70853 282978 70919 282981
rect 70228 282976 70919 282978
rect 70228 282920 70858 282976
rect 70914 282920 70919 282976
rect 70228 282918 70919 282920
rect 70228 282916 70234 282918
rect 70853 282915 70919 282918
rect 81985 282978 82051 282981
rect 82629 282980 82695 282981
rect 83457 282980 83523 282981
rect 82629 282978 82676 282980
rect 81985 282976 82676 282978
rect 81985 282920 81990 282976
rect 82046 282920 82634 282976
rect 81985 282918 82676 282920
rect 81985 282915 82051 282918
rect 82629 282916 82676 282918
rect 82740 282916 82746 282980
rect 83406 282916 83412 282980
rect 83476 282978 83523 282980
rect 86309 282978 86375 282981
rect 86718 282978 86724 282980
rect 83476 282976 83568 282978
rect 83518 282920 83568 282976
rect 83476 282918 83568 282920
rect 86309 282976 86724 282978
rect 86309 282920 86314 282976
rect 86370 282920 86724 282976
rect 86309 282918 86724 282920
rect 83476 282916 83523 282918
rect 82629 282915 82695 282916
rect 83457 282915 83523 282916
rect 86309 282915 86375 282918
rect 86718 282916 86724 282918
rect 86788 282916 86794 282980
rect 88742 282916 88748 282980
rect 88812 282978 88818 282980
rect 89069 282978 89135 282981
rect 88812 282976 89135 282978
rect 88812 282920 89074 282976
rect 89130 282920 89135 282976
rect 88812 282918 89135 282920
rect 88812 282916 88818 282918
rect 89069 282915 89135 282918
rect 90725 282978 90791 282981
rect 98913 282978 98979 282981
rect 90725 282976 98979 282978
rect 90725 282920 90730 282976
rect 90786 282920 98918 282976
rect 98974 282920 98979 282976
rect 90725 282918 98979 282920
rect 90725 282915 90791 282918
rect 98913 282915 98979 282918
rect 259361 282842 259427 282845
rect 253460 282840 259427 282842
rect 253460 282784 259366 282840
rect 259422 282784 259427 282840
rect 253460 282782 259427 282784
rect 259361 282779 259427 282782
rect 100845 282706 100911 282709
rect 98716 282704 100911 282706
rect 98716 282648 100850 282704
rect 100906 282648 100911 282704
rect 98716 282646 100911 282648
rect 100845 282643 100911 282646
rect 191465 282434 191531 282437
rect 255497 282434 255563 282437
rect 191465 282432 193660 282434
rect 191465 282376 191470 282432
rect 191526 282376 193660 282432
rect 191465 282374 193660 282376
rect 253460 282432 255563 282434
rect 253460 282376 255502 282432
rect 255558 282376 255563 282432
rect 253460 282374 255563 282376
rect 191465 282371 191531 282374
rect 255497 282371 255563 282374
rect 258717 282298 258783 282301
rect 259453 282298 259519 282301
rect 258717 282296 259519 282298
rect 258717 282240 258722 282296
rect 258778 282240 259458 282296
rect 259514 282240 259519 282296
rect 258717 282238 259519 282240
rect 258717 282235 258783 282238
rect 259453 282235 259519 282238
rect 67265 282162 67331 282165
rect 260097 282162 260163 282165
rect 270585 282162 270651 282165
rect 292665 282162 292731 282165
rect 67265 282160 68908 282162
rect 67265 282104 67270 282160
rect 67326 282104 68908 282160
rect 67265 282102 68908 282104
rect 260097 282160 292731 282162
rect 260097 282104 260102 282160
rect 260158 282104 270590 282160
rect 270646 282104 292670 282160
rect 292726 282104 292731 282160
rect 260097 282102 292731 282104
rect 67265 282099 67331 282102
rect 260097 282099 260163 282102
rect 270585 282099 270651 282102
rect 292665 282099 292731 282102
rect 255405 282026 255471 282029
rect 253460 282024 255471 282026
rect 253460 281968 255410 282024
rect 255466 281968 255471 282024
rect 253460 281966 255471 281968
rect 255405 281963 255471 281966
rect 100753 281890 100819 281893
rect 98716 281888 100819 281890
rect 98716 281832 100758 281888
rect 100814 281832 100819 281888
rect 98716 281830 100819 281832
rect 100753 281827 100819 281830
rect 103329 281482 103395 281485
rect 115289 281482 115355 281485
rect 255405 281482 255471 281485
rect 103329 281480 115355 281482
rect 103329 281424 103334 281480
rect 103390 281424 115294 281480
rect 115350 281424 115355 281480
rect 103329 281422 115355 281424
rect 253460 281480 255471 281482
rect 253460 281424 255410 281480
rect 255466 281424 255471 281480
rect 253460 281422 255471 281424
rect 103329 281419 103395 281422
rect 115289 281419 115355 281422
rect 255405 281419 255471 281422
rect 270585 281482 270651 281485
rect 273253 281482 273319 281485
rect 270585 281480 273319 281482
rect 270585 281424 270590 281480
rect 270646 281424 273258 281480
rect 273314 281424 273319 281480
rect 270585 281422 273319 281424
rect 270585 281419 270651 281422
rect 273253 281419 273319 281422
rect 67265 281346 67331 281349
rect 67541 281346 67607 281349
rect 191465 281346 191531 281349
rect 67265 281344 68908 281346
rect 67265 281288 67270 281344
rect 67326 281288 67546 281344
rect 67602 281288 68908 281344
rect 67265 281286 68908 281288
rect 191465 281344 193660 281346
rect 191465 281288 191470 281344
rect 191526 281288 193660 281344
rect 191465 281286 193660 281288
rect 67265 281283 67331 281286
rect 67541 281283 67607 281286
rect 191465 281283 191531 281286
rect 100845 281074 100911 281077
rect 259637 281074 259703 281077
rect 262581 281074 262647 281077
rect 98716 281072 100911 281074
rect 98716 281016 100850 281072
rect 100906 281016 100911 281072
rect 98716 281014 100911 281016
rect 253460 281072 262647 281074
rect 253460 281016 259642 281072
rect 259698 281016 262586 281072
rect 262642 281016 262647 281072
rect 253460 281014 262647 281016
rect 100845 281011 100911 281014
rect 259637 281011 259703 281014
rect 262581 281011 262647 281014
rect 270585 280666 270651 280669
rect 253460 280664 270651 280666
rect 253460 280608 270590 280664
rect 270646 280608 270651 280664
rect 253460 280606 270651 280608
rect 270585 280603 270651 280606
rect 65926 280468 65932 280532
rect 65996 280530 66002 280532
rect 65996 280470 68908 280530
rect 65996 280468 66002 280470
rect 99966 280258 99972 280260
rect -960 279972 480 280212
rect 98716 280198 99972 280258
rect 99966 280196 99972 280198
rect 100036 280258 100042 280260
rect 103329 280258 103395 280261
rect 100036 280256 103395 280258
rect 100036 280200 103334 280256
rect 103390 280200 103395 280256
rect 100036 280198 103395 280200
rect 100036 280196 100042 280198
rect 103329 280195 103395 280198
rect 191465 280258 191531 280261
rect 255497 280258 255563 280261
rect 191465 280256 193660 280258
rect 191465 280200 191470 280256
rect 191526 280200 193660 280256
rect 191465 280198 193660 280200
rect 253460 280256 255563 280258
rect 253460 280200 255502 280256
rect 255558 280200 255563 280256
rect 253460 280198 255563 280200
rect 191465 280195 191531 280198
rect 255497 280195 255563 280198
rect 259453 279850 259519 279853
rect 253460 279848 267750 279850
rect 253460 279792 259458 279848
rect 259514 279792 267750 279848
rect 253460 279790 267750 279792
rect 259453 279787 259519 279790
rect 65885 279714 65951 279717
rect 263961 279714 264027 279717
rect 65885 279712 68908 279714
rect 65885 279656 65890 279712
rect 65946 279656 68908 279712
rect 65885 279654 68908 279656
rect 253430 279712 264027 279714
rect 253430 279656 263966 279712
rect 264022 279656 264027 279712
rect 253430 279654 264027 279656
rect 65885 279651 65951 279654
rect 100753 279442 100819 279445
rect 98716 279440 100819 279442
rect 98716 279384 100758 279440
rect 100814 279384 100819 279440
rect 253430 279412 253490 279654
rect 263961 279651 264027 279654
rect 267690 279442 267750 279790
rect 274817 279442 274883 279445
rect 267690 279440 274883 279442
rect 98716 279382 100819 279384
rect 267690 279384 274822 279440
rect 274878 279384 274883 279440
rect 267690 279382 274883 279384
rect 100753 279379 100819 279382
rect 274817 279379 274883 279382
rect 191465 279170 191531 279173
rect 191465 279168 193660 279170
rect 191465 279112 191470 279168
rect 191526 279112 193660 279168
rect 191465 279110 193660 279112
rect 191465 279107 191531 279110
rect 255405 279034 255471 279037
rect 253460 279032 255471 279034
rect 253460 278976 255410 279032
rect 255466 278976 255471 279032
rect 253460 278974 255471 278976
rect 255405 278971 255471 278974
rect 66805 278898 66871 278901
rect 66805 278896 68908 278898
rect 66805 278840 66810 278896
rect 66866 278840 68908 278896
rect 66805 278838 68908 278840
rect 66805 278835 66871 278838
rect 101254 278626 101260 278628
rect 98716 278566 101260 278626
rect 101254 278564 101260 278566
rect 101324 278564 101330 278628
rect 255405 278490 255471 278493
rect 253460 278488 255471 278490
rect 253460 278432 255410 278488
rect 255466 278432 255471 278488
rect 253460 278430 255471 278432
rect 255405 278427 255471 278430
rect 67541 278084 67607 278085
rect 67541 278082 67588 278084
rect 67460 278080 67588 278082
rect 67652 278082 67658 278084
rect 191465 278082 191531 278085
rect 256877 278082 256943 278085
rect 67460 278024 67546 278080
rect 67460 278022 67588 278024
rect 67541 278020 67588 278022
rect 67652 278022 68908 278082
rect 191465 278080 193660 278082
rect 191465 278024 191470 278080
rect 191526 278024 193660 278080
rect 191465 278022 193660 278024
rect 253460 278080 256943 278082
rect 253460 278024 256882 278080
rect 256938 278024 256943 278080
rect 253460 278022 256943 278024
rect 67652 278020 67658 278022
rect 67541 278019 67607 278020
rect 191465 278019 191531 278022
rect 256877 278019 256943 278022
rect 100753 277810 100819 277813
rect 98716 277808 100819 277810
rect 98716 277752 100758 277808
rect 100814 277752 100819 277808
rect 98716 277750 100819 277752
rect 100753 277747 100819 277750
rect 255497 277674 255563 277677
rect 253460 277672 255563 277674
rect 253460 277616 255502 277672
rect 255558 277616 255563 277672
rect 253460 277614 255563 277616
rect 255497 277611 255563 277614
rect 67817 277266 67883 277269
rect 255497 277266 255563 277269
rect 67817 277264 68908 277266
rect 67817 277208 67822 277264
rect 67878 277208 68908 277264
rect 67817 277206 68908 277208
rect 253460 277264 255563 277266
rect 253460 277208 255502 277264
rect 255558 277208 255563 277264
rect 253460 277206 255563 277208
rect 67817 277203 67883 277206
rect 255497 277203 255563 277206
rect 262305 277130 262371 277133
rect 253430 277128 262371 277130
rect 253430 277072 262310 277128
rect 262366 277072 262371 277128
rect 253430 277070 262371 277072
rect 101029 276994 101095 276997
rect 98716 276992 101095 276994
rect 98716 276936 101034 276992
rect 101090 276936 101095 276992
rect 98716 276934 101095 276936
rect 101029 276931 101095 276934
rect 190637 276994 190703 276997
rect 190637 276992 193660 276994
rect 190637 276936 190642 276992
rect 190698 276936 193660 276992
rect 190637 276934 193660 276936
rect 190637 276931 190703 276934
rect 253430 276828 253490 277070
rect 262305 277067 262371 277070
rect 66897 276450 66963 276453
rect 255405 276450 255471 276453
rect 66897 276448 68908 276450
rect 66897 276392 66902 276448
rect 66958 276392 68908 276448
rect 66897 276390 68908 276392
rect 253460 276448 255471 276450
rect 253460 276392 255410 276448
rect 255466 276392 255471 276448
rect 253460 276390 255471 276392
rect 66897 276387 66963 276390
rect 255405 276387 255471 276390
rect 100845 276178 100911 276181
rect 98716 276176 100911 276178
rect 98716 276120 100850 276176
rect 100906 276120 100911 276176
rect 98716 276118 100911 276120
rect 100845 276115 100911 276118
rect 273253 276042 273319 276045
rect 276013 276042 276079 276045
rect 253460 276040 276079 276042
rect 253460 275984 273258 276040
rect 273314 275984 276018 276040
rect 276074 275984 276079 276040
rect 253460 275982 276079 275984
rect 273253 275979 273319 275982
rect 276013 275979 276079 275982
rect 191557 275906 191623 275909
rect 191557 275904 193660 275906
rect 191557 275848 191562 275904
rect 191618 275848 193660 275904
rect 191557 275846 193660 275848
rect 191557 275843 191623 275846
rect 68878 275090 68938 275604
rect 255497 275498 255563 275501
rect 253460 275496 255563 275498
rect 253460 275440 255502 275496
rect 255558 275440 255563 275496
rect 253460 275438 255563 275440
rect 255497 275435 255563 275438
rect 100937 275362 101003 275365
rect 98716 275360 101003 275362
rect 98716 275304 100942 275360
rect 100998 275304 101003 275360
rect 98716 275302 101003 275304
rect 100937 275299 101003 275302
rect 193806 275300 193812 275364
rect 193876 275300 193882 275364
rect 101029 275226 101095 275229
rect 103830 275226 103836 275228
rect 101029 275224 103836 275226
rect 101029 275168 101034 275224
rect 101090 275168 103836 275224
rect 101029 275166 103836 275168
rect 101029 275163 101095 275166
rect 103830 275164 103836 275166
rect 103900 275226 103906 275228
rect 117497 275226 117563 275229
rect 103900 275224 117563 275226
rect 103900 275168 117502 275224
rect 117558 275168 117563 275224
rect 103900 275166 117563 275168
rect 103900 275164 103906 275166
rect 117497 275163 117563 275166
rect 64830 275030 68938 275090
rect 57789 274818 57855 274821
rect 64830 274818 64890 275030
rect 57789 274816 64890 274818
rect 57789 274760 57794 274816
rect 57850 274760 64890 274816
rect 57789 274758 64890 274760
rect 66437 274818 66503 274821
rect 66437 274816 68908 274818
rect 66437 274760 66442 274816
rect 66498 274760 68908 274816
rect 66437 274758 68908 274760
rect 57789 274755 57855 274758
rect 66437 274755 66503 274758
rect 185342 274620 185348 274684
rect 185412 274682 185418 274684
rect 193814 274682 193874 275300
rect 255405 275090 255471 275093
rect 253460 275088 255471 275090
rect 253460 275032 255410 275088
rect 255466 275032 255471 275088
rect 253460 275030 255471 275032
rect 255405 275027 255471 275030
rect 270493 274682 270559 274685
rect 185412 274622 193874 274682
rect 253460 274680 270559 274682
rect 253460 274624 270498 274680
rect 270554 274624 270559 274680
rect 253460 274622 270559 274624
rect 185412 274620 185418 274622
rect 270493 274619 270559 274622
rect 100845 274546 100911 274549
rect 98716 274544 100911 274546
rect 98716 274488 100850 274544
rect 100906 274488 100911 274544
rect 98716 274486 100911 274488
rect 100845 274483 100911 274486
rect 255405 274274 255471 274277
rect 253460 274272 255471 274274
rect 253460 274216 255410 274272
rect 255466 274216 255471 274272
rect 253460 274214 255471 274216
rect 255405 274211 255471 274214
rect 68878 273458 68938 273972
rect 255497 273866 255563 273869
rect 270677 273866 270743 273869
rect 282913 273866 282979 273869
rect 253460 273864 255563 273866
rect 253460 273808 255502 273864
rect 255558 273808 255563 273864
rect 253460 273806 255563 273808
rect 255497 273803 255563 273806
rect 258030 273864 282979 273866
rect 258030 273808 270682 273864
rect 270738 273808 282918 273864
rect 282974 273808 282979 273864
rect 258030 273806 282979 273808
rect 101397 273730 101463 273733
rect 98716 273728 101463 273730
rect 98716 273672 101402 273728
rect 101458 273672 101463 273728
rect 98716 273670 101463 273672
rect 101397 273667 101463 273670
rect 190821 273730 190887 273733
rect 190821 273728 193660 273730
rect 190821 273672 190826 273728
rect 190882 273672 193660 273728
rect 190821 273670 193660 273672
rect 190821 273667 190887 273670
rect 258030 273594 258090 273806
rect 270677 273803 270743 273806
rect 282913 273803 282979 273806
rect 64830 273398 68938 273458
rect 253430 273534 258090 273594
rect 253430 273428 253490 273534
rect 61101 273322 61167 273325
rect 61929 273322 61995 273325
rect 64830 273322 64890 273398
rect 61101 273320 64890 273322
rect 61101 273264 61106 273320
rect 61162 273264 61934 273320
rect 61990 273264 64890 273320
rect 61101 273262 64890 273264
rect 61101 273259 61167 273262
rect 61929 273259 61995 273262
rect 66805 273186 66871 273189
rect 255405 273186 255471 273189
rect 272057 273186 272123 273189
rect 66805 273184 68908 273186
rect 66805 273128 66810 273184
rect 66866 273128 68908 273184
rect 66805 273126 68908 273128
rect 255405 273184 272123 273186
rect 255405 273128 255410 273184
rect 255466 273128 272062 273184
rect 272118 273128 272123 273184
rect 255405 273126 272123 273128
rect 66805 273123 66871 273126
rect 255405 273123 255471 273126
rect 272057 273123 272123 273126
rect 100845 272914 100911 272917
rect 98716 272912 100911 272914
rect 98716 272856 100850 272912
rect 100906 272856 100911 272912
rect 98716 272854 100911 272856
rect 100845 272851 100911 272854
rect 253430 272778 253490 272884
rect 253430 272718 258090 272778
rect 191557 272642 191623 272645
rect 191557 272640 193660 272642
rect 191557 272584 191562 272640
rect 191618 272584 193660 272640
rect 191557 272582 193660 272584
rect 191557 272579 191623 272582
rect 104709 272506 104775 272509
rect 138841 272506 138907 272509
rect 98686 272504 138907 272506
rect 98686 272448 104714 272504
rect 104770 272448 138846 272504
rect 138902 272448 138907 272504
rect 98686 272446 138907 272448
rect 66069 272370 66135 272373
rect 66621 272370 66687 272373
rect 66069 272368 68908 272370
rect 66069 272312 66074 272368
rect 66130 272312 66626 272368
rect 66682 272312 68908 272368
rect 66069 272310 68908 272312
rect 66069 272307 66135 272310
rect 66621 272307 66687 272310
rect 98686 272068 98746 272446
rect 104709 272443 104775 272446
rect 138841 272443 138907 272446
rect 144177 272506 144243 272509
rect 155166 272506 155172 272508
rect 144177 272504 155172 272506
rect 144177 272448 144182 272504
rect 144238 272448 155172 272504
rect 144177 272446 155172 272448
rect 144177 272443 144243 272446
rect 155166 272444 155172 272446
rect 155236 272444 155242 272508
rect 255497 272506 255563 272509
rect 253460 272504 255563 272506
rect 253460 272448 255502 272504
rect 255558 272448 255563 272504
rect 253460 272446 255563 272448
rect 258030 272506 258090 272718
rect 269389 272506 269455 272509
rect 258030 272504 269455 272506
rect 258030 272448 269394 272504
rect 269450 272448 269455 272504
rect 258030 272446 269455 272448
rect 255497 272443 255563 272446
rect 269389 272443 269455 272446
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 255405 272098 255471 272101
rect 253460 272096 255471 272098
rect 253460 272040 255410 272096
rect 255466 272040 255471 272096
rect 583520 272084 584960 272174
rect 253460 272038 255471 272040
rect 255405 272035 255471 272038
rect 59077 271962 59143 271965
rect 66805 271962 66871 271965
rect 59077 271960 66871 271962
rect 59077 271904 59082 271960
rect 59138 271904 66810 271960
rect 66866 271904 66871 271960
rect 59077 271902 66871 271904
rect 59077 271899 59143 271902
rect 66805 271899 66871 271902
rect 255497 271826 255563 271829
rect 276105 271826 276171 271829
rect 277669 271826 277735 271829
rect 255497 271824 277735 271826
rect 255497 271768 255502 271824
rect 255558 271768 276110 271824
rect 276166 271768 277674 271824
rect 277730 271768 277735 271824
rect 255497 271766 277735 271768
rect 255497 271763 255563 271766
rect 276105 271763 276171 271766
rect 277669 271763 277735 271766
rect 255313 271690 255379 271693
rect 253460 271688 255379 271690
rect 253460 271632 255318 271688
rect 255374 271632 255379 271688
rect 253460 271630 255379 271632
rect 255313 271627 255379 271630
rect 191557 271554 191623 271557
rect 191557 271552 193660 271554
rect 68878 271010 68938 271524
rect 191557 271496 191562 271552
rect 191618 271496 193660 271552
rect 191557 271494 193660 271496
rect 191557 271491 191623 271494
rect 99465 271282 99531 271285
rect 101489 271282 101555 271285
rect 255405 271282 255471 271285
rect 98716 271280 101555 271282
rect 98716 271224 99470 271280
rect 99526 271224 101494 271280
rect 101550 271224 101555 271280
rect 98716 271222 101555 271224
rect 253460 271280 255471 271282
rect 253460 271224 255410 271280
rect 255466 271224 255471 271280
rect 253460 271222 255471 271224
rect 99465 271219 99531 271222
rect 101489 271219 101555 271222
rect 255405 271219 255471 271222
rect 255773 271146 255839 271149
rect 270769 271146 270835 271149
rect 280153 271146 280219 271149
rect 255773 271144 280219 271146
rect 255773 271088 255778 271144
rect 255834 271088 270774 271144
rect 270830 271088 280158 271144
rect 280214 271088 280219 271144
rect 255773 271086 280219 271088
rect 255773 271083 255839 271086
rect 270769 271083 270835 271086
rect 280153 271083 280219 271086
rect 64830 270950 68938 271010
rect 61837 270738 61903 270741
rect 64830 270738 64890 270950
rect 255497 270874 255563 270877
rect 253460 270872 255563 270874
rect 253460 270816 255502 270872
rect 255558 270816 255563 270872
rect 253460 270814 255563 270816
rect 255497 270811 255563 270814
rect 61837 270736 64890 270738
rect 61837 270680 61842 270736
rect 61898 270680 64890 270736
rect 61837 270678 64890 270680
rect 66529 270738 66595 270741
rect 66529 270736 68908 270738
rect 66529 270680 66534 270736
rect 66590 270680 68908 270736
rect 66529 270678 68908 270680
rect 61837 270675 61903 270678
rect 66529 270675 66595 270678
rect 255313 270602 255379 270605
rect 262397 270602 262463 270605
rect 255313 270600 262463 270602
rect 255313 270544 255318 270600
rect 255374 270544 262402 270600
rect 262458 270544 262463 270600
rect 255313 270542 262463 270544
rect 255313 270539 255379 270542
rect 262397 270539 262463 270542
rect 100845 270466 100911 270469
rect 98716 270464 100911 270466
rect 98716 270408 100850 270464
rect 100906 270408 100911 270464
rect 98716 270406 100911 270408
rect 100845 270403 100911 270406
rect 173249 270466 173315 270469
rect 176510 270466 176516 270468
rect 173249 270464 176516 270466
rect 173249 270408 173254 270464
rect 173310 270408 176516 270464
rect 173249 270406 176516 270408
rect 173249 270403 173315 270406
rect 176510 270404 176516 270406
rect 176580 270466 176586 270468
rect 189073 270466 189139 270469
rect 176580 270464 189139 270466
rect 176580 270408 189078 270464
rect 189134 270408 189139 270464
rect 176580 270406 189139 270408
rect 176580 270404 176586 270406
rect 189073 270403 189139 270406
rect 191465 270466 191531 270469
rect 262213 270466 262279 270469
rect 263726 270466 263732 270468
rect 191465 270464 193660 270466
rect 191465 270408 191470 270464
rect 191526 270408 193660 270464
rect 262213 270464 263732 270466
rect 191465 270406 193660 270408
rect 191465 270403 191531 270406
rect 253430 270194 253490 270436
rect 262213 270408 262218 270464
rect 262274 270408 263732 270464
rect 262213 270406 263732 270408
rect 262213 270403 262279 270406
rect 263726 270404 263732 270406
rect 263796 270404 263802 270468
rect 262213 270194 262279 270197
rect 253430 270192 262279 270194
rect 253430 270136 262218 270192
rect 262274 270136 262279 270192
rect 253430 270134 262279 270136
rect 262213 270131 262279 270134
rect 66805 269922 66871 269925
rect 255405 269922 255471 269925
rect 66805 269920 68908 269922
rect 66805 269864 66810 269920
rect 66866 269864 68908 269920
rect 66805 269862 68908 269864
rect 253460 269920 255471 269922
rect 253460 269864 255410 269920
rect 255466 269864 255471 269920
rect 253460 269862 255471 269864
rect 66805 269859 66871 269862
rect 255405 269859 255471 269862
rect 165470 269724 165476 269788
rect 165540 269786 165546 269788
rect 178677 269786 178743 269789
rect 165540 269784 178743 269786
rect 165540 269728 178682 269784
rect 178738 269728 178743 269784
rect 165540 269726 178743 269728
rect 165540 269724 165546 269726
rect 178677 269723 178743 269726
rect 98686 269242 98746 269620
rect 191557 269378 191623 269381
rect 253430 269378 253490 269484
rect 266537 269378 266603 269381
rect 273621 269378 273687 269381
rect 191557 269376 193660 269378
rect 191557 269320 191562 269376
rect 191618 269320 193660 269376
rect 191557 269318 193660 269320
rect 253430 269376 273687 269378
rect 253430 269320 266542 269376
rect 266598 269320 273626 269376
rect 273682 269320 273687 269376
rect 253430 269318 273687 269320
rect 191557 269315 191623 269318
rect 266537 269315 266603 269318
rect 273621 269315 273687 269318
rect 108297 269242 108363 269245
rect 98686 269240 108363 269242
rect 98686 269184 108302 269240
rect 108358 269184 108363 269240
rect 98686 269182 108363 269184
rect 108297 269179 108363 269182
rect 189073 269242 189139 269245
rect 191465 269242 191531 269245
rect 189073 269240 191531 269242
rect 189073 269184 189078 269240
rect 189134 269184 191470 269240
rect 191526 269184 191531 269240
rect 189073 269182 191531 269184
rect 189073 269179 189139 269182
rect 191465 269179 191531 269182
rect 255497 269106 255563 269109
rect 253460 269104 255563 269106
rect 65885 268562 65951 268565
rect 68878 268562 68938 269076
rect 253460 269048 255502 269104
rect 255558 269048 255563 269104
rect 253460 269046 255563 269048
rect 255497 269043 255563 269046
rect 64830 268560 68938 268562
rect 64830 268504 65890 268560
rect 65946 268504 68938 268560
rect 64830 268502 68938 268504
rect 49601 268426 49667 268429
rect 64830 268426 64890 268502
rect 65885 268499 65951 268502
rect 49601 268424 64890 268426
rect 49601 268368 49606 268424
rect 49662 268368 64890 268424
rect 49601 268366 64890 268368
rect 49601 268363 49667 268366
rect 66805 268290 66871 268293
rect 98686 268290 98746 268804
rect 253430 268562 253490 268668
rect 291377 268562 291443 268565
rect 253430 268560 291443 268562
rect 253430 268504 291382 268560
rect 291438 268504 291443 268560
rect 253430 268502 291443 268504
rect 291377 268499 291443 268502
rect 191557 268290 191623 268293
rect 255773 268290 255839 268293
rect 66805 268288 68908 268290
rect 66805 268232 66810 268288
rect 66866 268232 68908 268288
rect 66805 268230 68908 268232
rect 98686 268230 103530 268290
rect 66805 268227 66871 268230
rect 100845 268018 100911 268021
rect 98716 268016 100911 268018
rect 98716 267960 100850 268016
rect 100906 267960 100911 268016
rect 98716 267958 100911 267960
rect 100845 267955 100911 267958
rect 103470 267882 103530 268230
rect 191557 268288 193660 268290
rect 191557 268232 191562 268288
rect 191618 268232 193660 268288
rect 191557 268230 193660 268232
rect 253460 268288 255839 268290
rect 253460 268232 255778 268288
rect 255834 268232 255839 268288
rect 253460 268230 255839 268232
rect 191557 268227 191623 268230
rect 255773 268227 255839 268230
rect 115289 267882 115355 267885
rect 255405 267882 255471 267885
rect 103470 267880 115355 267882
rect 103470 267824 115294 267880
rect 115350 267824 115355 267880
rect 103470 267822 115355 267824
rect 253460 267880 255471 267882
rect 253460 267824 255410 267880
rect 255466 267824 255471 267880
rect 253460 267822 255471 267824
rect 115289 267819 115355 267822
rect 255405 267819 255471 267822
rect 255405 267474 255471 267477
rect 253460 267472 255471 267474
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 68878 266930 68938 267444
rect 253460 267416 255410 267472
rect 255466 267416 255471 267472
rect 253460 267414 255471 267416
rect 255405 267411 255471 267414
rect 98686 267066 98746 267172
rect 106089 267066 106155 267069
rect 98686 267064 106155 267066
rect 98686 267008 106094 267064
rect 106150 267008 106155 267064
rect 98686 267006 106155 267008
rect 106089 267003 106155 267006
rect 64830 266870 68938 266930
rect 58341 266522 58407 266525
rect 59169 266522 59235 266525
rect 64830 266522 64890 266870
rect 65977 266658 66043 266661
rect 65977 266656 68908 266658
rect 65977 266600 65982 266656
rect 66038 266600 68908 266656
rect 65977 266598 68908 266600
rect 65977 266595 66043 266598
rect 58341 266520 64890 266522
rect 58341 266464 58346 266520
rect 58402 266464 59174 266520
rect 59230 266464 64890 266520
rect 58341 266462 64890 266464
rect 58341 266459 58407 266462
rect 59169 266459 59235 266462
rect 101029 266386 101095 266389
rect 98716 266384 101095 266386
rect 98716 266328 101034 266384
rect 101090 266328 101095 266384
rect 98716 266326 101095 266328
rect 101029 266323 101095 266326
rect 106089 266386 106155 266389
rect 108297 266386 108363 266389
rect 106089 266384 108363 266386
rect 106089 266328 106094 266384
rect 106150 266328 108302 266384
rect 108358 266328 108363 266384
rect 106089 266326 108363 266328
rect 106089 266323 106155 266326
rect 108297 266323 108363 266326
rect 158621 266386 158687 266389
rect 162853 266386 162919 266389
rect 193630 266386 193690 267172
rect 260966 267004 260972 267068
rect 261036 267066 261042 267068
rect 288382 267066 288388 267068
rect 261036 267006 288388 267066
rect 261036 267004 261042 267006
rect 288382 267004 288388 267006
rect 288452 267004 288458 267068
rect 256877 266930 256943 266933
rect 253460 266928 256943 266930
rect 253460 266872 256882 266928
rect 256938 266872 256943 266928
rect 253460 266870 256943 266872
rect 256877 266867 256943 266870
rect 259637 266522 259703 266525
rect 253460 266520 259703 266522
rect 253460 266464 259642 266520
rect 259698 266464 259703 266520
rect 253460 266462 259703 266464
rect 259637 266459 259703 266462
rect 158621 266384 193690 266386
rect 158621 266328 158626 266384
rect 158682 266328 162858 266384
rect 162914 266328 193690 266384
rect 158621 266326 193690 266328
rect 158621 266323 158687 266326
rect 162853 266323 162919 266326
rect 191649 266114 191715 266117
rect 255313 266114 255379 266117
rect 191649 266112 193660 266114
rect 191649 266056 191654 266112
rect 191710 266056 193660 266112
rect 252908 266112 255379 266114
rect 252908 266084 255318 266112
rect 191649 266054 193660 266056
rect 252878 266056 255318 266084
rect 255374 266056 255379 266112
rect 252878 266054 255379 266056
rect 191649 266051 191715 266054
rect 252878 265980 252938 266054
rect 255313 266051 255379 266054
rect 252870 265916 252876 265980
rect 252940 265916 252946 265980
rect 68878 265298 68938 265812
rect 255405 265706 255471 265709
rect 253460 265704 255471 265706
rect 253460 265648 255410 265704
rect 255466 265648 255471 265704
rect 253460 265646 255471 265648
rect 255405 265643 255471 265646
rect 100845 265570 100911 265573
rect 98716 265568 100911 265570
rect 98716 265512 100850 265568
rect 100906 265512 100911 265568
rect 98716 265510 100911 265512
rect 100845 265507 100911 265510
rect 262438 265508 262444 265572
rect 262508 265570 262514 265572
rect 274817 265570 274883 265573
rect 262508 265568 274883 265570
rect 262508 265512 274822 265568
rect 274878 265512 274883 265568
rect 262508 265510 274883 265512
rect 262508 265508 262514 265510
rect 274817 265507 274883 265510
rect 64830 265238 68938 265298
rect 50797 265026 50863 265029
rect 57881 265026 57947 265029
rect 64830 265026 64890 265238
rect 253430 265162 253490 265268
rect 262438 265162 262444 265164
rect 253430 265102 262444 265162
rect 262438 265100 262444 265102
rect 262508 265100 262514 265164
rect 50797 265024 64890 265026
rect 50797 264968 50802 265024
rect 50858 264968 57886 265024
rect 57942 264968 64890 265024
rect 50797 264966 64890 264968
rect 66805 265026 66871 265029
rect 190637 265026 190703 265029
rect 66805 265024 68908 265026
rect 66805 264968 66810 265024
rect 66866 264968 68908 265024
rect 66805 264966 68908 264968
rect 190637 265024 193660 265026
rect 190637 264968 190642 265024
rect 190698 264968 193660 265024
rect 190637 264966 193660 264968
rect 50797 264963 50863 264966
rect 57881 264963 57947 264966
rect 66805 264963 66871 264966
rect 190637 264963 190703 264966
rect 100937 264754 101003 264757
rect 98716 264752 101003 264754
rect 98716 264696 100942 264752
rect 100998 264696 101003 264752
rect 98716 264694 101003 264696
rect 100937 264691 101003 264694
rect 253430 264618 253490 264860
rect 253430 264558 258090 264618
rect 255497 264346 255563 264349
rect 253460 264344 255563 264346
rect 253460 264288 255502 264344
rect 255558 264288 255563 264344
rect 253460 264286 255563 264288
rect 255497 264283 255563 264286
rect 66621 264210 66687 264213
rect 258030 264210 258090 264558
rect 288525 264210 288591 264213
rect 66621 264208 68908 264210
rect 66621 264152 66626 264208
rect 66682 264152 68908 264208
rect 66621 264150 68908 264152
rect 258030 264208 288591 264210
rect 258030 264152 288530 264208
rect 288586 264152 288591 264208
rect 258030 264150 288591 264152
rect 66621 264147 66687 264150
rect 288525 264147 288591 264150
rect 192017 263938 192083 263941
rect 255405 263938 255471 263941
rect 192017 263936 193660 263938
rect 98686 263666 98746 263908
rect 192017 263880 192022 263936
rect 192078 263880 193660 263936
rect 192017 263878 193660 263880
rect 253460 263936 255471 263938
rect 253460 263880 255410 263936
rect 255466 263880 255471 263936
rect 253460 263878 255471 263880
rect 192017 263875 192083 263878
rect 255405 263875 255471 263878
rect 109769 263666 109835 263669
rect 98686 263664 109835 263666
rect 98686 263608 109774 263664
rect 109830 263608 109835 263664
rect 98686 263606 109835 263608
rect 109769 263603 109835 263606
rect 260741 263530 260807 263533
rect 253460 263528 260807 263530
rect 253460 263472 260746 263528
rect 260802 263472 260807 263528
rect 253460 263470 260807 263472
rect 260741 263467 260807 263470
rect 285121 263530 285187 263533
rect 288709 263530 288775 263533
rect 285121 263528 288775 263530
rect 285121 263472 285126 263528
rect 285182 263472 288714 263528
rect 288770 263472 288775 263528
rect 285121 263470 288775 263472
rect 285121 263467 285187 263470
rect 288709 263467 288775 263470
rect 67081 263394 67147 263397
rect 67449 263394 67515 263397
rect 67081 263392 68908 263394
rect 67081 263336 67086 263392
rect 67142 263336 67454 263392
rect 67510 263336 68908 263392
rect 67081 263334 68908 263336
rect 67081 263331 67147 263334
rect 67449 263331 67515 263334
rect 100845 263122 100911 263125
rect 255497 263122 255563 263125
rect 98716 263120 100911 263122
rect 98716 263064 100850 263120
rect 100906 263064 100911 263120
rect 98716 263062 100911 263064
rect 253460 263120 255563 263122
rect 253460 263064 255502 263120
rect 255558 263064 255563 263120
rect 253460 263062 255563 263064
rect 100845 263059 100911 263062
rect 255497 263059 255563 263062
rect 191649 262850 191715 262853
rect 281574 262850 281580 262852
rect 191649 262848 193660 262850
rect 191649 262792 191654 262848
rect 191710 262792 193660 262848
rect 191649 262790 193660 262792
rect 253430 262790 281580 262850
rect 191649 262787 191715 262790
rect 253430 262684 253490 262790
rect 281574 262788 281580 262790
rect 281644 262850 281650 262852
rect 281717 262850 281783 262853
rect 281644 262848 281783 262850
rect 281644 262792 281722 262848
rect 281778 262792 281783 262848
rect 281644 262790 281783 262792
rect 281644 262788 281650 262790
rect 281717 262787 281783 262790
rect 263869 262716 263935 262717
rect 263869 262714 263916 262716
rect 263824 262712 263916 262714
rect 263824 262656 263874 262712
rect 263824 262654 263916 262656
rect 263869 262652 263916 262654
rect 263980 262652 263986 262716
rect 263869 262651 263935 262652
rect 66897 262578 66963 262581
rect 66897 262576 68908 262578
rect 66897 262520 66902 262576
rect 66958 262520 68908 262576
rect 66897 262518 68908 262520
rect 66897 262515 66963 262518
rect 268285 262442 268351 262445
rect 270718 262442 270724 262444
rect 268285 262440 270724 262442
rect 268285 262384 268290 262440
rect 268346 262384 270724 262440
rect 268285 262382 270724 262384
rect 268285 262379 268351 262382
rect 270718 262380 270724 262382
rect 270788 262380 270794 262444
rect 100017 262306 100083 262309
rect 101121 262306 101187 262309
rect 255405 262306 255471 262309
rect 98716 262304 101187 262306
rect 98716 262248 100022 262304
rect 100078 262248 101126 262304
rect 101182 262248 101187 262304
rect 98716 262246 101187 262248
rect 253460 262304 255471 262306
rect 253460 262248 255410 262304
rect 255466 262248 255471 262304
rect 253460 262246 255471 262248
rect 100017 262243 100083 262246
rect 101121 262243 101187 262246
rect 255405 262243 255471 262246
rect 261477 262306 261543 262309
rect 284477 262306 284543 262309
rect 285121 262306 285187 262309
rect 261477 262304 285187 262306
rect 261477 262248 261482 262304
rect 261538 262248 284482 262304
rect 284538 262248 285126 262304
rect 285182 262248 285187 262304
rect 261477 262246 285187 262248
rect 261477 262243 261543 262246
rect 284477 262243 284543 262246
rect 285121 262243 285187 262246
rect 273662 262108 273668 262172
rect 273732 262170 273738 262172
rect 278957 262170 279023 262173
rect 273732 262168 279023 262170
rect 273732 262112 278962 262168
rect 279018 262112 279023 262168
rect 273732 262110 279023 262112
rect 273732 262108 273738 262110
rect 278957 262107 279023 262110
rect 255405 261898 255471 261901
rect 253460 261896 255471 261898
rect 253460 261840 255410 261896
rect 255466 261840 255471 261896
rect 253460 261838 255471 261840
rect 255405 261835 255471 261838
rect 191649 261762 191715 261765
rect 191649 261760 193660 261762
rect 68878 261218 68938 261732
rect 191649 261704 191654 261760
rect 191710 261704 193660 261760
rect 191649 261702 193660 261704
rect 191649 261699 191715 261702
rect 100845 261490 100911 261493
rect 98716 261488 100911 261490
rect 98716 261432 100850 261488
rect 100906 261432 100911 261488
rect 98716 261430 100911 261432
rect 100845 261427 100911 261430
rect 101029 261490 101095 261493
rect 155401 261490 155467 261493
rect 101029 261488 155467 261490
rect 101029 261432 101034 261488
rect 101090 261432 155406 261488
rect 155462 261432 155467 261488
rect 101029 261430 155467 261432
rect 101029 261427 101095 261430
rect 155401 261427 155467 261430
rect 263542 261428 263548 261492
rect 263612 261490 263618 261492
rect 284334 261490 284340 261492
rect 263612 261430 284340 261490
rect 263612 261428 263618 261430
rect 284334 261428 284340 261430
rect 284404 261428 284410 261492
rect 64830 261158 68938 261218
rect 253430 261218 253490 261324
rect 273662 261218 273668 261220
rect 253430 261158 273668 261218
rect 60549 261082 60615 261085
rect 61745 261082 61811 261085
rect 64830 261082 64890 261158
rect 273662 261156 273668 261158
rect 273732 261156 273738 261220
rect 60549 261080 64890 261082
rect 60549 261024 60554 261080
rect 60610 261024 61750 261080
rect 61806 261024 64890 261080
rect 60549 261022 64890 261024
rect 255313 261082 255379 261085
rect 263542 261082 263548 261084
rect 255313 261080 263548 261082
rect 255313 261024 255318 261080
rect 255374 261024 263548 261080
rect 255313 261022 263548 261024
rect 60549 261019 60615 261022
rect 61745 261019 61811 261022
rect 255313 261019 255379 261022
rect 263542 261020 263548 261022
rect 263612 261020 263618 261084
rect 66253 260946 66319 260949
rect 255497 260946 255563 260949
rect 66253 260944 68908 260946
rect 66253 260888 66258 260944
rect 66314 260888 68908 260944
rect 66253 260886 68908 260888
rect 253460 260944 255563 260946
rect 253460 260888 255502 260944
rect 255558 260888 255563 260944
rect 253460 260886 255563 260888
rect 66253 260883 66319 260886
rect 255497 260883 255563 260886
rect 100845 260674 100911 260677
rect 98716 260672 100911 260674
rect 98716 260616 100850 260672
rect 100906 260616 100911 260672
rect 98716 260614 100911 260616
rect 100845 260611 100911 260614
rect 191373 260674 191439 260677
rect 191373 260672 193660 260674
rect 191373 260616 191378 260672
rect 191434 260616 193660 260672
rect 191373 260614 193660 260616
rect 191373 260611 191439 260614
rect 167637 260538 167703 260541
rect 168966 260538 168972 260540
rect 167637 260536 168972 260538
rect 167637 260480 167642 260536
rect 167698 260480 168972 260536
rect 167637 260478 168972 260480
rect 167637 260475 167703 260478
rect 168966 260476 168972 260478
rect 169036 260538 169042 260540
rect 169293 260538 169359 260541
rect 255405 260538 255471 260541
rect 169036 260536 169359 260538
rect 169036 260480 169298 260536
rect 169354 260480 169359 260536
rect 169036 260478 169359 260480
rect 253460 260536 255471 260538
rect 253460 260480 255410 260536
rect 255466 260480 255471 260536
rect 253460 260478 255471 260480
rect 169036 260476 169042 260478
rect 169293 260475 169359 260478
rect 255405 260475 255471 260478
rect 260741 260538 260807 260541
rect 260966 260538 260972 260540
rect 260741 260536 260972 260538
rect 260741 260480 260746 260536
rect 260802 260480 260972 260536
rect 260741 260478 260972 260480
rect 260741 260475 260807 260478
rect 260966 260476 260972 260478
rect 261036 260476 261042 260540
rect 265249 260266 265315 260269
rect 273294 260266 273300 260268
rect 265249 260264 273300 260266
rect 265249 260208 265254 260264
rect 265310 260208 273300 260264
rect 265249 260206 273300 260208
rect 265249 260203 265315 260206
rect 273294 260204 273300 260206
rect 273364 260204 273370 260268
rect 67725 260130 67791 260133
rect 67725 260128 68908 260130
rect 67725 260072 67730 260128
rect 67786 260072 68908 260128
rect 67725 260070 68908 260072
rect 67725 260067 67791 260070
rect 159950 260068 159956 260132
rect 160020 260130 160026 260132
rect 176653 260130 176719 260133
rect 295333 260130 295399 260133
rect 160020 260128 176719 260130
rect 160020 260072 176658 260128
rect 176714 260072 176719 260128
rect 267690 260128 295399 260130
rect 160020 260070 176719 260072
rect 160020 260068 160026 260070
rect 176653 260067 176719 260070
rect 253430 259994 253490 260100
rect 267690 260072 295338 260128
rect 295394 260072 295399 260128
rect 267690 260070 295399 260072
rect 263726 259994 263732 259996
rect 253430 259934 263732 259994
rect 263726 259932 263732 259934
rect 263796 259994 263802 259996
rect 267690 259994 267750 260070
rect 295333 260067 295399 260070
rect 263796 259934 267750 259994
rect 263796 259932 263802 259934
rect 101949 259858 102015 259861
rect 98716 259856 102015 259858
rect 98716 259800 101954 259856
rect 102010 259800 102015 259856
rect 98716 259798 102015 259800
rect 101949 259795 102015 259798
rect 255313 259722 255379 259725
rect 253460 259720 255379 259722
rect 253460 259664 255318 259720
rect 255374 259664 255379 259720
rect 253460 259662 255379 259664
rect 255313 259659 255379 259662
rect 191649 259586 191715 259589
rect 191649 259584 193660 259586
rect 191649 259528 191654 259584
rect 191710 259528 193660 259584
rect 191649 259526 193660 259528
rect 191649 259523 191715 259526
rect 271086 259388 271092 259452
rect 271156 259450 271162 259452
rect 276422 259450 276428 259452
rect 271156 259390 276428 259450
rect 271156 259388 271162 259390
rect 276422 259388 276428 259390
rect 276492 259388 276498 259452
rect 68185 258770 68251 258773
rect 68878 258770 68938 259284
rect 253430 259178 253490 259284
rect 265157 259178 265223 259181
rect 253430 259176 265223 259178
rect 253430 259120 265162 259176
rect 265218 259120 265223 259176
rect 253430 259118 265223 259120
rect 265157 259115 265223 259118
rect 99373 259042 99439 259045
rect 98716 259040 99439 259042
rect 98716 258984 99378 259040
rect 99434 258984 99439 259040
rect 98716 258982 99439 258984
rect 99373 258979 99439 258982
rect 258390 258906 258396 258908
rect 253460 258846 258396 258906
rect 258390 258844 258396 258846
rect 258460 258844 258466 258908
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 98361 258770 98427 258773
rect 68185 258768 68938 258770
rect 68185 258712 68190 258768
rect 68246 258712 68938 258768
rect 68185 258710 68938 258712
rect 98318 258768 98427 258770
rect 98318 258712 98366 258768
rect 98422 258712 98427 258768
rect 583520 258756 584960 258846
rect 68185 258707 68251 258710
rect 98318 258707 98427 258712
rect 66805 258498 66871 258501
rect 66805 258496 68908 258498
rect 66805 258440 66810 258496
rect 66866 258440 68908 258496
rect 66805 258438 68908 258440
rect 66805 258435 66871 258438
rect 98318 258196 98378 258707
rect 190453 258090 190519 258093
rect 190453 258088 190562 258090
rect 190453 258032 190458 258088
rect 190514 258032 190562 258088
rect 190453 258027 190562 258032
rect 144821 257954 144887 257957
rect 171133 257954 171199 257957
rect 144821 257952 171199 257954
rect 144821 257896 144826 257952
rect 144882 257896 171138 257952
rect 171194 257896 171199 257952
rect 144821 257894 171199 257896
rect 190502 257954 190562 258027
rect 193630 257954 193690 258468
rect 255405 258362 255471 258365
rect 271086 258362 271092 258364
rect 253460 258360 255471 258362
rect 253460 258304 255410 258360
rect 255466 258304 255471 258360
rect 253460 258302 255471 258304
rect 255405 258299 255471 258302
rect 256374 258302 271092 258362
rect 256374 257954 256434 258302
rect 271086 258300 271092 258302
rect 271156 258300 271162 258364
rect 258073 258226 258139 258229
rect 285622 258226 285628 258228
rect 258073 258224 285628 258226
rect 258073 258168 258078 258224
rect 258134 258168 285628 258224
rect 258073 258166 285628 258168
rect 258073 258163 258139 258166
rect 274774 257957 274834 258166
rect 285622 258164 285628 258166
rect 285692 258164 285698 258228
rect 190502 257894 193690 257954
rect 253460 257894 256434 257954
rect 274725 257952 274834 257957
rect 274725 257896 274730 257952
rect 274786 257896 274834 257952
rect 274725 257894 274834 257896
rect 144821 257891 144887 257894
rect 171133 257891 171199 257894
rect 274725 257891 274791 257894
rect 66253 257682 66319 257685
rect 66253 257680 68908 257682
rect 66253 257624 66258 257680
rect 66314 257624 68908 257680
rect 66253 257622 68908 257624
rect 66253 257619 66319 257622
rect 255313 257546 255379 257549
rect 253460 257544 255379 257546
rect 253460 257488 255318 257544
rect 255374 257488 255379 257544
rect 253460 257486 255379 257488
rect 255313 257483 255379 257486
rect 101397 257410 101463 257413
rect 98716 257408 101463 257410
rect 98716 257352 101402 257408
rect 101458 257352 101463 257408
rect 98716 257350 101463 257352
rect 101397 257347 101463 257350
rect 190637 257410 190703 257413
rect 190637 257408 193660 257410
rect 190637 257352 190642 257408
rect 190698 257352 193660 257408
rect 190637 257350 193660 257352
rect 190637 257347 190703 257350
rect 178677 257274 178743 257277
rect 185577 257274 185643 257277
rect 262438 257274 262444 257276
rect 178677 257272 185643 257274
rect 178677 257216 178682 257272
rect 178738 257216 185582 257272
rect 185638 257216 185643 257272
rect 178677 257214 185643 257216
rect 178677 257211 178743 257214
rect 185577 257211 185643 257214
rect 258030 257214 262444 257274
rect 255405 257138 255471 257141
rect 253460 257136 255471 257138
rect 253460 257080 255410 257136
rect 255466 257080 255471 257136
rect 253460 257078 255471 257080
rect 255405 257075 255471 257078
rect 67357 256866 67423 256869
rect 67357 256864 68908 256866
rect 67357 256808 67362 256864
rect 67418 256808 68908 256864
rect 67357 256806 68908 256808
rect 67357 256803 67423 256806
rect 258030 256730 258090 257214
rect 262438 257212 262444 257214
rect 262508 257274 262514 257276
rect 285857 257274 285923 257277
rect 262508 257272 285923 257274
rect 262508 257216 285862 257272
rect 285918 257216 285923 257272
rect 262508 257214 285923 257216
rect 262508 257212 262514 257214
rect 285857 257211 285923 257214
rect 253460 256670 258090 256730
rect 100937 256594 101003 256597
rect 98716 256592 101003 256594
rect 98716 256536 100942 256592
rect 100998 256536 101003 256592
rect 98716 256534 101003 256536
rect 100937 256531 101003 256534
rect 191649 256322 191715 256325
rect 255497 256322 255563 256325
rect 191649 256320 193660 256322
rect 191649 256264 191654 256320
rect 191710 256264 193660 256320
rect 191649 256262 193660 256264
rect 253460 256320 255563 256322
rect 253460 256264 255502 256320
rect 255558 256264 255563 256320
rect 253460 256262 255563 256264
rect 191649 256259 191715 256262
rect 255497 256259 255563 256262
rect 68878 255506 68938 256020
rect 173934 255988 173940 256052
rect 174004 256050 174010 256052
rect 175181 256050 175247 256053
rect 174004 256048 175247 256050
rect 174004 255992 175186 256048
rect 175242 255992 175247 256048
rect 174004 255990 175247 255992
rect 174004 255988 174010 255990
rect 175181 255987 175247 255990
rect 100702 255778 100708 255780
rect 98716 255718 100708 255778
rect 100702 255716 100708 255718
rect 100772 255778 100778 255780
rect 100845 255778 100911 255781
rect 258073 255778 258139 255781
rect 100772 255776 100911 255778
rect 100772 255720 100850 255776
rect 100906 255720 100911 255776
rect 100772 255718 100911 255720
rect 253460 255776 258139 255778
rect 253460 255720 258078 255776
rect 258134 255720 258139 255776
rect 253460 255718 258139 255720
rect 100772 255716 100778 255718
rect 100845 255715 100911 255718
rect 258073 255715 258139 255718
rect 64830 255446 68938 255506
rect 63401 255370 63467 255373
rect 64638 255370 64644 255372
rect 63401 255368 64644 255370
rect 63401 255312 63406 255368
rect 63462 255312 64644 255368
rect 63401 255310 64644 255312
rect 63401 255307 63467 255310
rect 64638 255308 64644 255310
rect 64708 255370 64714 255372
rect 64830 255370 64890 255446
rect 255405 255370 255471 255373
rect 64708 255310 64890 255370
rect 253460 255368 255471 255370
rect 253460 255312 255410 255368
rect 255466 255312 255471 255368
rect 253460 255310 255471 255312
rect 64708 255308 64714 255310
rect 255405 255307 255471 255310
rect 66805 255234 66871 255237
rect 191005 255234 191071 255237
rect 66805 255232 68908 255234
rect 66805 255176 66810 255232
rect 66866 255176 68908 255232
rect 66805 255174 68908 255176
rect 191005 255232 193660 255234
rect 191005 255176 191010 255232
rect 191066 255176 193660 255232
rect 191005 255174 193660 255176
rect 66805 255171 66871 255174
rect 191005 255171 191071 255174
rect 100845 254962 100911 254965
rect 255497 254962 255563 254965
rect 98716 254960 100911 254962
rect 98716 254904 100850 254960
rect 100906 254904 100911 254960
rect 98716 254902 100911 254904
rect 253460 254960 255563 254962
rect 253460 254904 255502 254960
rect 255558 254904 255563 254960
rect 253460 254902 255563 254904
rect 100845 254899 100911 254902
rect 255497 254899 255563 254902
rect 255405 254554 255471 254557
rect 253460 254552 255471 254554
rect 253460 254496 255410 254552
rect 255466 254496 255471 254552
rect 253460 254494 255471 254496
rect 255405 254491 255471 254494
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 56317 254146 56383 254149
rect 56501 254146 56567 254149
rect 68878 254146 68938 254388
rect 56317 254144 68938 254146
rect 56317 254088 56322 254144
rect 56378 254088 56506 254144
rect 56562 254088 68938 254144
rect 181437 254146 181503 254149
rect 188838 254146 188844 254148
rect 181437 254144 188844 254146
rect 56317 254086 68938 254088
rect 56317 254083 56383 254086
rect 56501 254083 56567 254086
rect 98686 254010 98746 254116
rect 181437 254088 181442 254144
rect 181498 254088 188844 254144
rect 181437 254086 188844 254088
rect 181437 254083 181503 254086
rect 188838 254084 188844 254086
rect 188908 254146 188914 254148
rect 188908 254086 193660 254146
rect 188908 254084 188914 254086
rect 112621 254010 112687 254013
rect 98686 254008 112687 254010
rect 98686 253952 112626 254008
rect 112682 253952 112687 254008
rect 98686 253950 112687 253952
rect 112621 253947 112687 253950
rect 175774 253948 175780 254012
rect 175844 254010 175850 254012
rect 177757 254010 177823 254013
rect 175844 254008 177823 254010
rect 175844 253952 177762 254008
rect 177818 253952 177823 254008
rect 175844 253950 177823 253952
rect 175844 253948 175850 253950
rect 177757 253947 177823 253950
rect 178534 253948 178540 254012
rect 178604 254010 178610 254012
rect 180149 254010 180215 254013
rect 178604 254008 180215 254010
rect 178604 253952 180154 254008
rect 180210 253952 180215 254008
rect 178604 253950 180215 253952
rect 253430 254010 253490 254116
rect 254025 254010 254091 254013
rect 261109 254010 261175 254013
rect 253430 254008 261175 254010
rect 253430 253952 254030 254008
rect 254086 253952 261114 254008
rect 261170 253952 261175 254008
rect 253430 253950 261175 253952
rect 178604 253948 178610 253950
rect 180149 253947 180215 253950
rect 254025 253947 254091 253950
rect 261109 253947 261175 253950
rect 162117 253874 162183 253877
rect 173566 253874 173572 253876
rect 162117 253872 173572 253874
rect 162117 253816 162122 253872
rect 162178 253816 173572 253872
rect 162117 253814 173572 253816
rect 162117 253811 162183 253814
rect 173566 253812 173572 253814
rect 173636 253874 173642 253876
rect 189073 253874 189139 253877
rect 173636 253872 189139 253874
rect 173636 253816 189078 253872
rect 189134 253816 189139 253872
rect 173636 253814 189139 253816
rect 173636 253812 173642 253814
rect 189073 253811 189139 253814
rect 283097 253874 283163 253877
rect 287094 253874 287100 253876
rect 283097 253872 287100 253874
rect 283097 253816 283102 253872
rect 283158 253816 287100 253872
rect 283097 253814 287100 253816
rect 283097 253811 283163 253814
rect 287094 253812 287100 253814
rect 287164 253812 287170 253876
rect 256734 253738 256740 253740
rect 253460 253678 256740 253738
rect 256734 253676 256740 253678
rect 256804 253676 256810 253740
rect 66989 253602 67055 253605
rect 66989 253600 68908 253602
rect 66989 253544 66994 253600
rect 67050 253544 68908 253600
rect 66989 253542 68908 253544
rect 66989 253539 67055 253542
rect 100845 253330 100911 253333
rect 255497 253330 255563 253333
rect 98716 253328 100911 253330
rect 98716 253272 100850 253328
rect 100906 253272 100911 253328
rect 98716 253270 100911 253272
rect 253460 253328 255563 253330
rect 253460 253272 255502 253328
rect 255558 253272 255563 253328
rect 253460 253270 255563 253272
rect 100845 253267 100911 253270
rect 255497 253267 255563 253270
rect 62113 252786 62179 252789
rect 63401 252786 63467 252789
rect 62113 252784 68908 252786
rect 62113 252728 62118 252784
rect 62174 252728 63406 252784
rect 63462 252728 68908 252784
rect 62113 252726 68908 252728
rect 62113 252723 62179 252726
rect 63401 252723 63467 252726
rect 189073 252650 189139 252653
rect 193630 252650 193690 253028
rect 255405 252786 255471 252789
rect 253460 252784 255471 252786
rect 253460 252728 255410 252784
rect 255466 252728 255471 252784
rect 253460 252726 255471 252728
rect 255405 252723 255471 252726
rect 189073 252648 193690 252650
rect 189073 252592 189078 252648
rect 189134 252592 193690 252648
rect 189073 252590 193690 252592
rect 189073 252587 189139 252590
rect 101254 252514 101260 252516
rect 98716 252454 101260 252514
rect 101254 252452 101260 252454
rect 101324 252452 101330 252516
rect 254945 252514 255011 252517
rect 265934 252514 265940 252516
rect 254945 252512 265940 252514
rect 254945 252456 254950 252512
rect 255006 252456 265940 252512
rect 254945 252454 265940 252456
rect 254945 252451 255011 252454
rect 265934 252452 265940 252454
rect 266004 252452 266010 252516
rect 253430 252242 253490 252348
rect 266629 252242 266695 252245
rect 253430 252240 267750 252242
rect 253430 252184 266634 252240
rect 266690 252184 267750 252240
rect 253430 252182 267750 252184
rect 266629 252179 266695 252182
rect 265065 252106 265131 252109
rect 265750 252106 265756 252108
rect 265065 252104 265756 252106
rect 265065 252048 265070 252104
rect 265126 252048 265756 252104
rect 265065 252046 265756 252048
rect 265065 252043 265131 252046
rect 265750 252044 265756 252046
rect 265820 252044 265826 252108
rect 66805 251970 66871 251973
rect 191005 251970 191071 251973
rect 255405 251970 255471 251973
rect 66805 251968 68908 251970
rect 66805 251912 66810 251968
rect 66866 251912 68908 251968
rect 66805 251910 68908 251912
rect 191005 251968 193660 251970
rect 191005 251912 191010 251968
rect 191066 251912 193660 251968
rect 191005 251910 193660 251912
rect 253460 251968 255471 251970
rect 253460 251912 255410 251968
rect 255466 251912 255471 251968
rect 253460 251910 255471 251912
rect 66805 251907 66871 251910
rect 191005 251907 191071 251910
rect 255405 251907 255471 251910
rect 267690 251834 267750 252182
rect 582465 251834 582531 251837
rect 267690 251832 582531 251834
rect 267690 251776 582470 251832
rect 582526 251776 582531 251832
rect 267690 251774 582531 251776
rect 582465 251771 582531 251774
rect 98134 251292 98194 251668
rect 254025 251562 254091 251565
rect 254945 251562 255011 251565
rect 253460 251560 255011 251562
rect 253460 251504 254030 251560
rect 254086 251504 254950 251560
rect 255006 251504 255011 251560
rect 253460 251502 255011 251504
rect 254025 251499 254091 251502
rect 254945 251499 255011 251502
rect 98126 251228 98132 251292
rect 98196 251228 98202 251292
rect 67725 251154 67791 251157
rect 255497 251154 255563 251157
rect 273110 251154 273116 251156
rect 67725 251152 68908 251154
rect 67725 251096 67730 251152
rect 67786 251096 68908 251152
rect 67725 251094 68908 251096
rect 253460 251152 255563 251154
rect 253460 251096 255502 251152
rect 255558 251096 255563 251152
rect 253460 251094 255563 251096
rect 67725 251091 67791 251094
rect 255497 251091 255563 251094
rect 258030 251094 273116 251154
rect 258030 251018 258090 251094
rect 273110 251092 273116 251094
rect 273180 251092 273186 251156
rect 253430 250958 258090 251018
rect 100845 250882 100911 250885
rect 98716 250880 100911 250882
rect 98716 250824 100850 250880
rect 100906 250824 100911 250880
rect 98716 250822 100911 250824
rect 100845 250819 100911 250822
rect 191649 250882 191715 250885
rect 191649 250880 193660 250882
rect 191649 250824 191654 250880
rect 191710 250824 193660 250880
rect 191649 250822 193660 250824
rect 191649 250819 191715 250822
rect 253430 250716 253490 250958
rect 170397 250474 170463 250477
rect 186313 250474 186379 250477
rect 186814 250474 186820 250476
rect 170397 250472 186820 250474
rect 170397 250416 170402 250472
rect 170458 250416 186318 250472
rect 186374 250416 186820 250472
rect 170397 250414 186820 250416
rect 170397 250411 170463 250414
rect 186313 250411 186379 250414
rect 186814 250412 186820 250414
rect 186884 250412 186890 250476
rect 66805 250338 66871 250341
rect 255405 250338 255471 250341
rect 66805 250336 68908 250338
rect 66805 250280 66810 250336
rect 66866 250280 68908 250336
rect 66805 250278 68908 250280
rect 253460 250336 255471 250338
rect 253460 250280 255410 250336
rect 255466 250280 255471 250336
rect 253460 250278 255471 250280
rect 66805 250275 66871 250278
rect 255405 250275 255471 250278
rect 100937 250066 101003 250069
rect 98716 250064 101003 250066
rect 98716 250008 100942 250064
rect 100998 250008 101003 250064
rect 98716 250006 101003 250008
rect 100937 250003 101003 250006
rect 267917 250068 267983 250069
rect 267917 250064 267964 250068
rect 268028 250066 268034 250068
rect 267917 250008 267922 250064
rect 267917 250004 267964 250008
rect 268028 250006 268074 250066
rect 268028 250004 268034 250006
rect 267917 250003 267983 250004
rect 191005 249794 191071 249797
rect 254209 249794 254275 249797
rect 191005 249792 193660 249794
rect 191005 249736 191010 249792
rect 191066 249736 193660 249792
rect 191005 249734 193660 249736
rect 253460 249792 254275 249794
rect 253460 249736 254214 249792
rect 254270 249736 254275 249792
rect 253460 249734 254275 249736
rect 191005 249731 191071 249734
rect 254209 249731 254275 249734
rect 67817 249522 67883 249525
rect 67817 249520 68908 249522
rect 67817 249464 67822 249520
rect 67878 249464 68908 249520
rect 67817 249462 68908 249464
rect 67817 249459 67883 249462
rect 255497 249386 255563 249389
rect 253460 249384 255563 249386
rect 253460 249328 255502 249384
rect 255558 249328 255563 249384
rect 253460 249326 255563 249328
rect 255497 249323 255563 249326
rect 99557 249250 99623 249253
rect 98716 249248 99623 249250
rect 98716 249192 99562 249248
rect 99618 249192 99623 249248
rect 98716 249190 99623 249192
rect 99557 249187 99623 249190
rect 176193 249114 176259 249117
rect 191782 249114 191788 249116
rect 176193 249112 191788 249114
rect 176193 249056 176198 249112
rect 176254 249056 191788 249112
rect 176193 249054 191788 249056
rect 176193 249051 176259 249054
rect 191782 249052 191788 249054
rect 191852 249052 191858 249116
rect 255405 248978 255471 248981
rect 253460 248976 255471 248978
rect 253460 248920 255410 248976
rect 255466 248920 255471 248976
rect 253460 248918 255471 248920
rect 255405 248915 255471 248918
rect 66437 248706 66503 248709
rect 66437 248704 68908 248706
rect 66437 248648 66442 248704
rect 66498 248648 68908 248704
rect 66437 248646 68908 248648
rect 66437 248643 66503 248646
rect 188286 248508 188292 248572
rect 188356 248570 188362 248572
rect 191557 248570 191623 248573
rect 193630 248570 193690 248676
rect 255313 248570 255379 248573
rect 188356 248568 193690 248570
rect 188356 248512 191562 248568
rect 191618 248512 193690 248568
rect 188356 248510 193690 248512
rect 253460 248568 255379 248570
rect 253460 248512 255318 248568
rect 255374 248512 255379 248568
rect 253460 248510 255379 248512
rect 188356 248508 188362 248510
rect 191557 248507 191623 248510
rect 255313 248507 255379 248510
rect 100845 248434 100911 248437
rect 98716 248432 100911 248434
rect 98716 248376 100850 248432
rect 100906 248376 100911 248432
rect 98716 248374 100911 248376
rect 100845 248371 100911 248374
rect 255497 248434 255563 248437
rect 270769 248434 270835 248437
rect 582465 248434 582531 248437
rect 255497 248432 582531 248434
rect 255497 248376 255502 248432
rect 255558 248376 270774 248432
rect 270830 248376 582470 248432
rect 582526 248376 582531 248432
rect 255497 248374 582531 248376
rect 255497 248371 255563 248374
rect 270769 248371 270835 248374
rect 582465 248371 582531 248374
rect 255497 248162 255563 248165
rect 253460 248160 255563 248162
rect 253460 248104 255502 248160
rect 255558 248104 255563 248160
rect 253460 248102 255563 248104
rect 255497 248099 255563 248102
rect 66805 247890 66871 247893
rect 66805 247888 68908 247890
rect 66805 247832 66810 247888
rect 66866 247832 68908 247888
rect 66805 247830 68908 247832
rect 66805 247827 66871 247830
rect 255405 247754 255471 247757
rect 253460 247752 255471 247754
rect 253460 247696 255410 247752
rect 255466 247696 255471 247752
rect 253460 247694 255471 247696
rect 255405 247691 255471 247694
rect 265065 247754 265131 247757
rect 266486 247754 266492 247756
rect 265065 247752 266492 247754
rect 265065 247696 265070 247752
rect 265126 247696 266492 247752
rect 265065 247694 266492 247696
rect 265065 247691 265131 247694
rect 266486 247692 266492 247694
rect 266556 247692 266562 247756
rect 191741 247618 191807 247621
rect 191741 247616 193660 247618
rect 98134 247077 98194 247588
rect 191741 247560 191746 247616
rect 191802 247560 193660 247616
rect 191741 247558 193660 247560
rect 191741 247555 191807 247558
rect 182081 247482 182147 247485
rect 192334 247482 192340 247484
rect 182081 247480 192340 247482
rect 182081 247424 182086 247480
rect 182142 247424 192340 247480
rect 182081 247422 192340 247424
rect 182081 247419 182147 247422
rect 192334 247420 192340 247422
rect 192404 247420 192410 247484
rect 66662 247012 66668 247076
rect 66732 247074 66738 247076
rect 66732 247014 68908 247074
rect 98085 247072 98194 247077
rect 98085 247016 98090 247072
rect 98146 247016 98194 247072
rect 98085 247014 98194 247016
rect 253430 247074 253490 247180
rect 253430 247014 255330 247074
rect 66732 247012 66738 247014
rect 98085 247011 98151 247014
rect 255270 246938 255330 247014
rect 255270 246878 258090 246938
rect 104249 246802 104315 246805
rect 255497 246802 255563 246805
rect 98716 246800 104315 246802
rect 98716 246744 104254 246800
rect 104310 246744 104315 246800
rect 98716 246742 104315 246744
rect 253460 246800 255563 246802
rect 253460 246744 255502 246800
rect 255558 246744 255563 246800
rect 253460 246742 255563 246744
rect 104249 246739 104315 246742
rect 255497 246739 255563 246742
rect 67449 246258 67515 246261
rect 67449 246256 68908 246258
rect 67449 246200 67454 246256
rect 67510 246200 68908 246256
rect 67449 246198 68908 246200
rect 67449 246195 67515 246198
rect 100661 245986 100727 245989
rect 98716 245984 100727 245986
rect 98716 245928 100666 245984
rect 100722 245928 100727 245984
rect 98716 245926 100727 245928
rect 100661 245923 100727 245926
rect 187693 245850 187759 245853
rect 188981 245850 189047 245853
rect 193438 245850 193444 245852
rect 187693 245848 193444 245850
rect 187693 245792 187698 245848
rect 187754 245792 188986 245848
rect 189042 245792 193444 245848
rect 187693 245790 193444 245792
rect 187693 245787 187759 245790
rect 188981 245787 189047 245790
rect 193438 245788 193444 245790
rect 193508 245788 193514 245852
rect 184790 245652 184796 245716
rect 184860 245714 184866 245716
rect 189073 245714 189139 245717
rect 193630 245714 193690 246500
rect 254117 246394 254183 246397
rect 255313 246394 255379 246397
rect 253460 246392 255379 246394
rect 253460 246336 254122 246392
rect 254178 246336 255318 246392
rect 255374 246336 255379 246392
rect 253460 246334 255379 246336
rect 258030 246394 258090 246878
rect 259494 246394 259500 246396
rect 258030 246334 259500 246394
rect 254117 246331 254183 246334
rect 255313 246331 255379 246334
rect 259494 246332 259500 246334
rect 259564 246394 259570 246396
rect 280286 246394 280292 246396
rect 259564 246334 280292 246394
rect 259564 246332 259570 246334
rect 280286 246332 280292 246334
rect 280356 246332 280362 246396
rect 258165 246258 258231 246261
rect 279417 246258 279483 246261
rect 258030 246256 279483 246258
rect 258030 246200 258170 246256
rect 258226 246200 279422 246256
rect 279478 246200 279483 246256
rect 258030 246198 279483 246200
rect 258030 246122 258090 246198
rect 258165 246195 258231 246198
rect 279417 246195 279483 246198
rect 253430 246062 258090 246122
rect 253430 245956 253490 246062
rect 184860 245712 193690 245714
rect 184860 245656 189078 245712
rect 189134 245656 193690 245712
rect 184860 245654 193690 245656
rect 184860 245652 184866 245654
rect 189073 245651 189139 245654
rect 254526 245652 254532 245716
rect 254596 245714 254602 245716
rect 256734 245714 256740 245716
rect 254596 245654 256740 245714
rect 254596 245652 254602 245654
rect 256734 245652 256740 245654
rect 256804 245652 256810 245716
rect 60457 245578 60523 245581
rect 66846 245578 66852 245580
rect 60457 245576 66852 245578
rect 60457 245520 60462 245576
rect 60518 245520 66852 245576
rect 60457 245518 66852 245520
rect 60457 245515 60523 245518
rect 66846 245516 66852 245518
rect 66916 245516 66922 245580
rect 255405 245578 255471 245581
rect 253460 245576 255471 245578
rect 253460 245520 255410 245576
rect 255466 245520 255471 245576
rect 253460 245518 255471 245520
rect 255405 245515 255471 245518
rect 582465 245578 582531 245581
rect 583520 245578 584960 245668
rect 582465 245576 584960 245578
rect 582465 245520 582470 245576
rect 582526 245520 584960 245576
rect 582465 245518 584960 245520
rect 582465 245515 582531 245518
rect 66110 245380 66116 245444
rect 66180 245442 66186 245444
rect 66180 245382 68908 245442
rect 583520 245428 584960 245518
rect 66180 245380 66186 245382
rect 100845 245170 100911 245173
rect 98716 245168 100911 245170
rect 98716 245112 100850 245168
rect 100906 245112 100911 245168
rect 98716 245110 100911 245112
rect 100845 245107 100911 245110
rect 173709 244626 173775 244629
rect 193630 244626 193690 245412
rect 255405 245170 255471 245173
rect 253460 245168 255471 245170
rect 253460 245112 255410 245168
rect 255466 245112 255471 245168
rect 253460 245110 255471 245112
rect 255405 245107 255471 245110
rect 173709 244624 193690 244626
rect 69430 244356 69490 244596
rect 173709 244568 173714 244624
rect 173770 244568 193690 244624
rect 173709 244566 193690 244568
rect 173709 244563 173775 244566
rect 253062 244493 253122 244732
rect 253013 244488 253122 244493
rect 253013 244432 253018 244488
rect 253074 244432 253122 244488
rect 253013 244430 253122 244432
rect 253013 244427 253079 244430
rect 69422 244292 69428 244356
rect 69492 244292 69498 244356
rect 101029 244354 101095 244357
rect 98716 244352 101095 244354
rect 98716 244296 101034 244352
rect 101090 244296 101095 244352
rect 98716 244294 101095 244296
rect 101029 244291 101095 244294
rect 162669 244354 162735 244357
rect 173157 244354 173223 244357
rect 173709 244354 173775 244357
rect 162669 244352 162778 244354
rect 162669 244296 162674 244352
rect 162730 244296 162778 244352
rect 162669 244291 162778 244296
rect 173157 244352 173775 244354
rect 173157 244296 173162 244352
rect 173218 244296 173714 244352
rect 173770 244296 173775 244352
rect 173157 244294 173775 244296
rect 173157 244291 173223 244294
rect 173709 244291 173775 244294
rect 191281 244354 191347 244357
rect 191649 244354 191715 244357
rect 191281 244352 193660 244354
rect 191281 244296 191286 244352
rect 191342 244296 191654 244352
rect 191710 244296 193660 244352
rect 191281 244294 193660 244296
rect 191281 244291 191347 244294
rect 191649 244291 191715 244294
rect 162718 244218 162778 244291
rect 193673 244218 193739 244221
rect 255497 244218 255563 244221
rect 267774 244218 267780 244220
rect 162718 244216 193739 244218
rect 162718 244160 193678 244216
rect 193734 244160 193739 244216
rect 162718 244158 193739 244160
rect 253460 244216 255563 244218
rect 253460 244160 255502 244216
rect 255558 244160 255563 244216
rect 253460 244158 255563 244160
rect 193673 244155 193739 244158
rect 255497 244155 255563 244158
rect 258030 244158 267780 244218
rect 66713 243810 66779 243813
rect 254117 243810 254183 243813
rect 258030 243810 258090 244158
rect 267774 244156 267780 244158
rect 267844 244156 267850 244220
rect 269614 244156 269620 244220
rect 269684 244218 269690 244220
rect 270401 244218 270467 244221
rect 277158 244218 277164 244220
rect 269684 244216 277164 244218
rect 269684 244160 270406 244216
rect 270462 244160 277164 244216
rect 269684 244158 277164 244160
rect 269684 244156 269690 244158
rect 270401 244155 270467 244158
rect 277158 244156 277164 244158
rect 277228 244156 277234 244220
rect 66713 243808 68908 243810
rect 66713 243752 66718 243808
rect 66774 243752 68908 243808
rect 66713 243750 68908 243752
rect 253460 243808 258090 243810
rect 253460 243752 254122 243808
rect 254178 243752 258090 243808
rect 253460 243750 258090 243752
rect 66713 243747 66779 243750
rect 254117 243747 254183 243750
rect 100845 243538 100911 243541
rect 98716 243536 100911 243538
rect 98716 243480 100850 243536
rect 100906 243480 100911 243536
rect 98716 243478 100911 243480
rect 100845 243475 100911 243478
rect 148593 243538 148659 243541
rect 193254 243538 193260 243540
rect 148593 243536 193260 243538
rect 148593 243480 148598 243536
rect 148654 243480 193260 243536
rect 148593 243478 193260 243480
rect 148593 243475 148659 243478
rect 193254 243476 193260 243478
rect 193324 243476 193330 243540
rect 255865 243402 255931 243405
rect 256734 243402 256740 243404
rect 253460 243400 256740 243402
rect 253460 243344 255870 243400
rect 255926 243344 256740 243400
rect 253460 243342 256740 243344
rect 255865 243339 255931 243342
rect 256734 243340 256740 243342
rect 256804 243340 256810 243404
rect 66846 242932 66852 242996
rect 66916 242994 66922 242996
rect 189717 242994 189783 242997
rect 193630 242994 193690 243236
rect 253606 243204 253612 243268
rect 253676 243266 253682 243268
rect 256785 243266 256851 243269
rect 253676 243264 256851 243266
rect 253676 243208 256790 243264
rect 256846 243208 256851 243264
rect 253676 243206 256851 243208
rect 253676 243204 253682 243206
rect 256785 243203 256851 243206
rect 66916 242934 68908 242994
rect 189717 242992 193690 242994
rect 189717 242936 189722 242992
rect 189778 242936 193690 242992
rect 189717 242934 193690 242936
rect 66916 242932 66922 242934
rect 189717 242931 189783 242934
rect 252878 242861 252938 242964
rect 191833 242860 191899 242861
rect 191782 242858 191788 242860
rect 191742 242798 191788 242858
rect 191852 242856 191899 242860
rect 191894 242800 191899 242856
rect 191782 242796 191788 242798
rect 191852 242796 191899 242800
rect 252878 242856 252987 242861
rect 252878 242800 252926 242856
rect 252982 242800 252987 242856
rect 252878 242798 252987 242800
rect 191833 242795 191899 242796
rect 252921 242795 252987 242798
rect 100845 242722 100911 242725
rect 98716 242720 100911 242722
rect 98716 242664 100850 242720
rect 100906 242664 100911 242720
rect 98716 242662 100911 242664
rect 100845 242659 100911 242662
rect 254209 242586 254275 242589
rect 253460 242584 254275 242586
rect 253460 242528 254214 242584
rect 254270 242528 254275 242584
rect 253460 242526 254275 242528
rect 254209 242523 254275 242526
rect 186221 242450 186287 242453
rect 193581 242450 193647 242453
rect 186221 242448 193647 242450
rect 186221 242392 186226 242448
rect 186282 242392 193586 242448
rect 193642 242392 193647 242448
rect 186221 242390 193647 242392
rect 186221 242387 186287 242390
rect 193581 242387 193647 242390
rect 256785 242314 256851 242317
rect 269062 242314 269068 242316
rect 253430 242312 269068 242314
rect 253430 242256 256790 242312
rect 256846 242256 269068 242312
rect 253430 242254 269068 242256
rect 66805 242178 66871 242181
rect 66805 242176 68908 242178
rect 66805 242120 66810 242176
rect 66866 242120 68908 242176
rect 66805 242118 68908 242120
rect 66805 242115 66871 242118
rect 180558 242116 180564 242180
rect 180628 242178 180634 242180
rect 186313 242178 186379 242181
rect 180628 242176 186379 242178
rect 180628 242120 186318 242176
rect 186374 242120 186379 242176
rect 180628 242118 186379 242120
rect 180628 242116 180634 242118
rect 186313 242115 186379 242118
rect 191741 242178 191807 242181
rect 191741 242176 193660 242178
rect 191741 242120 191746 242176
rect 191802 242120 193660 242176
rect 253430 242148 253490 242254
rect 256785 242251 256851 242254
rect 269062 242252 269068 242254
rect 269132 242252 269138 242316
rect 284293 242178 284359 242181
rect 258030 242176 284359 242178
rect 191741 242118 193660 242120
rect 258030 242120 284298 242176
rect 284354 242120 284359 242176
rect 258030 242118 284359 242120
rect 191741 242115 191807 242118
rect 193254 241980 193260 242044
rect 193324 242042 193330 242044
rect 194501 242042 194567 242045
rect 193324 242040 194567 242042
rect 193324 241984 194506 242040
rect 194562 241984 194567 242040
rect 193324 241982 194567 241984
rect 193324 241980 193330 241982
rect 194501 241979 194567 241982
rect 250161 242042 250227 242045
rect 251030 242042 251036 242044
rect 250161 242040 251036 242042
rect 250161 241984 250166 242040
rect 250222 241984 251036 242040
rect 250161 241982 251036 241984
rect 250161 241979 250227 241982
rect 251030 241980 251036 241982
rect 251100 241980 251106 242044
rect 251766 241980 251772 242044
rect 251836 242042 251842 242044
rect 252921 242042 252987 242045
rect 258030 242042 258090 242118
rect 284293 242115 284359 242118
rect 251836 242040 252987 242042
rect 251836 241984 252926 242040
rect 252982 241984 252987 242040
rect 251836 241982 252987 241984
rect 251836 241980 251842 241982
rect 252921 241979 252987 241982
rect 253430 241982 258090 242042
rect 71129 241770 71195 241773
rect 71630 241770 71636 241772
rect 71129 241768 71636 241770
rect 71129 241712 71134 241768
rect 71190 241712 71636 241768
rect 71129 241710 71636 241712
rect 71129 241707 71195 241710
rect 71630 241708 71636 241710
rect 71700 241708 71706 241772
rect 74901 241770 74967 241773
rect 75678 241770 75684 241772
rect 74901 241768 75684 241770
rect 74901 241712 74906 241768
rect 74962 241712 75684 241768
rect 74901 241710 75684 241712
rect 74901 241707 74967 241710
rect 75678 241708 75684 241710
rect 75748 241708 75754 241772
rect 76649 241770 76715 241773
rect 77150 241770 77156 241772
rect 76649 241768 77156 241770
rect 76649 241712 76654 241768
rect 76710 241712 77156 241768
rect 76649 241710 77156 241712
rect 76649 241707 76715 241710
rect 77150 241708 77156 241710
rect 77220 241708 77226 241772
rect 77661 241770 77727 241773
rect 78397 241772 78463 241773
rect 78070 241770 78076 241772
rect 77661 241768 78076 241770
rect 77661 241712 77666 241768
rect 77722 241712 78076 241768
rect 77661 241710 78076 241712
rect 77661 241707 77727 241710
rect 78070 241708 78076 241710
rect 78140 241708 78146 241772
rect 78397 241770 78444 241772
rect 78352 241768 78444 241770
rect 78352 241712 78402 241768
rect 78352 241710 78444 241712
rect 78397 241708 78444 241710
rect 78508 241708 78514 241772
rect 79869 241770 79935 241773
rect 81985 241772 82051 241773
rect 80646 241770 80652 241772
rect 79869 241768 80652 241770
rect 79869 241712 79874 241768
rect 79930 241712 80652 241768
rect 79869 241710 80652 241712
rect 78397 241707 78463 241708
rect 79869 241707 79935 241710
rect 80646 241708 80652 241710
rect 80716 241708 80722 241772
rect 81934 241708 81940 241772
rect 82004 241770 82051 241772
rect 83733 241770 83799 241773
rect 84510 241770 84516 241772
rect 82004 241768 82096 241770
rect 82046 241712 82096 241768
rect 82004 241710 82096 241712
rect 83733 241768 84516 241770
rect 83733 241712 83738 241768
rect 83794 241712 84516 241768
rect 83733 241710 84516 241712
rect 82004 241708 82051 241710
rect 81985 241707 82051 241708
rect 83733 241707 83799 241710
rect 84510 241708 84516 241710
rect 84580 241708 84586 241772
rect 85941 241770 86007 241773
rect 86585 241772 86651 241773
rect 85941 241768 86418 241770
rect 85941 241712 85946 241768
rect 86002 241712 86418 241768
rect 85941 241710 86418 241712
rect 85941 241707 86007 241710
rect 86358 241634 86418 241710
rect 86534 241708 86540 241772
rect 86604 241770 86651 241772
rect 86604 241768 86696 241770
rect 86646 241712 86696 241768
rect 86604 241710 86696 241712
rect 86604 241708 86651 241710
rect 91134 241708 91140 241772
rect 91204 241770 91210 241772
rect 91553 241770 91619 241773
rect 91204 241768 91619 241770
rect 91204 241712 91558 241768
rect 91614 241712 91619 241768
rect 91204 241710 91619 241712
rect 91204 241708 91210 241710
rect 86585 241707 86651 241708
rect 91553 241707 91619 241710
rect 88006 241634 88012 241636
rect 86358 241574 88012 241634
rect 88006 241572 88012 241574
rect 88076 241572 88082 241636
rect 90265 241634 90331 241637
rect 90817 241634 90883 241637
rect 91502 241634 91508 241636
rect 90265 241632 91508 241634
rect 90265 241576 90270 241632
rect 90326 241576 90822 241632
rect 90878 241576 91508 241632
rect 90265 241574 91508 241576
rect 90265 241571 90331 241574
rect 90817 241571 90883 241574
rect 91502 241572 91508 241574
rect 91572 241572 91578 241636
rect 98686 241634 98746 241876
rect 253430 241740 253490 241982
rect 151169 241634 151235 241637
rect 98686 241632 151235 241634
rect 98686 241576 151174 241632
rect 151230 241576 151235 241632
rect 98686 241574 151235 241576
rect 151169 241571 151235 241574
rect 68870 241436 68876 241500
rect 68940 241498 68946 241500
rect 69289 241498 69355 241501
rect 69565 241498 69631 241501
rect 68940 241496 69631 241498
rect 68940 241440 69294 241496
rect 69350 241440 69570 241496
rect 69626 241440 69631 241496
rect 68940 241438 69631 241440
rect 68940 241436 68946 241438
rect 69289 241435 69355 241438
rect 69565 241435 69631 241438
rect 71313 241498 71379 241501
rect 128997 241498 129063 241501
rect 187049 241498 187115 241501
rect 187550 241498 187556 241500
rect 71313 241496 132510 241498
rect 71313 241440 71318 241496
rect 71374 241440 129002 241496
rect 129058 241440 132510 241496
rect 71313 241438 132510 241440
rect 71313 241435 71379 241438
rect 128997 241435 129063 241438
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 132450 240954 132510 241438
rect 187049 241496 187556 241498
rect 187049 241440 187054 241496
rect 187110 241440 187556 241496
rect 187049 241438 187556 241440
rect 187049 241435 187115 241438
rect 187550 241436 187556 241438
rect 187620 241498 187626 241500
rect 258390 241498 258396 241500
rect 187620 241438 258396 241498
rect 187620 241436 187626 241438
rect 258390 241436 258396 241438
rect 258460 241436 258466 241500
rect 193673 241362 193739 241365
rect 234613 241362 234679 241365
rect 235533 241362 235599 241365
rect 193673 241360 235599 241362
rect 193673 241304 193678 241360
rect 193734 241304 234618 241360
rect 234674 241304 235538 241360
rect 235594 241304 235599 241360
rect 193673 241302 235599 241304
rect 193673 241299 193739 241302
rect 234613 241299 234679 241302
rect 235533 241299 235599 241302
rect 181529 241090 181595 241093
rect 196617 241090 196683 241093
rect 181529 241088 196683 241090
rect 181529 241032 181534 241088
rect 181590 241032 196622 241088
rect 196678 241032 196683 241088
rect 181529 241030 196683 241032
rect 181529 241027 181595 241030
rect 196617 241027 196683 241030
rect 243537 240954 243603 240957
rect 253606 240954 253612 240956
rect 132450 240894 180810 240954
rect 65885 240818 65951 240821
rect 156689 240818 156755 240821
rect 65885 240816 156755 240818
rect 65885 240760 65890 240816
rect 65946 240760 156694 240816
rect 156750 240760 156755 240816
rect 65885 240758 156755 240760
rect 180750 240818 180810 240894
rect 243537 240952 253612 240954
rect 243537 240896 243542 240952
rect 243598 240896 253612 240952
rect 243537 240894 253612 240896
rect 243537 240891 243603 240894
rect 253606 240892 253612 240894
rect 253676 240892 253682 240956
rect 184841 240818 184907 240821
rect 258257 240818 258323 240821
rect 180750 240816 258323 240818
rect 180750 240760 184846 240816
rect 184902 240760 258262 240816
rect 258318 240760 258323 240816
rect 180750 240758 258323 240760
rect 65885 240755 65951 240758
rect 156689 240755 156755 240758
rect 184841 240755 184907 240758
rect 258257 240755 258323 240758
rect 71630 240076 71636 240140
rect 71700 240138 71706 240140
rect 71773 240138 71839 240141
rect 71700 240136 71839 240138
rect 71700 240080 71778 240136
rect 71834 240080 71839 240136
rect 71700 240078 71839 240080
rect 71700 240076 71706 240078
rect 71773 240075 71839 240078
rect 73470 240076 73476 240140
rect 73540 240138 73546 240140
rect 74441 240138 74507 240141
rect 73540 240136 74507 240138
rect 73540 240080 74446 240136
rect 74502 240080 74507 240136
rect 73540 240078 74507 240080
rect 73540 240076 73546 240078
rect 74441 240075 74507 240078
rect 75126 240076 75132 240140
rect 75196 240138 75202 240140
rect 75453 240138 75519 240141
rect 75196 240136 75519 240138
rect 75196 240080 75458 240136
rect 75514 240080 75519 240136
rect 75196 240078 75519 240080
rect 75196 240076 75202 240078
rect 75453 240075 75519 240078
rect 77661 240138 77727 240141
rect 78397 240138 78463 240141
rect 77661 240136 78463 240138
rect 77661 240080 77666 240136
rect 77722 240080 78402 240136
rect 78458 240080 78463 240136
rect 77661 240078 78463 240080
rect 77661 240075 77727 240078
rect 78397 240075 78463 240078
rect 88006 240076 88012 240140
rect 88076 240138 88082 240140
rect 88425 240138 88491 240141
rect 91093 240140 91159 240141
rect 91093 240138 91140 240140
rect 88076 240136 88491 240138
rect 88076 240080 88430 240136
rect 88486 240080 88491 240136
rect 88076 240078 88491 240080
rect 91048 240136 91140 240138
rect 91048 240080 91098 240136
rect 91048 240078 91140 240080
rect 88076 240076 88082 240078
rect 88425 240075 88491 240078
rect 91093 240076 91140 240078
rect 91204 240076 91210 240140
rect 91093 240075 91159 240076
rect 72918 239940 72924 240004
rect 72988 240002 72994 240004
rect 73521 240002 73587 240005
rect 72988 240000 73587 240002
rect 72988 239944 73526 240000
rect 73582 239944 73587 240000
rect 72988 239942 73587 239944
rect 72988 239940 72994 239942
rect 73521 239939 73587 239942
rect 89621 240002 89687 240005
rect 178769 240002 178835 240005
rect 211797 240002 211863 240005
rect 89621 240000 211863 240002
rect 89621 239944 89626 240000
rect 89682 239944 178774 240000
rect 178830 239944 211802 240000
rect 211858 239944 211863 240000
rect 89621 239942 211863 239944
rect 89621 239939 89687 239942
rect 178769 239939 178835 239942
rect 211797 239939 211863 239942
rect 72785 239866 72851 239869
rect 171225 239866 171291 239869
rect 172513 239866 172579 239869
rect 72785 239864 172579 239866
rect 72785 239808 72790 239864
rect 72846 239808 171230 239864
rect 171286 239808 172518 239864
rect 172574 239808 172579 239864
rect 72785 239806 172579 239808
rect 72785 239803 72851 239806
rect 171225 239803 171291 239806
rect 172513 239803 172579 239806
rect 189901 239866 189967 239869
rect 251817 239866 251883 239869
rect 189901 239864 251883 239866
rect 189901 239808 189906 239864
rect 189962 239808 251822 239864
rect 251878 239808 251883 239864
rect 189901 239806 251883 239808
rect 189901 239803 189967 239806
rect 251817 239803 251883 239806
rect 252461 239730 252527 239733
rect 254526 239730 254532 239732
rect 252461 239728 254532 239730
rect 252461 239672 252466 239728
rect 252522 239672 254532 239728
rect 252461 239670 254532 239672
rect 252461 239667 252527 239670
rect 254526 239668 254532 239670
rect 254596 239668 254602 239732
rect 246297 239594 246363 239597
rect 254117 239594 254183 239597
rect 246297 239592 254183 239594
rect 246297 239536 246302 239592
rect 246358 239536 254122 239592
rect 254178 239536 254183 239592
rect 246297 239534 254183 239536
rect 246297 239531 246363 239534
rect 254117 239531 254183 239534
rect 50889 239458 50955 239461
rect 72877 239458 72943 239461
rect 50889 239456 72943 239458
rect 50889 239400 50894 239456
rect 50950 239400 72882 239456
rect 72938 239400 72943 239456
rect 50889 239398 72943 239400
rect 50889 239395 50955 239398
rect 72877 239395 72943 239398
rect 91921 239458 91987 239461
rect 103513 239458 103579 239461
rect 91921 239456 103579 239458
rect 91921 239400 91926 239456
rect 91982 239400 103518 239456
rect 103574 239400 103579 239456
rect 91921 239398 103579 239400
rect 91921 239395 91987 239398
rect 103513 239395 103579 239398
rect 172513 239458 172579 239461
rect 247493 239458 247559 239461
rect 172513 239456 247559 239458
rect 172513 239400 172518 239456
rect 172574 239400 247498 239456
rect 247554 239400 247559 239456
rect 172513 239398 247559 239400
rect 172513 239395 172579 239398
rect 247493 239395 247559 239398
rect 250529 239458 250595 239461
rect 261109 239458 261175 239461
rect 250529 239456 261175 239458
rect 250529 239400 250534 239456
rect 250590 239400 261114 239456
rect 261170 239400 261175 239456
rect 250529 239398 261175 239400
rect 250529 239395 250595 239398
rect 261109 239395 261175 239398
rect 68870 238852 68876 238916
rect 68940 238914 68946 238916
rect 76557 238914 76623 238917
rect 68940 238912 76623 238914
rect 68940 238856 76562 238912
rect 76618 238856 76623 238912
rect 68940 238854 76623 238856
rect 68940 238852 68946 238854
rect 76557 238851 76623 238854
rect 77150 238580 77156 238644
rect 77220 238642 77226 238644
rect 77293 238642 77359 238645
rect 77220 238640 77359 238642
rect 77220 238584 77298 238640
rect 77354 238584 77359 238640
rect 77220 238582 77359 238584
rect 77220 238580 77226 238582
rect 77293 238579 77359 238582
rect 84285 238642 84351 238645
rect 137369 238642 137435 238645
rect 84285 238640 137435 238642
rect 84285 238584 84290 238640
rect 84346 238584 137374 238640
rect 137430 238584 137435 238640
rect 84285 238582 137435 238584
rect 84285 238579 84351 238582
rect 137369 238579 137435 238582
rect 165061 238642 165127 238645
rect 266537 238642 266603 238645
rect 165061 238640 266603 238642
rect 165061 238584 165066 238640
rect 165122 238584 266542 238640
rect 266598 238584 266603 238640
rect 165061 238582 266603 238584
rect 165061 238579 165127 238582
rect 266537 238579 266603 238582
rect 80145 238506 80211 238509
rect 107009 238506 107075 238509
rect 80145 238504 107075 238506
rect 80145 238448 80150 238504
rect 80206 238448 107014 238504
rect 107070 238448 107075 238504
rect 80145 238446 107075 238448
rect 80145 238443 80211 238446
rect 107009 238443 107075 238446
rect 82905 238370 82971 238373
rect 106181 238370 106247 238373
rect 82905 238368 106247 238370
rect 82905 238312 82910 238368
rect 82966 238312 106186 238368
rect 106242 238312 106247 238368
rect 82905 238310 106247 238312
rect 82905 238307 82971 238310
rect 106181 238307 106247 238310
rect 194501 238098 194567 238101
rect 216673 238098 216739 238101
rect 194501 238096 216739 238098
rect 194501 238040 194506 238096
rect 194562 238040 216678 238096
rect 216734 238040 216739 238096
rect 194501 238038 216739 238040
rect 194501 238035 194567 238038
rect 216673 238035 216739 238038
rect 49601 237962 49667 237965
rect 80145 237962 80211 237965
rect 49601 237960 80211 237962
rect 49601 237904 49606 237960
rect 49662 237904 80150 237960
rect 80206 237904 80211 237960
rect 49601 237902 80211 237904
rect 49601 237899 49667 237902
rect 80145 237899 80211 237902
rect 137369 237962 137435 237965
rect 179229 237962 179295 237965
rect 137369 237960 179295 237962
rect 137369 237904 137374 237960
rect 137430 237904 179234 237960
rect 179290 237904 179295 237960
rect 137369 237902 179295 237904
rect 137369 237899 137435 237902
rect 179229 237899 179295 237902
rect 182909 237962 182975 237965
rect 197353 237962 197419 237965
rect 182909 237960 197419 237962
rect 182909 237904 182914 237960
rect 182970 237904 197358 237960
rect 197414 237904 197419 237960
rect 182909 237902 197419 237904
rect 182909 237899 182975 237902
rect 197353 237899 197419 237902
rect 215385 237962 215451 237965
rect 254209 237962 254275 237965
rect 215385 237960 254275 237962
rect 215385 237904 215390 237960
rect 215446 237904 254214 237960
rect 254270 237904 254275 237960
rect 215385 237902 254275 237904
rect 215385 237899 215451 237902
rect 254209 237899 254275 237902
rect 106181 237418 106247 237421
rect 109033 237418 109099 237421
rect 106181 237416 109099 237418
rect 106181 237360 106186 237416
rect 106242 237360 109038 237416
rect 109094 237360 109099 237416
rect 106181 237358 109099 237360
rect 106181 237355 106247 237358
rect 109033 237355 109099 237358
rect 94773 237282 94839 237285
rect 169753 237284 169819 237285
rect 169702 237282 169708 237284
rect 94773 237280 169708 237282
rect 169772 237282 169819 237284
rect 216673 237282 216739 237285
rect 217961 237282 218027 237285
rect 256734 237282 256740 237284
rect 169772 237280 169900 237282
rect 94773 237224 94778 237280
rect 94834 237224 169708 237280
rect 169814 237224 169900 237280
rect 94773 237222 169708 237224
rect 94773 237219 94839 237222
rect 169702 237220 169708 237222
rect 169772 237222 169900 237224
rect 216673 237280 256740 237282
rect 216673 237224 216678 237280
rect 216734 237224 217966 237280
rect 218022 237224 256740 237280
rect 216673 237222 256740 237224
rect 169772 237220 169819 237222
rect 169753 237219 169819 237220
rect 216673 237219 216739 237222
rect 217961 237219 218027 237222
rect 256734 237220 256740 237222
rect 256804 237220 256810 237284
rect 103513 236738 103579 236741
rect 121545 236738 121611 236741
rect 103513 236736 121611 236738
rect 103513 236680 103518 236736
rect 103574 236680 121550 236736
rect 121606 236680 121611 236736
rect 103513 236678 121611 236680
rect 103513 236675 103579 236678
rect 121545 236675 121611 236678
rect 231117 236738 231183 236741
rect 266302 236738 266308 236740
rect 231117 236736 266308 236738
rect 231117 236680 231122 236736
rect 231178 236680 266308 236736
rect 231117 236678 266308 236680
rect 231117 236675 231183 236678
rect 266302 236676 266308 236678
rect 266372 236676 266378 236740
rect 77569 236602 77635 236605
rect 106038 236602 106044 236604
rect 77569 236600 106044 236602
rect 77569 236544 77574 236600
rect 77630 236544 106044 236600
rect 77569 236542 106044 236544
rect 77569 236539 77635 236542
rect 106038 236540 106044 236542
rect 106108 236602 106114 236604
rect 110505 236602 110571 236605
rect 106108 236600 110571 236602
rect 106108 236544 110510 236600
rect 110566 236544 110571 236600
rect 106108 236542 110571 236544
rect 106108 236540 106114 236542
rect 110505 236539 110571 236542
rect 127709 236602 127775 236605
rect 200757 236602 200823 236605
rect 256785 236602 256851 236605
rect 127709 236600 256851 236602
rect 127709 236544 127714 236600
rect 127770 236544 200762 236600
rect 200818 236544 256790 236600
rect 256846 236544 256851 236600
rect 127709 236542 256851 236544
rect 127709 236539 127775 236542
rect 200757 236539 200823 236542
rect 256785 236539 256851 236542
rect 92381 236466 92447 236469
rect 93894 236466 93900 236468
rect 92381 236464 93900 236466
rect 92381 236408 92386 236464
rect 92442 236408 93900 236464
rect 92381 236406 93900 236408
rect 92381 236403 92447 236406
rect 93894 236404 93900 236406
rect 93964 236404 93970 236468
rect 13813 236058 13879 236061
rect 91093 236058 91159 236061
rect 13813 236056 91159 236058
rect 13813 236000 13818 236056
rect 13874 236000 91098 236056
rect 91154 236000 91159 236056
rect 13813 235998 91159 236000
rect 13813 235995 13879 235998
rect 91093 235995 91159 235998
rect 182541 236058 182607 236061
rect 196709 236058 196775 236061
rect 182541 236056 196775 236058
rect 182541 236000 182546 236056
rect 182602 236000 196714 236056
rect 196770 236000 196775 236056
rect 182541 235998 196775 236000
rect 182541 235995 182607 235998
rect 196709 235995 196775 235998
rect 61745 235922 61811 235925
rect 158713 235922 158779 235925
rect 61745 235920 158779 235922
rect 61745 235864 61750 235920
rect 61806 235864 158718 235920
rect 158774 235864 158779 235920
rect 61745 235862 158779 235864
rect 61745 235859 61811 235862
rect 158713 235859 158779 235862
rect 168281 235922 168347 235925
rect 269389 235922 269455 235925
rect 168281 235920 269455 235922
rect 168281 235864 168286 235920
rect 168342 235864 269394 235920
rect 269450 235864 269455 235920
rect 168281 235862 269455 235864
rect 168281 235859 168347 235862
rect 269389 235859 269455 235862
rect 69606 235724 69612 235788
rect 69676 235786 69682 235788
rect 125133 235786 125199 235789
rect 69676 235784 125199 235786
rect 69676 235728 125138 235784
rect 125194 235728 125199 235784
rect 69676 235726 125199 235728
rect 69676 235724 69682 235726
rect 125133 235723 125199 235726
rect 169109 235786 169175 235789
rect 169661 235786 169727 235789
rect 237373 235786 237439 235789
rect 169109 235784 237439 235786
rect 169109 235728 169114 235784
rect 169170 235728 169666 235784
rect 169722 235728 237378 235784
rect 237434 235728 237439 235784
rect 169109 235726 237439 235728
rect 169109 235723 169175 235726
rect 169661 235723 169727 235726
rect 237373 235723 237439 235726
rect 22737 235242 22803 235245
rect 191281 235242 191347 235245
rect 22737 235240 191347 235242
rect 22737 235184 22742 235240
rect 22798 235184 191286 235240
rect 191342 235184 191347 235240
rect 22737 235182 191347 235184
rect 22737 235179 22803 235182
rect 191281 235179 191347 235182
rect 250437 235242 250503 235245
rect 262254 235242 262260 235244
rect 250437 235240 262260 235242
rect 250437 235184 250442 235240
rect 250498 235184 262260 235240
rect 250437 235182 262260 235184
rect 250437 235179 250503 235182
rect 262254 235180 262260 235182
rect 262324 235180 262330 235244
rect 267089 235242 267155 235245
rect 273478 235242 273484 235244
rect 267089 235240 273484 235242
rect 267089 235184 267094 235240
rect 267150 235184 273484 235240
rect 267089 235182 273484 235184
rect 267089 235179 267155 235182
rect 273478 235180 273484 235182
rect 273548 235180 273554 235244
rect 158713 234698 158779 234701
rect 159633 234698 159699 234701
rect 158713 234696 159699 234698
rect 158713 234640 158718 234696
rect 158774 234640 159638 234696
rect 159694 234640 159699 234696
rect 158713 234638 159699 234640
rect 158713 234635 158779 234638
rect 159633 234635 159699 234638
rect 167729 234698 167795 234701
rect 168281 234698 168347 234701
rect 167729 234696 168347 234698
rect 167729 234640 167734 234696
rect 167790 234640 168286 234696
rect 168342 234640 168347 234696
rect 167729 234638 168347 234640
rect 167729 234635 167795 234638
rect 168281 234635 168347 234638
rect 160134 234500 160140 234564
rect 160204 234562 160210 234564
rect 161054 234562 161060 234564
rect 160204 234502 161060 234562
rect 160204 234500 160210 234502
rect 161054 234500 161060 234502
rect 161124 234562 161130 234564
rect 187141 234562 187207 234565
rect 161124 234560 187207 234562
rect 161124 234504 187146 234560
rect 187202 234504 187207 234560
rect 161124 234502 187207 234504
rect 161124 234500 161130 234502
rect 187141 234499 187207 234502
rect 196617 234562 196683 234565
rect 265750 234562 265756 234564
rect 196617 234560 265756 234562
rect 196617 234504 196622 234560
rect 196678 234504 265756 234560
rect 196617 234502 265756 234504
rect 196617 234499 196683 234502
rect 265750 234500 265756 234502
rect 265820 234500 265826 234564
rect 188889 234426 188955 234429
rect 247033 234426 247099 234429
rect 188889 234424 247099 234426
rect 188889 234368 188894 234424
rect 188950 234368 247038 234424
rect 247094 234368 247099 234424
rect 188889 234366 247099 234368
rect 188889 234363 188955 234366
rect 247033 234363 247099 234366
rect 94129 234154 94195 234157
rect 107653 234154 107719 234157
rect 118785 234154 118851 234157
rect 94129 234152 118851 234154
rect 94129 234096 94134 234152
rect 94190 234096 107658 234152
rect 107714 234096 118790 234152
rect 118846 234096 118851 234152
rect 94129 234094 118851 234096
rect 94129 234091 94195 234094
rect 107653 234091 107719 234094
rect 118785 234091 118851 234094
rect 71773 234018 71839 234021
rect 123477 234018 123543 234021
rect 71773 234016 123543 234018
rect 71773 233960 71778 234016
rect 71834 233960 123482 234016
rect 123538 233960 123543 234016
rect 71773 233958 123543 233960
rect 71773 233955 71839 233958
rect 123477 233955 123543 233958
rect 124213 234018 124279 234021
rect 188429 234018 188495 234021
rect 124213 234016 188495 234018
rect 124213 233960 124218 234016
rect 124274 233960 188434 234016
rect 188490 233960 188495 234016
rect 124213 233958 188495 233960
rect 124213 233955 124279 233958
rect 188429 233955 188495 233958
rect 38653 233882 38719 233885
rect 160134 233882 160140 233884
rect 38653 233880 160140 233882
rect 38653 233824 38658 233880
rect 38714 233824 160140 233880
rect 38653 233822 160140 233824
rect 38653 233819 38719 233822
rect 160134 233820 160140 233822
rect 160204 233820 160210 233884
rect 67449 233202 67515 233205
rect 104157 233202 104223 233205
rect 67449 233200 104223 233202
rect 67449 233144 67454 233200
rect 67510 233144 104162 233200
rect 104218 233144 104223 233200
rect 67449 233142 104223 233144
rect 67449 233139 67515 233142
rect 104157 233139 104223 233142
rect 197353 233202 197419 233205
rect 198641 233202 198707 233205
rect 266629 233202 266695 233205
rect 197353 233200 266695 233202
rect 197353 233144 197358 233200
rect 197414 233144 198646 233200
rect 198702 233144 266634 233200
rect 266690 233144 266695 233200
rect 197353 233142 266695 233144
rect 197353 233139 197419 233142
rect 198641 233139 198707 233142
rect 266629 233139 266695 233142
rect 112713 232522 112779 232525
rect 203609 232522 203675 232525
rect 112713 232520 203675 232522
rect 112713 232464 112718 232520
rect 112774 232464 203614 232520
rect 203670 232464 203675 232520
rect 112713 232462 203675 232464
rect 112713 232459 112779 232462
rect 203609 232459 203675 232462
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 166901 231842 166967 231845
rect 267958 231842 267964 231844
rect 166901 231840 267964 231842
rect 166901 231784 166906 231840
rect 166962 231784 267964 231840
rect 166901 231782 267964 231784
rect 166901 231779 166967 231782
rect 267958 231780 267964 231782
rect 268028 231780 268034 231844
rect 181529 231162 181595 231165
rect 260966 231162 260972 231164
rect 181529 231160 260972 231162
rect 181529 231104 181534 231160
rect 181590 231104 260972 231160
rect 181529 231102 260972 231104
rect 181529 231099 181595 231102
rect 260966 231100 260972 231102
rect 261036 231100 261042 231164
rect 93894 230420 93900 230484
rect 93964 230482 93970 230484
rect 100753 230482 100819 230485
rect 93964 230480 100819 230482
rect 93964 230424 100758 230480
rect 100814 230424 100819 230480
rect 93964 230422 100819 230424
rect 93964 230420 93970 230422
rect 100753 230419 100819 230422
rect 193806 230420 193812 230484
rect 193876 230482 193882 230484
rect 222193 230482 222259 230485
rect 193876 230480 222259 230482
rect 193876 230424 222198 230480
rect 222254 230424 222259 230480
rect 193876 230422 222259 230424
rect 193876 230420 193882 230422
rect 222193 230419 222259 230422
rect 228357 230074 228423 230077
rect 251766 230074 251772 230076
rect 228357 230072 251772 230074
rect 228357 230016 228362 230072
rect 228418 230016 251772 230072
rect 228357 230014 251772 230016
rect 228357 230011 228423 230014
rect 251766 230012 251772 230014
rect 251836 230012 251842 230076
rect 213126 229876 213132 229940
rect 213196 229938 213202 229940
rect 252686 229938 252692 229940
rect 213196 229878 252692 229938
rect 213196 229876 213202 229878
rect 252686 229876 252692 229878
rect 252756 229876 252762 229940
rect 180241 229802 180307 229805
rect 231945 229802 232011 229805
rect 263726 229802 263732 229804
rect 180241 229800 263732 229802
rect 180241 229744 180246 229800
rect 180302 229744 231950 229800
rect 232006 229744 263732 229800
rect 180241 229742 263732 229744
rect 180241 229739 180307 229742
rect 231945 229739 232011 229742
rect 263726 229740 263732 229742
rect 263796 229740 263802 229804
rect 248321 228442 248387 228445
rect 258165 228442 258231 228445
rect 248321 228440 258231 228442
rect 248321 228384 248326 228440
rect 248382 228384 258170 228440
rect 258226 228384 258231 228440
rect 248321 228382 258231 228384
rect 248321 228379 248387 228382
rect 258165 228379 258231 228382
rect 148501 228306 148567 228309
rect 235993 228306 236059 228309
rect 262489 228306 262555 228309
rect 148501 228304 262555 228306
rect 148501 228248 148506 228304
rect 148562 228248 235998 228304
rect 236054 228248 262494 228304
rect 262550 228248 262555 228304
rect 148501 228246 262555 228248
rect 148501 228243 148567 228246
rect 235993 228243 236059 228246
rect 262489 228243 262555 228246
rect -960 227884 480 228124
rect 203609 227626 203675 227629
rect 280153 227626 280219 227629
rect 203609 227624 280219 227626
rect 203609 227568 203614 227624
rect 203670 227568 280158 227624
rect 280214 227568 280219 227624
rect 203609 227566 280219 227568
rect 203609 227563 203675 227566
rect 280153 227563 280219 227566
rect 115197 226946 115263 226949
rect 236637 226946 236703 226949
rect 115197 226944 236703 226946
rect 115197 226888 115202 226944
rect 115258 226888 236642 226944
rect 236698 226888 236703 226944
rect 115197 226886 236703 226888
rect 115197 226883 115263 226886
rect 236637 226883 236703 226886
rect 66662 226204 66668 226268
rect 66732 226266 66738 226268
rect 270585 226266 270651 226269
rect 66732 226264 270651 226266
rect 66732 226208 270590 226264
rect 270646 226208 270651 226264
rect 66732 226206 270651 226208
rect 66732 226204 66738 226206
rect 270585 226203 270651 226206
rect 171777 224906 171843 224909
rect 248321 224906 248387 224909
rect 249057 224906 249123 224909
rect 171777 224904 249123 224906
rect 171777 224848 171782 224904
rect 171838 224848 248326 224904
rect 248382 224848 249062 224904
rect 249118 224848 249123 224904
rect 171777 224846 249123 224848
rect 171777 224843 171843 224846
rect 248321 224843 248387 224846
rect 249057 224843 249123 224846
rect 211797 224226 211863 224229
rect 215334 224226 215340 224228
rect 211797 224224 215340 224226
rect 211797 224168 211802 224224
rect 211858 224168 215340 224224
rect 211797 224166 215340 224168
rect 211797 224163 211863 224166
rect 215334 224164 215340 224166
rect 215404 224164 215410 224228
rect 97942 223484 97948 223548
rect 98012 223546 98018 223548
rect 98729 223546 98795 223549
rect 98012 223544 98795 223546
rect 98012 223488 98734 223544
rect 98790 223488 98795 223544
rect 98012 223486 98795 223488
rect 98012 223484 98018 223486
rect 98729 223483 98795 223486
rect 98729 222322 98795 222325
rect 213269 222322 213335 222325
rect 98729 222320 213335 222322
rect 98729 222264 98734 222320
rect 98790 222264 213274 222320
rect 213330 222264 213335 222320
rect 98729 222262 213335 222264
rect 98729 222259 98795 222262
rect 213269 222259 213335 222262
rect 210417 222186 210483 222189
rect 211061 222186 211127 222189
rect 262438 222186 262444 222188
rect 210417 222184 262444 222186
rect 210417 222128 210422 222184
rect 210478 222128 211066 222184
rect 211122 222128 262444 222184
rect 210417 222126 262444 222128
rect 210417 222123 210483 222126
rect 211061 222123 211127 222126
rect 262438 222124 262444 222126
rect 262508 222124 262514 222188
rect 270585 222186 270651 222189
rect 271086 222186 271092 222188
rect 270585 222184 271092 222186
rect 270585 222128 270590 222184
rect 270646 222128 271092 222184
rect 270585 222126 271092 222128
rect 270585 222123 270651 222126
rect 271086 222124 271092 222126
rect 271156 222124 271162 222188
rect 192334 221988 192340 222052
rect 192404 222050 192410 222052
rect 231853 222050 231919 222053
rect 233141 222050 233207 222053
rect 192404 222048 233207 222050
rect 192404 221992 231858 222048
rect 231914 221992 233146 222048
rect 233202 221992 233207 222048
rect 192404 221990 233207 221992
rect 192404 221988 192410 221990
rect 231853 221987 231919 221990
rect 233141 221987 233207 221990
rect 62021 221506 62087 221509
rect 185577 221506 185643 221509
rect 62021 221504 185643 221506
rect 62021 221448 62026 221504
rect 62082 221448 185582 221504
rect 185638 221448 185643 221504
rect 62021 221446 185643 221448
rect 62021 221443 62087 221446
rect 185577 221443 185643 221446
rect 83549 220146 83615 220149
rect 104157 220146 104223 220149
rect 83549 220144 104223 220146
rect 83549 220088 83554 220144
rect 83610 220088 104162 220144
rect 104218 220088 104223 220144
rect 83549 220086 104223 220088
rect 83549 220083 83615 220086
rect 104157 220083 104223 220086
rect 151169 220146 151235 220149
rect 256601 220146 256667 220149
rect 151169 220144 256667 220146
rect 151169 220088 151174 220144
rect 151230 220088 256606 220144
rect 256662 220088 256667 220144
rect 151169 220086 256667 220088
rect 151169 220083 151235 220086
rect 256601 220083 256667 220086
rect 256601 219330 256667 219333
rect 266486 219330 266492 219332
rect 256601 219328 266492 219330
rect 256601 219272 256606 219328
rect 256662 219272 266492 219328
rect 256601 219270 266492 219272
rect 256601 219267 256667 219270
rect 266486 219268 266492 219270
rect 266556 219268 266562 219332
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 56409 218650 56475 218653
rect 163497 218650 163563 218653
rect 56409 218648 163563 218650
rect 56409 218592 56414 218648
rect 56470 218592 163502 218648
rect 163558 218592 163563 218648
rect 56409 218590 163563 218592
rect 56409 218587 56475 218590
rect 163497 218587 163563 218590
rect 247033 217290 247099 217293
rect 248321 217290 248387 217293
rect 259494 217290 259500 217292
rect 247033 217288 259500 217290
rect 247033 217232 247038 217288
rect 247094 217232 248326 217288
rect 248382 217232 259500 217288
rect 247033 217230 259500 217232
rect 247033 217227 247099 217230
rect 248321 217227 248387 217230
rect 259494 217228 259500 217230
rect 259564 217228 259570 217292
rect 101254 216684 101260 216748
rect 101324 216746 101330 216748
rect 101489 216746 101555 216749
rect 285121 216746 285187 216749
rect 101324 216744 285187 216746
rect 101324 216688 101494 216744
rect 101550 216688 285126 216744
rect 285182 216688 285187 216744
rect 101324 216686 285187 216688
rect 101324 216684 101330 216686
rect 101489 216683 101555 216686
rect 285121 216683 285187 216686
rect 204897 216610 204963 216613
rect 263869 216610 263935 216613
rect 204897 216608 263935 216610
rect 204897 216552 204902 216608
rect 204958 216552 263874 216608
rect 263930 216552 263935 216608
rect 204897 216550 263935 216552
rect 204897 216547 204963 216550
rect 263869 216547 263935 216550
rect 2773 215930 2839 215933
rect 189809 215930 189875 215933
rect 2773 215928 189875 215930
rect 2773 215872 2778 215928
rect 2834 215872 189814 215928
rect 189870 215872 189875 215928
rect 2773 215870 189875 215872
rect 2773 215867 2839 215870
rect 189809 215867 189875 215870
rect 204897 215386 204963 215389
rect 205541 215386 205607 215389
rect 204897 215384 205607 215386
rect 204897 215328 204902 215384
rect 204958 215328 205546 215384
rect 205602 215328 205607 215384
rect 204897 215326 205607 215328
rect 204897 215323 204963 215326
rect 205541 215323 205607 215326
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 52361 214570 52427 214573
rect 195973 214570 196039 214573
rect 196617 214570 196683 214573
rect 52361 214568 196683 214570
rect 52361 214512 52366 214568
rect 52422 214512 195978 214568
rect 196034 214512 196622 214568
rect 196678 214512 196683 214568
rect 52361 214510 196683 214512
rect 52361 214507 52427 214510
rect 195973 214507 196039 214510
rect 196617 214507 196683 214510
rect 233877 213210 233943 213213
rect 284477 213210 284543 213213
rect 233877 213208 284543 213210
rect 233877 213152 233882 213208
rect 233938 213152 284482 213208
rect 284538 213152 284543 213208
rect 233877 213150 284543 213152
rect 233877 213147 233943 213150
rect 284477 213147 284543 213150
rect 85573 211850 85639 211853
rect 94078 211850 94084 211852
rect 85573 211848 94084 211850
rect 85573 211792 85578 211848
rect 85634 211792 94084 211848
rect 85573 211790 94084 211792
rect 85573 211787 85639 211790
rect 94078 211788 94084 211790
rect 94148 211788 94154 211852
rect 68870 210972 68876 211036
rect 68940 211034 68946 211036
rect 138013 211034 138079 211037
rect 68940 211032 138079 211034
rect 68940 210976 138018 211032
rect 138074 210976 138079 211032
rect 68940 210974 138079 210976
rect 68940 210972 68946 210974
rect 138013 210971 138079 210974
rect 172329 211034 172395 211037
rect 250529 211034 250595 211037
rect 172329 211032 250595 211034
rect 172329 210976 172334 211032
rect 172390 210976 250534 211032
rect 250590 210976 250595 211032
rect 172329 210974 250595 210976
rect 172329 210971 172395 210974
rect 250529 210971 250595 210974
rect 220077 210898 220143 210901
rect 269614 210898 269620 210900
rect 220077 210896 269620 210898
rect 220077 210840 220082 210896
rect 220138 210840 269620 210896
rect 220077 210838 269620 210840
rect 220077 210835 220143 210838
rect 269614 210836 269620 210838
rect 269684 210836 269690 210900
rect 71630 209612 71636 209676
rect 71700 209674 71706 209676
rect 277669 209674 277735 209677
rect 71700 209672 277735 209674
rect 71700 209616 277674 209672
rect 277730 209616 277735 209672
rect 71700 209614 277735 209616
rect 71700 209612 71706 209614
rect 277669 209611 277735 209614
rect 236637 206954 236703 206957
rect 265065 206954 265131 206957
rect 236637 206952 265131 206954
rect 236637 206896 236642 206952
rect 236698 206896 265070 206952
rect 265126 206896 265131 206952
rect 236637 206894 265131 206896
rect 236637 206891 236703 206894
rect 265065 206891 265131 206894
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 120073 205050 120139 205053
rect 185342 205050 185348 205052
rect 120073 205048 185348 205050
rect 120073 204992 120078 205048
rect 120134 204992 185348 205048
rect 120073 204990 185348 204992
rect 120073 204987 120139 204990
rect 185342 204988 185348 204990
rect 185412 204988 185418 205052
rect 66110 204852 66116 204916
rect 66180 204914 66186 204916
rect 181529 204914 181595 204917
rect 66180 204912 181595 204914
rect 66180 204856 181534 204912
rect 181590 204856 181595 204912
rect 66180 204854 181595 204856
rect 66180 204852 66186 204854
rect 181529 204851 181595 204854
rect 159633 204234 159699 204237
rect 267089 204234 267155 204237
rect 159633 204232 267155 204234
rect 159633 204176 159638 204232
rect 159694 204176 267094 204232
rect 267150 204176 267155 204232
rect 159633 204174 267155 204176
rect 159633 204171 159699 204174
rect 267089 204171 267155 204174
rect 256141 203554 256207 203557
rect 273662 203554 273668 203556
rect 256141 203552 273668 203554
rect 256141 203496 256146 203552
rect 256202 203496 273668 203552
rect 256141 203494 273668 203496
rect 256141 203491 256207 203494
rect 273662 203492 273668 203494
rect 273732 203492 273738 203556
rect 35985 202194 36051 202197
rect 188286 202194 188292 202196
rect 35985 202192 188292 202194
rect 35985 202136 35990 202192
rect 36046 202136 188292 202192
rect 35985 202134 188292 202136
rect 35985 202131 36051 202134
rect 188286 202132 188292 202134
rect 188356 202132 188362 202196
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 65926 192476 65932 192540
rect 65996 192538 66002 192540
rect 128997 192538 129063 192541
rect 65996 192536 129063 192538
rect 65996 192480 129002 192536
rect 129058 192480 129063 192536
rect 65996 192478 129063 192480
rect 65996 192476 66002 192478
rect 128997 192475 129063 192478
rect 214649 192538 214715 192541
rect 223614 192538 223620 192540
rect 214649 192536 223620 192538
rect 214649 192480 214654 192536
rect 214710 192480 223620 192536
rect 214649 192478 223620 192480
rect 214649 192475 214715 192478
rect 223614 192476 223620 192478
rect 223684 192476 223690 192540
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 211797 189682 211863 189685
rect 263542 189682 263548 189684
rect 211797 189680 263548 189682
rect 211797 189624 211802 189680
rect 211858 189624 263548 189680
rect 211797 189622 263548 189624
rect 211797 189619 211863 189622
rect 263542 189620 263548 189622
rect 263612 189620 263618 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 193765 182882 193831 182885
rect 226374 182882 226380 182884
rect 193765 182880 226380 182882
rect 193765 182824 193770 182880
rect 193826 182824 226380 182880
rect 193765 182822 226380 182824
rect 193765 182819 193831 182822
rect 226374 182820 226380 182822
rect 226444 182820 226450 182884
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 83406 177244 83412 177308
rect 83476 177306 83482 177308
rect 83549 177306 83615 177309
rect 207013 177306 207079 177309
rect 83476 177304 207079 177306
rect 83476 177248 83554 177304
rect 83610 177248 207018 177304
rect 207074 177248 207079 177304
rect 83476 177246 207079 177248
rect 83476 177244 83482 177246
rect 83549 177243 83615 177246
rect 207013 177243 207079 177246
rect 82169 176762 82235 176765
rect 82670 176762 82676 176764
rect 82169 176760 82676 176762
rect 82169 176704 82174 176760
rect 82230 176704 82676 176760
rect 82169 176702 82676 176704
rect 82169 176699 82235 176702
rect 82670 176700 82676 176702
rect 82740 176762 82746 176764
rect 205817 176762 205883 176765
rect 82740 176760 205883 176762
rect 82740 176704 205822 176760
rect 205878 176704 205883 176760
rect 82740 176702 205883 176704
rect 82740 176700 82746 176702
rect 205817 176699 205883 176702
rect 207013 176762 207079 176765
rect 207657 176762 207723 176765
rect 207013 176760 207723 176762
rect 207013 176704 207018 176760
rect 207074 176704 207662 176760
rect 207718 176704 207723 176760
rect 207013 176702 207723 176704
rect 207013 176699 207079 176702
rect 207657 176699 207723 176702
rect 76966 176564 76972 176628
rect 77036 176626 77042 176628
rect 172421 176626 172487 176629
rect 77036 176624 172487 176626
rect 77036 176568 172426 176624
rect 172482 176568 172487 176624
rect 77036 176566 172487 176568
rect 77036 176564 77042 176566
rect 172421 176563 172487 176566
rect 75913 176218 75979 176221
rect 76966 176218 76972 176220
rect 75913 176216 76972 176218
rect 75913 176160 75918 176216
rect 75974 176160 76972 176216
rect 75913 176158 76972 176160
rect 75913 176155 75979 176158
rect 76966 176156 76972 176158
rect 77036 176156 77042 176220
rect -960 175796 480 176036
rect 189942 174524 189948 174588
rect 190012 174586 190018 174588
rect 248965 174586 249031 174589
rect 190012 174584 249031 174586
rect 190012 174528 248970 174584
rect 249026 174528 249031 174584
rect 190012 174526 249031 174528
rect 190012 174524 190018 174526
rect 248965 174523 249031 174526
rect 86309 172410 86375 172413
rect 86718 172410 86724 172412
rect 86309 172408 86724 172410
rect 86309 172352 86314 172408
rect 86370 172352 86724 172408
rect 86309 172350 86724 172352
rect 86309 172347 86375 172350
rect 86718 172348 86724 172350
rect 86788 172348 86794 172412
rect 86309 171186 86375 171189
rect 210417 171186 210483 171189
rect 86309 171184 210483 171186
rect 86309 171128 86314 171184
rect 86370 171128 210422 171184
rect 210478 171128 210483 171184
rect 86309 171126 210483 171128
rect 86309 171123 86375 171126
rect 210417 171123 210483 171126
rect 188286 168948 188292 169012
rect 188356 169010 188362 169012
rect 256141 169010 256207 169013
rect 188356 169008 256207 169010
rect 188356 168952 256146 169008
rect 256202 168952 256207 169008
rect 188356 168950 256207 168952
rect 188356 168948 188362 168950
rect 256141 168947 256207 168950
rect 89713 167106 89779 167109
rect 220077 167106 220143 167109
rect 89713 167104 220143 167106
rect 89713 167048 89718 167104
rect 89774 167048 220082 167104
rect 220138 167048 220143 167104
rect 89713 167046 220143 167048
rect 89713 167043 89779 167046
rect 220077 167043 220143 167046
rect 582833 165882 582899 165885
rect 583520 165882 584960 165972
rect 582833 165880 584960 165882
rect 582833 165824 582838 165880
rect 582894 165824 584960 165880
rect 582833 165822 584960 165824
rect 582833 165819 582899 165822
rect 122097 165746 122163 165749
rect 229093 165746 229159 165749
rect 122097 165744 229159 165746
rect 122097 165688 122102 165744
rect 122158 165688 229098 165744
rect 229154 165688 229159 165744
rect 583520 165732 584960 165822
rect 122097 165686 229159 165688
rect 122097 165683 122163 165686
rect 229093 165683 229159 165686
rect 86953 164522 87019 164525
rect 95969 164522 96035 164525
rect 86953 164520 96035 164522
rect 86953 164464 86958 164520
rect 87014 164464 95974 164520
rect 96030 164464 96035 164520
rect 86953 164462 96035 164464
rect 86953 164459 87019 164462
rect 95969 164459 96035 164462
rect 77937 164386 78003 164389
rect 189942 164386 189948 164388
rect 77937 164384 189948 164386
rect 77937 164328 77942 164384
rect 77998 164328 189948 164384
rect 77937 164326 189948 164328
rect 77937 164323 78003 164326
rect 189942 164324 189948 164326
rect 190012 164324 190018 164388
rect 215937 164386 216003 164389
rect 190410 164384 216003 164386
rect 190410 164328 215942 164384
rect 215998 164328 216003 164384
rect 190410 164326 216003 164328
rect 95969 164250 96035 164253
rect 190410 164250 190470 164326
rect 215937 164323 216003 164326
rect 95969 164248 190470 164250
rect 95969 164192 95974 164248
rect 96030 164192 190470 164248
rect 95969 164190 190470 164192
rect 95969 164187 96035 164190
rect 197261 163434 197327 163437
rect 211654 163434 211660 163436
rect 197261 163432 211660 163434
rect 197261 163376 197266 163432
rect 197322 163376 211660 163432
rect 197261 163374 211660 163376
rect 197261 163371 197327 163374
rect 211654 163372 211660 163374
rect 211724 163372 211730 163436
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 142981 162890 143047 162893
rect 231945 162890 232011 162893
rect 142981 162888 232011 162890
rect 142981 162832 142986 162888
rect 143042 162832 231950 162888
rect 232006 162832 232011 162888
rect 142981 162830 232011 162832
rect 142981 162827 143047 162830
rect 231945 162827 232011 162830
rect 66161 162754 66227 162757
rect 154481 162754 154547 162757
rect 66161 162752 154547 162754
rect 66161 162696 66166 162752
rect 66222 162696 154486 162752
rect 154542 162696 154547 162752
rect 66161 162694 154547 162696
rect 66161 162691 66227 162694
rect 154481 162691 154547 162694
rect 236085 162754 236151 162757
rect 236637 162754 236703 162757
rect 236085 162752 236703 162754
rect 236085 162696 236090 162752
rect 236146 162696 236642 162752
rect 236698 162696 236703 162752
rect 236085 162694 236703 162696
rect 236085 162691 236151 162694
rect 236637 162691 236703 162694
rect 114001 161530 114067 161533
rect 236085 161530 236151 161533
rect 114001 161528 236151 161530
rect 114001 161472 114006 161528
rect 114062 161472 236090 161528
rect 236146 161472 236151 161528
rect 114001 161470 236151 161472
rect 114001 161467 114067 161470
rect 236085 161467 236151 161470
rect 59077 160714 59143 160717
rect 158069 160714 158135 160717
rect 59077 160712 158135 160714
rect 59077 160656 59082 160712
rect 59138 160656 158074 160712
rect 158130 160656 158135 160712
rect 59077 160654 158135 160656
rect 59077 160651 59143 160654
rect 158069 160651 158135 160654
rect 138749 160170 138815 160173
rect 227713 160170 227779 160173
rect 228357 160170 228423 160173
rect 138749 160168 228423 160170
rect 138749 160112 138754 160168
rect 138810 160112 227718 160168
rect 227774 160112 228362 160168
rect 228418 160112 228423 160168
rect 138749 160110 228423 160112
rect 138749 160107 138815 160110
rect 227713 160107 227779 160110
rect 228357 160107 228423 160110
rect 213269 159354 213335 159357
rect 281758 159354 281764 159356
rect 213269 159352 281764 159354
rect 213269 159296 213274 159352
rect 213330 159296 281764 159352
rect 213269 159294 281764 159296
rect 213269 159291 213335 159294
rect 281758 159292 281764 159294
rect 281828 159354 281834 159356
rect 316033 159354 316099 159357
rect 281828 159352 316099 159354
rect 281828 159296 316038 159352
rect 316094 159296 316099 159352
rect 281828 159294 316099 159296
rect 281828 159292 281834 159294
rect 316033 159291 316099 159294
rect 154481 158810 154547 158813
rect 234613 158810 234679 158813
rect 154481 158808 234679 158810
rect 154481 158752 154486 158808
rect 154542 158752 234618 158808
rect 234674 158752 234679 158808
rect 154481 158750 234679 158752
rect 154481 158747 154547 158750
rect 234613 158747 234679 158750
rect 198641 158130 198707 158133
rect 205582 158130 205588 158132
rect 198641 158128 205588 158130
rect 198641 158072 198646 158128
rect 198702 158072 205588 158128
rect 198641 158070 205588 158072
rect 198641 158067 198707 158070
rect 205582 158068 205588 158070
rect 205652 158068 205658 158132
rect 192477 157994 192543 157997
rect 200614 157994 200620 157996
rect 192477 157992 200620 157994
rect 192477 157936 192482 157992
rect 192538 157936 200620 157992
rect 192477 157934 200620 157936
rect 192477 157931 192543 157934
rect 200614 157932 200620 157934
rect 200684 157932 200690 157996
rect 72417 157450 72483 157453
rect 193213 157450 193279 157453
rect 193857 157450 193923 157453
rect 72417 157448 193923 157450
rect 72417 157392 72422 157448
rect 72478 157392 193218 157448
rect 193274 157392 193862 157448
rect 193918 157392 193923 157448
rect 72417 157390 193923 157392
rect 72417 157387 72483 157390
rect 193213 157387 193279 157390
rect 193857 157387 193923 157390
rect 196065 157450 196131 157453
rect 196617 157450 196683 157453
rect 303613 157450 303679 157453
rect 196065 157448 303679 157450
rect 196065 157392 196070 157448
rect 196126 157392 196622 157448
rect 196678 157392 303618 157448
rect 303674 157392 303679 157448
rect 196065 157390 303679 157392
rect 196065 157387 196131 157390
rect 196617 157387 196683 157390
rect 303613 157387 303679 157390
rect 240317 156634 240383 156637
rect 276238 156634 276244 156636
rect 238710 156632 276244 156634
rect 238710 156576 240322 156632
rect 240378 156576 276244 156632
rect 238710 156574 276244 156576
rect 175917 156226 175983 156229
rect 238710 156226 238770 156574
rect 240317 156571 240383 156574
rect 276238 156572 276244 156574
rect 276308 156572 276314 156636
rect 175917 156224 238770 156226
rect 175917 156168 175922 156224
rect 175978 156168 238770 156224
rect 175917 156166 238770 156168
rect 175917 156163 175983 156166
rect 82997 156090 83063 156093
rect 211153 156090 211219 156093
rect 82997 156088 211219 156090
rect 82997 156032 83002 156088
rect 83058 156032 211158 156088
rect 211214 156032 211219 156088
rect 82997 156030 211219 156032
rect 82997 156027 83063 156030
rect 211153 156027 211219 156030
rect 70393 155954 70459 155957
rect 71037 155954 71103 155957
rect 70393 155952 71103 155954
rect 70393 155896 70398 155952
rect 70454 155896 71042 155952
rect 71098 155896 71103 155952
rect 70393 155894 71103 155896
rect 70393 155891 70459 155894
rect 71037 155891 71103 155894
rect 205541 155954 205607 155957
rect 209814 155954 209820 155956
rect 205541 155952 209820 155954
rect 205541 155896 205546 155952
rect 205602 155896 209820 155952
rect 205541 155894 209820 155896
rect 205541 155891 205607 155894
rect 209814 155892 209820 155894
rect 209884 155892 209890 155956
rect 70393 154866 70459 154869
rect 188429 154866 188495 154869
rect 70393 154864 188495 154866
rect 70393 154808 70398 154864
rect 70454 154808 188434 154864
rect 188490 154808 188495 154864
rect 70393 154806 188495 154808
rect 70393 154803 70459 154806
rect 188429 154803 188495 154806
rect 153929 154730 153995 154733
rect 222193 154730 222259 154733
rect 153929 154728 222259 154730
rect 153929 154672 153934 154728
rect 153990 154672 222198 154728
rect 222254 154672 222259 154728
rect 153929 154670 222259 154672
rect 153929 154667 153995 154670
rect 222193 154667 222259 154670
rect 187509 154594 187575 154597
rect 252829 154594 252895 154597
rect 187509 154592 252895 154594
rect 187509 154536 187514 154592
rect 187570 154536 252834 154592
rect 252890 154536 252895 154592
rect 187509 154534 252895 154536
rect 187509 154531 187575 154534
rect 252829 154531 252895 154534
rect 193990 153852 193996 153916
rect 194060 153914 194066 153916
rect 215293 153914 215359 153917
rect 194060 153912 215359 153914
rect 194060 153856 215298 153912
rect 215354 153856 215359 153912
rect 194060 153854 215359 153856
rect 194060 153852 194066 153854
rect 215293 153851 215359 153854
rect 148593 153778 148659 153781
rect 200757 153778 200823 153781
rect 233325 153778 233391 153781
rect 148593 153776 233391 153778
rect 148593 153720 148598 153776
rect 148654 153720 200762 153776
rect 200818 153720 233330 153776
rect 233386 153720 233391 153776
rect 148593 153718 233391 153720
rect 148593 153715 148659 153718
rect 200757 153715 200823 153718
rect 233325 153715 233391 153718
rect 66069 153234 66135 153237
rect 159541 153234 159607 153237
rect 66069 153232 159607 153234
rect 66069 153176 66074 153232
rect 66130 153176 159546 153232
rect 159602 153176 159607 153232
rect 66069 153174 159607 153176
rect 66069 153171 66135 153174
rect 159541 153171 159607 153174
rect 244365 153098 244431 153101
rect 245009 153098 245075 153101
rect 244365 153096 245075 153098
rect 244365 153040 244370 153096
rect 244426 153040 245014 153096
rect 245070 153040 245075 153096
rect 244365 153038 245075 153040
rect 244365 153035 244431 153038
rect 245009 153035 245075 153038
rect 582649 152690 582715 152693
rect 583520 152690 584960 152780
rect 582649 152688 584960 152690
rect 582649 152632 582654 152688
rect 582710 152632 584960 152688
rect 582649 152630 584960 152632
rect 582649 152627 582715 152630
rect 583520 152540 584960 152630
rect 27705 152418 27771 152421
rect 189073 152418 189139 152421
rect 27705 152416 189139 152418
rect 27705 152360 27710 152416
rect 27766 152360 189078 152416
rect 189134 152360 189139 152416
rect 27705 152358 189139 152360
rect 27705 152355 27771 152358
rect 189073 152355 189139 152358
rect 145649 151874 145715 151877
rect 244365 151874 244431 151877
rect 145649 151872 244431 151874
rect 145649 151816 145654 151872
rect 145710 151816 244370 151872
rect 244426 151816 244431 151872
rect 145649 151814 244431 151816
rect 145649 151811 145715 151814
rect 244365 151811 244431 151814
rect 208485 151194 208551 151197
rect 281625 151194 281691 151197
rect 208485 151192 281691 151194
rect 208485 151136 208490 151192
rect 208546 151136 281630 151192
rect 281686 151136 281691 151192
rect 208485 151134 281691 151136
rect 208485 151131 208551 151134
rect 281625 151131 281691 151134
rect 88241 151058 88307 151061
rect 100753 151058 100819 151061
rect 88241 151056 100819 151058
rect 88241 151000 88246 151056
rect 88302 151000 100758 151056
rect 100814 151000 100819 151056
rect 88241 150998 100819 151000
rect 88241 150995 88307 150998
rect 100753 150995 100819 150998
rect 102777 151058 102843 151061
rect 211061 151058 211127 151061
rect 227662 151058 227668 151060
rect 102777 151056 227668 151058
rect 102777 151000 102782 151056
rect 102838 151000 211066 151056
rect 211122 151000 227668 151056
rect 102777 150998 227668 151000
rect 102777 150995 102843 150998
rect 211061 150995 211127 150998
rect 227662 150996 227668 150998
rect 227732 150996 227738 151060
rect 67357 150650 67423 150653
rect 104249 150650 104315 150653
rect 67357 150648 104315 150650
rect 67357 150592 67362 150648
rect 67418 150592 104254 150648
rect 104310 150592 104315 150648
rect 67357 150590 104315 150592
rect 67357 150587 67423 150590
rect 104249 150587 104315 150590
rect 102961 150514 103027 150517
rect 230013 150514 230079 150517
rect 102961 150512 230079 150514
rect 102961 150456 102966 150512
rect 103022 150456 230018 150512
rect 230074 150456 230079 150512
rect 102961 150454 230079 150456
rect 102961 150451 103027 150454
rect 230013 150451 230079 150454
rect -960 149834 480 149924
rect 4245 149834 4311 149837
rect -960 149832 4311 149834
rect -960 149776 4250 149832
rect 4306 149776 4311 149832
rect -960 149774 4311 149776
rect -960 149684 480 149774
rect 4245 149771 4311 149774
rect 74717 149698 74783 149701
rect 88977 149698 89043 149701
rect 74717 149696 89043 149698
rect 74717 149640 74722 149696
rect 74778 149640 88982 149696
rect 89038 149640 89043 149696
rect 74717 149638 89043 149640
rect 74717 149635 74783 149638
rect 88977 149635 89043 149638
rect 204437 149698 204503 149701
rect 211797 149698 211863 149701
rect 204437 149696 211863 149698
rect 204437 149640 204442 149696
rect 204498 149640 211802 149696
rect 211858 149640 211863 149696
rect 204437 149638 211863 149640
rect 204437 149635 204503 149638
rect 211797 149635 211863 149638
rect 219433 149562 219499 149565
rect 220169 149562 220235 149565
rect 200070 149560 220235 149562
rect 200070 149504 219438 149560
rect 219494 149504 220174 149560
rect 220230 149504 220235 149560
rect 200070 149502 220235 149504
rect 96286 149228 96292 149292
rect 96356 149290 96362 149292
rect 100702 149290 100708 149292
rect 96356 149230 100708 149290
rect 96356 149228 96362 149230
rect 100702 149228 100708 149230
rect 100772 149228 100778 149292
rect 136081 149290 136147 149293
rect 200070 149290 200130 149502
rect 219433 149499 219499 149502
rect 220169 149499 220235 149502
rect 136081 149288 200130 149290
rect 136081 149232 136086 149288
rect 136142 149232 200130 149288
rect 136081 149230 200130 149232
rect 136081 149227 136147 149230
rect 43989 149154 44055 149157
rect 192334 149154 192340 149156
rect 43989 149152 192340 149154
rect 43989 149096 43994 149152
rect 44050 149096 192340 149152
rect 43989 149094 192340 149096
rect 43989 149091 44055 149094
rect 192334 149092 192340 149094
rect 192404 149092 192410 149156
rect 192477 149154 192543 149157
rect 240041 149154 240107 149157
rect 192477 149152 240107 149154
rect 192477 149096 192482 149152
rect 192538 149096 240046 149152
rect 240102 149096 240107 149152
rect 192477 149094 240107 149096
rect 192477 149091 192543 149094
rect 240041 149091 240107 149094
rect 194542 148276 194548 148340
rect 194612 148338 194618 148340
rect 201585 148338 201651 148341
rect 239397 148338 239463 148341
rect 194612 148336 239463 148338
rect 194612 148280 201590 148336
rect 201646 148280 239402 148336
rect 239458 148280 239463 148336
rect 194612 148278 239463 148280
rect 194612 148276 194618 148278
rect 201585 148275 201651 148278
rect 239397 148275 239463 148278
rect 89161 147794 89227 147797
rect 218329 147794 218395 147797
rect 89161 147792 218395 147794
rect 89161 147736 89166 147792
rect 89222 147736 218334 147792
rect 218390 147736 218395 147792
rect 89161 147734 218395 147736
rect 89161 147731 89227 147734
rect 218329 147731 218395 147734
rect 55029 146978 55095 146981
rect 160921 146978 160987 146981
rect 55029 146976 160987 146978
rect 55029 146920 55034 146976
rect 55090 146920 160926 146976
rect 160982 146920 160987 146976
rect 55029 146918 160987 146920
rect 55029 146915 55095 146918
rect 160921 146915 160987 146918
rect 186957 146570 187023 146573
rect 230473 146570 230539 146573
rect 186957 146568 230539 146570
rect 186957 146512 186962 146568
rect 187018 146512 230478 146568
rect 230534 146512 230539 146568
rect 186957 146510 230539 146512
rect 186957 146507 187023 146510
rect 230473 146507 230539 146510
rect 188521 146434 188587 146437
rect 218789 146434 218855 146437
rect 188521 146432 218855 146434
rect 188521 146376 188526 146432
rect 188582 146376 218794 146432
rect 218850 146376 218855 146432
rect 188521 146374 218855 146376
rect 188521 146371 188587 146374
rect 218789 146371 218855 146374
rect 220077 146434 220143 146437
rect 583109 146434 583175 146437
rect 220077 146432 583175 146434
rect 220077 146376 220082 146432
rect 220138 146376 583114 146432
rect 583170 146376 583175 146432
rect 220077 146374 583175 146376
rect 220077 146371 220143 146374
rect 583109 146371 583175 146374
rect 176009 146298 176075 146301
rect 176561 146298 176627 146301
rect 176009 146296 176627 146298
rect 176009 146240 176014 146296
rect 176070 146240 176566 146296
rect 176622 146240 176627 146296
rect 176009 146238 176627 146240
rect 176009 146235 176075 146238
rect 176561 146235 176627 146238
rect 192334 146236 192340 146300
rect 192404 146298 192410 146300
rect 245101 146298 245167 146301
rect 192404 146296 245167 146298
rect 192404 146240 245106 146296
rect 245162 146240 245167 146296
rect 192404 146238 245167 146240
rect 192404 146236 192410 146238
rect 245101 146235 245167 146238
rect 92473 145618 92539 145621
rect 153929 145618 153995 145621
rect 92473 145616 153995 145618
rect 92473 145560 92478 145616
rect 92534 145560 153934 145616
rect 153990 145560 153995 145616
rect 92473 145558 153995 145560
rect 92473 145555 92539 145558
rect 153929 145555 153995 145558
rect 176009 145074 176075 145077
rect 207105 145074 207171 145077
rect 176009 145072 207171 145074
rect 176009 145016 176014 145072
rect 176070 145016 207110 145072
rect 207166 145016 207171 145072
rect 176009 145014 207171 145016
rect 176009 145011 176075 145014
rect 207105 145011 207171 145014
rect 61837 144938 61903 144941
rect 108481 144938 108547 144941
rect 61837 144936 108547 144938
rect 61837 144880 61842 144936
rect 61898 144880 108486 144936
rect 108542 144880 108547 144936
rect 61837 144878 108547 144880
rect 61837 144875 61903 144878
rect 108481 144875 108547 144878
rect 151169 144938 151235 144941
rect 229737 144938 229803 144941
rect 151169 144936 229803 144938
rect 151169 144880 151174 144936
rect 151230 144880 229742 144936
rect 229798 144880 229803 144936
rect 151169 144878 229803 144880
rect 151169 144875 151235 144878
rect 229737 144875 229803 144878
rect 86861 144802 86927 144805
rect 89846 144802 89852 144804
rect 86861 144800 89852 144802
rect 86861 144744 86866 144800
rect 86922 144744 89852 144800
rect 86861 144742 89852 144744
rect 86861 144739 86927 144742
rect 89846 144740 89852 144742
rect 89916 144740 89922 144804
rect 90817 144802 90883 144805
rect 92606 144802 92612 144804
rect 90817 144800 92612 144802
rect 90817 144744 90822 144800
rect 90878 144744 92612 144800
rect 90817 144742 92612 144744
rect 90817 144739 90883 144742
rect 92606 144740 92612 144742
rect 92676 144740 92682 144804
rect 97349 144802 97415 144805
rect 188337 144804 188403 144805
rect 99966 144802 99972 144804
rect 97349 144800 99972 144802
rect 97349 144744 97354 144800
rect 97410 144744 99972 144800
rect 97349 144742 99972 144744
rect 97349 144739 97415 144742
rect 99966 144740 99972 144742
rect 100036 144740 100042 144804
rect 188286 144740 188292 144804
rect 188356 144802 188403 144804
rect 188356 144800 188448 144802
rect 188398 144744 188448 144800
rect 188356 144742 188448 144744
rect 188356 144740 188403 144742
rect 188337 144739 188403 144740
rect 210509 144122 210575 144125
rect 285765 144122 285831 144125
rect 210509 144120 285831 144122
rect 210509 144064 210514 144120
rect 210570 144064 285770 144120
rect 285826 144064 285831 144120
rect 210509 144062 285831 144064
rect 210509 144059 210575 144062
rect 285765 144059 285831 144062
rect 67909 143850 67975 143853
rect 188337 143850 188403 143853
rect 67909 143848 188403 143850
rect 67909 143792 67914 143848
rect 67970 143792 188342 143848
rect 188398 143792 188403 143848
rect 67909 143790 188403 143792
rect 67909 143787 67975 143790
rect 188337 143787 188403 143790
rect 182909 143714 182975 143717
rect 224350 143714 224356 143716
rect 182909 143712 224356 143714
rect 182909 143656 182914 143712
rect 182970 143656 224356 143712
rect 182909 143654 224356 143656
rect 182909 143651 182975 143654
rect 224350 143652 224356 143654
rect 224420 143652 224426 143716
rect 86125 143578 86191 143581
rect 88742 143578 88748 143580
rect 86125 143576 88748 143578
rect 86125 143520 86130 143576
rect 86186 143520 88748 143576
rect 86125 143518 88748 143520
rect 86125 143515 86191 143518
rect 88742 143516 88748 143518
rect 88812 143516 88818 143580
rect 184381 143578 184447 143581
rect 223614 143578 223620 143580
rect 184381 143576 223620 143578
rect 184381 143520 184386 143576
rect 184442 143520 223620 143576
rect 184381 143518 223620 143520
rect 184381 143515 184447 143518
rect 223614 143516 223620 143518
rect 223684 143516 223690 143580
rect 68686 143380 68692 143444
rect 68756 143442 68762 143444
rect 69105 143442 69171 143445
rect 68756 143440 69171 143442
rect 68756 143384 69110 143440
rect 69166 143384 69171 143440
rect 68756 143382 69171 143384
rect 68756 143380 68762 143382
rect 69105 143379 69171 143382
rect 158713 143442 158779 143445
rect 159357 143442 159423 143445
rect 218237 143442 218303 143445
rect 158713 143440 218303 143442
rect 158713 143384 158718 143440
rect 158774 143384 159362 143440
rect 159418 143384 218242 143440
rect 218298 143384 218303 143440
rect 158713 143382 218303 143384
rect 158713 143379 158779 143382
rect 159357 143379 159423 143382
rect 218237 143379 218303 143382
rect 70158 143244 70164 143308
rect 70228 143306 70234 143308
rect 160737 143306 160803 143309
rect 207013 143306 207079 143309
rect 208117 143306 208183 143309
rect 70228 143304 161490 143306
rect 70228 143248 160742 143304
rect 160798 143248 161490 143304
rect 70228 143246 161490 143248
rect 70228 143244 70234 143246
rect 160737 143243 160803 143246
rect 69013 143034 69079 143037
rect 70158 143034 70164 143036
rect 69013 143032 70164 143034
rect 69013 142976 69018 143032
rect 69074 142976 70164 143032
rect 69013 142974 70164 142976
rect 69013 142971 69079 142974
rect 70158 142972 70164 142974
rect 70228 142972 70234 143036
rect 116853 142762 116919 142765
rect 158713 142762 158779 142765
rect 116853 142760 158779 142762
rect 116853 142704 116858 142760
rect 116914 142704 158718 142760
rect 158774 142704 158779 142760
rect 116853 142702 158779 142704
rect 161430 142762 161490 143246
rect 207013 143304 208183 143306
rect 207013 143248 207018 143304
rect 207074 143248 208122 143304
rect 208178 143248 208183 143304
rect 207013 143246 208183 143248
rect 207013 143243 207079 143246
rect 208117 143243 208183 143246
rect 193305 142900 193371 142901
rect 193254 142898 193260 142900
rect 193214 142838 193260 142898
rect 193324 142896 193371 142900
rect 193366 142840 193371 142896
rect 193254 142836 193260 142838
rect 193324 142836 193371 142840
rect 193305 142835 193371 142836
rect 194685 142762 194751 142765
rect 161430 142760 194751 142762
rect 161430 142704 194690 142760
rect 194746 142704 194751 142760
rect 161430 142702 194751 142704
rect 116853 142699 116919 142702
rect 158713 142699 158779 142702
rect 194685 142699 194751 142702
rect 212809 142490 212875 142493
rect 268377 142490 268443 142493
rect 212809 142488 268443 142490
rect 212809 142432 212814 142488
rect 212870 142432 268382 142488
rect 268438 142432 268443 142488
rect 212809 142430 268443 142432
rect 212809 142427 212875 142430
rect 268377 142427 268443 142430
rect 73286 142292 73292 142356
rect 73356 142354 73362 142356
rect 196617 142354 196683 142357
rect 73356 142352 196683 142354
rect 73356 142296 196622 142352
rect 196678 142296 196683 142352
rect 73356 142294 196683 142296
rect 73356 142292 73362 142294
rect 196617 142291 196683 142294
rect 221917 142354 221983 142357
rect 231209 142354 231275 142357
rect 221917 142352 231275 142354
rect 221917 142296 221922 142352
rect 221978 142296 231214 142352
rect 231270 142296 231275 142352
rect 221917 142294 231275 142296
rect 221917 142291 221983 142294
rect 231209 142291 231275 142294
rect 194685 142218 194751 142221
rect 197854 142218 197860 142220
rect 194685 142216 197860 142218
rect 194685 142160 194690 142216
rect 194746 142160 197860 142216
rect 194685 142158 197860 142160
rect 194685 142155 194751 142158
rect 197854 142156 197860 142158
rect 197924 142156 197930 142220
rect 84694 142020 84700 142084
rect 84764 142082 84770 142084
rect 84837 142082 84903 142085
rect 88425 142082 88491 142085
rect 84764 142080 88491 142082
rect 84764 142024 84842 142080
rect 84898 142024 88430 142080
rect 88486 142024 88491 142080
rect 84764 142022 88491 142024
rect 84764 142020 84770 142022
rect 84837 142019 84903 142022
rect 88425 142019 88491 142022
rect 79961 141402 80027 141405
rect 176009 141402 176075 141405
rect 79961 141400 176075 141402
rect 79961 141344 79966 141400
rect 80022 141344 176014 141400
rect 176070 141344 176075 141400
rect 79961 141342 176075 141344
rect 79961 141339 80027 141342
rect 176009 141339 176075 141342
rect 223757 141402 223823 141405
rect 234613 141402 234679 141405
rect 223757 141400 234679 141402
rect 223757 141344 223762 141400
rect 223818 141344 234618 141400
rect 234674 141344 234679 141400
rect 223757 141342 234679 141344
rect 223757 141339 223823 141342
rect 234613 141339 234679 141342
rect 204253 141130 204319 141133
rect 220169 141130 220235 141133
rect 224902 141130 224908 141132
rect 204253 141128 204362 141130
rect 204253 141072 204258 141128
rect 204314 141072 204362 141128
rect 204253 141067 204362 141072
rect 220169 141128 224908 141130
rect 220169 141072 220174 141128
rect 220230 141072 224908 141128
rect 220169 141070 224908 141072
rect 220169 141067 220235 141070
rect 224902 141068 224908 141070
rect 224972 141068 224978 141132
rect 204302 140994 204362 141067
rect 205449 140994 205515 140997
rect 266997 140994 267063 140997
rect 204302 140992 267063 140994
rect 204302 140936 205454 140992
rect 205510 140936 267002 140992
rect 267058 140936 267063 140992
rect 204302 140934 267063 140936
rect 205449 140931 205515 140934
rect 266997 140931 267063 140934
rect 76966 140796 76972 140860
rect 77036 140858 77042 140860
rect 82077 140858 82143 140861
rect 77036 140856 82143 140858
rect 77036 140800 82082 140856
rect 82138 140800 82143 140856
rect 77036 140798 82143 140800
rect 77036 140796 77042 140798
rect 82077 140795 82143 140798
rect 90817 140858 90883 140861
rect 93342 140858 93348 140860
rect 90817 140856 93348 140858
rect 90817 140800 90822 140856
rect 90878 140800 93348 140856
rect 90817 140798 93348 140800
rect 90817 140795 90883 140798
rect 93342 140796 93348 140798
rect 93412 140858 93418 140860
rect 219985 140858 220051 140861
rect 93412 140856 220051 140858
rect 93412 140800 219990 140856
rect 220046 140800 220051 140856
rect 93412 140798 220051 140800
rect 93412 140796 93418 140798
rect 219985 140795 220051 140798
rect 120165 140722 120231 140725
rect 211889 140722 211955 140725
rect 120165 140720 211955 140722
rect 120165 140664 120170 140720
rect 120226 140664 211894 140720
rect 211950 140664 211955 140720
rect 120165 140662 211955 140664
rect 120165 140659 120231 140662
rect 211889 140659 211955 140662
rect 209497 140586 209563 140589
rect 209998 140586 210004 140588
rect 209497 140584 210004 140586
rect 209497 140528 209502 140584
rect 209558 140528 210004 140584
rect 209497 140526 210004 140528
rect 209497 140523 209563 140526
rect 209998 140524 210004 140526
rect 210068 140524 210074 140588
rect 196566 140388 196572 140452
rect 196636 140450 196642 140452
rect 196801 140450 196867 140453
rect 196636 140448 196867 140450
rect 196636 140392 196806 140448
rect 196862 140392 196867 140448
rect 196636 140390 196867 140392
rect 196636 140388 196642 140390
rect 196801 140387 196867 140390
rect 202873 140450 202939 140453
rect 203190 140450 203196 140452
rect 202873 140448 203196 140450
rect 202873 140392 202878 140448
rect 202934 140392 203196 140448
rect 202873 140390 203196 140392
rect 202873 140387 202939 140390
rect 203190 140388 203196 140390
rect 203260 140450 203266 140452
rect 203517 140450 203583 140453
rect 208209 140452 208275 140453
rect 203260 140448 203583 140450
rect 203260 140392 203522 140448
rect 203578 140392 203583 140448
rect 203260 140390 203583 140392
rect 203260 140388 203266 140390
rect 203517 140387 203583 140390
rect 208158 140388 208164 140452
rect 208228 140450 208275 140452
rect 208228 140448 208320 140450
rect 208270 140392 208320 140448
rect 208228 140390 208320 140392
rect 208228 140388 208275 140390
rect 208209 140387 208275 140388
rect 84745 140042 84811 140045
rect 120165 140042 120231 140045
rect 84745 140040 120231 140042
rect 84745 139984 84750 140040
rect 84806 139984 120170 140040
rect 120226 139984 120231 140040
rect 84745 139982 120231 139984
rect 84745 139979 84811 139982
rect 120165 139979 120231 139982
rect 192937 139906 193003 139909
rect 227989 139906 228055 139909
rect 192937 139904 193660 139906
rect 192937 139848 192942 139904
rect 192998 139848 193660 139904
rect 192937 139846 193660 139848
rect 224940 139904 228055 139906
rect 224940 139848 227994 139904
rect 228050 139848 228055 139904
rect 224940 139846 228055 139848
rect 192937 139843 193003 139846
rect 227989 139843 228055 139846
rect 70209 139634 70275 139637
rect 71814 139634 71820 139636
rect 70209 139632 71820 139634
rect 70209 139576 70214 139632
rect 70270 139576 71820 139632
rect 70209 139574 71820 139576
rect 70209 139571 70275 139574
rect 71814 139572 71820 139574
rect 71884 139572 71890 139636
rect 59261 139498 59327 139501
rect 159357 139498 159423 139501
rect 159633 139498 159699 139501
rect 59261 139496 159699 139498
rect 59261 139440 59266 139496
rect 59322 139440 159362 139496
rect 159418 139440 159638 139496
rect 159694 139440 159699 139496
rect 59261 139438 159699 139440
rect 59261 139435 59327 139438
rect 159357 139435 159423 139438
rect 159633 139435 159699 139438
rect 73613 139362 73679 139365
rect 75310 139362 75316 139364
rect 73613 139360 75316 139362
rect 73613 139304 73618 139360
rect 73674 139304 75316 139360
rect 73613 139302 75316 139304
rect 73613 139299 73679 139302
rect 75310 139300 75316 139302
rect 75380 139300 75386 139364
rect 583017 139362 583083 139365
rect 583520 139362 584960 139452
rect 583017 139360 584960 139362
rect 583017 139304 583022 139360
rect 583078 139304 584960 139360
rect 583017 139302 584960 139304
rect 583017 139299 583083 139302
rect 583520 139212 584960 139302
rect 226333 139090 226399 139093
rect 224940 139088 226399 139090
rect 69422 138620 69428 138684
rect 69492 138682 69498 138684
rect 174537 138682 174603 138685
rect 69492 138680 174603 138682
rect 69492 138624 174542 138680
rect 174598 138624 174603 138680
rect 69492 138622 174603 138624
rect 69492 138620 69498 138622
rect 174537 138619 174603 138622
rect 190361 138682 190427 138685
rect 193254 138682 193260 138684
rect 190361 138680 193260 138682
rect 190361 138624 190366 138680
rect 190422 138624 193260 138680
rect 190361 138622 193260 138624
rect 190361 138619 190427 138622
rect 193254 138620 193260 138622
rect 193324 138620 193330 138684
rect 190269 138546 190335 138549
rect 193630 138546 193690 139060
rect 224940 139032 226338 139088
rect 226394 139032 226399 139088
rect 224940 139030 226399 139032
rect 226333 139027 226399 139030
rect 233325 138954 233391 138957
rect 224910 138952 233391 138954
rect 224910 138896 233330 138952
rect 233386 138896 233391 138952
rect 224910 138894 233391 138896
rect 194174 138756 194180 138820
rect 194244 138756 194250 138820
rect 190269 138544 193690 138546
rect 190269 138488 190274 138544
rect 190330 138488 193690 138544
rect 190269 138486 193690 138488
rect 190269 138483 190335 138486
rect 71313 138274 71379 138277
rect 73286 138274 73292 138276
rect 71313 138272 73292 138274
rect 71313 138216 71318 138272
rect 71374 138216 73292 138272
rect 71313 138214 73292 138216
rect 71313 138211 71379 138214
rect 73286 138212 73292 138214
rect 73356 138212 73362 138276
rect 194182 138244 194242 138756
rect 224910 138244 224970 138894
rect 233325 138891 233391 138894
rect 233325 138682 233391 138685
rect 582649 138682 582715 138685
rect 233325 138680 582715 138682
rect 233325 138624 233330 138680
rect 233386 138624 582654 138680
rect 582710 138624 582715 138680
rect 233325 138622 582715 138624
rect 233325 138619 233391 138622
rect 582649 138619 582715 138622
rect 61929 138138 61995 138141
rect 94865 138138 94931 138141
rect 61929 138136 94931 138138
rect 61929 138080 61934 138136
rect 61990 138080 94870 138136
rect 94926 138080 94931 138136
rect 61929 138078 94931 138080
rect 61929 138075 61995 138078
rect 94865 138075 94931 138078
rect 174537 138138 174603 138141
rect 176009 138138 176075 138141
rect 174537 138136 176075 138138
rect 174537 138080 174542 138136
rect 174598 138080 176014 138136
rect 176070 138080 176075 138136
rect 174537 138078 176075 138080
rect 174537 138075 174603 138078
rect 176009 138075 176075 138078
rect 79593 137322 79659 137325
rect 79910 137322 79916 137324
rect 79593 137320 79916 137322
rect 79593 137264 79598 137320
rect 79654 137264 79916 137320
rect 79593 137262 79916 137264
rect 79593 137259 79659 137262
rect 79910 137260 79916 137262
rect 79980 137260 79986 137324
rect 89069 137322 89135 137325
rect 116853 137322 116919 137325
rect 89069 137320 116919 137322
rect 89069 137264 89074 137320
rect 89130 137264 116858 137320
rect 116914 137264 116919 137320
rect 89069 137262 116919 137264
rect 89069 137259 89135 137262
rect 116853 137259 116919 137262
rect 64781 137050 64847 137053
rect 166441 137050 166507 137053
rect 64781 137048 166507 137050
rect 64781 136992 64786 137048
rect 64842 136992 166446 137048
rect 166502 136992 166507 137048
rect 64781 136990 166507 136992
rect 64781 136987 64847 136990
rect 166441 136987 166507 136990
rect 64689 136914 64755 136917
rect 91001 136914 91067 136917
rect 64689 136912 91067 136914
rect -960 136778 480 136868
rect 64689 136856 64694 136912
rect 64750 136856 91006 136912
rect 91062 136856 91067 136912
rect 64689 136854 91067 136856
rect 64689 136851 64755 136854
rect 91001 136851 91067 136854
rect 2865 136778 2931 136781
rect -960 136776 2931 136778
rect -960 136720 2870 136776
rect 2926 136720 2931 136776
rect -960 136718 2931 136720
rect -960 136628 480 136718
rect 2865 136715 2931 136718
rect 189993 136778 190059 136781
rect 193630 136778 193690 137428
rect 226701 137186 226767 137189
rect 224940 137184 226767 137186
rect 224940 137128 226706 137184
rect 226762 137128 226767 137184
rect 224940 137126 226767 137128
rect 226701 137123 226767 137126
rect 189993 136776 193690 136778
rect 189993 136720 189998 136776
rect 190054 136720 193690 136776
rect 189993 136718 193690 136720
rect 189993 136715 190059 136718
rect 78765 136642 78831 136645
rect 169661 136642 169727 136645
rect 225045 136642 225111 136645
rect 78765 136640 169727 136642
rect 78765 136584 78770 136640
rect 78826 136584 169666 136640
rect 169722 136584 169727 136640
rect 78765 136582 169727 136584
rect 78765 136579 78831 136582
rect 169661 136579 169727 136582
rect 224910 136640 225111 136642
rect 224910 136584 225050 136640
rect 225106 136584 225111 136640
rect 224910 136582 225111 136584
rect 155861 136506 155927 136509
rect 156689 136506 156755 136509
rect 155861 136504 156755 136506
rect 155861 136448 155866 136504
rect 155922 136448 156694 136504
rect 156750 136448 156755 136504
rect 155861 136446 156755 136448
rect 155861 136443 155927 136446
rect 156689 136443 156755 136446
rect 191741 136370 191807 136373
rect 224910 136370 224970 136582
rect 225045 136579 225111 136582
rect 226333 136370 226399 136373
rect 191741 136368 193660 136370
rect 191741 136312 191746 136368
rect 191802 136312 193660 136368
rect 224910 136368 226399 136370
rect 224910 136340 226338 136368
rect 191741 136310 193660 136312
rect 224940 136312 226338 136340
rect 226394 136312 226399 136368
rect 224940 136310 226399 136312
rect 191741 136307 191807 136310
rect 226333 136307 226399 136310
rect 57237 135962 57303 135965
rect 91093 135962 91159 135965
rect 91277 135962 91343 135965
rect 57237 135960 91343 135962
rect 57237 135904 57242 135960
rect 57298 135904 91098 135960
rect 91154 135904 91282 135960
rect 91338 135904 91343 135960
rect 57237 135902 91343 135904
rect 57237 135899 57303 135902
rect 91093 135899 91159 135902
rect 91277 135899 91343 135902
rect 111241 135962 111307 135965
rect 186957 135962 187023 135965
rect 111241 135960 187023 135962
rect 111241 135904 111246 135960
rect 111302 135904 186962 135960
rect 187018 135904 187023 135960
rect 111241 135902 187023 135904
rect 111241 135899 111307 135902
rect 186957 135899 187023 135902
rect 191741 135554 191807 135557
rect 226701 135554 226767 135557
rect 191741 135552 193660 135554
rect 191741 135496 191746 135552
rect 191802 135496 193660 135552
rect 191741 135494 193660 135496
rect 224940 135552 226767 135554
rect 224940 135496 226706 135552
rect 226762 135496 226767 135552
rect 224940 135494 226767 135496
rect 191741 135491 191807 135494
rect 226701 135491 226767 135494
rect 64505 135282 64571 135285
rect 155861 135282 155927 135285
rect 64505 135280 155927 135282
rect 64505 135224 64510 135280
rect 64566 135224 155866 135280
rect 155922 135224 155927 135280
rect 64505 135222 155927 135224
rect 64505 135219 64571 135222
rect 155861 135219 155927 135222
rect 69238 135084 69244 135148
rect 69308 135146 69314 135148
rect 70301 135146 70367 135149
rect 69308 135144 70367 135146
rect 69308 135088 70306 135144
rect 70362 135088 70367 135144
rect 69308 135086 70367 135088
rect 69308 135084 69314 135086
rect 70301 135083 70367 135086
rect 70301 135010 70367 135013
rect 69430 135008 70367 135010
rect 69430 134952 70306 135008
rect 70362 134952 70367 135008
rect 69430 134950 70367 134952
rect 69430 134436 69490 134950
rect 70301 134947 70367 134950
rect 73470 134812 73476 134876
rect 73540 134874 73546 134876
rect 74441 134874 74507 134877
rect 73540 134872 74507 134874
rect 73540 134816 74446 134872
rect 74502 134816 74507 134872
rect 73540 134814 74507 134816
rect 73540 134812 73546 134814
rect 74441 134811 74507 134814
rect 75310 134676 75316 134740
rect 75380 134738 75386 134740
rect 75637 134738 75703 134741
rect 75380 134736 75703 134738
rect 75380 134680 75642 134736
rect 75698 134680 75703 134736
rect 75380 134678 75703 134680
rect 75380 134676 75386 134678
rect 75637 134675 75703 134678
rect 93710 134676 93716 134740
rect 93780 134738 93786 134740
rect 94078 134738 94084 134740
rect 93780 134678 94084 134738
rect 93780 134676 93786 134678
rect 94078 134676 94084 134678
rect 94148 134676 94154 134740
rect 190453 134738 190519 134741
rect 226374 134738 226380 134740
rect 190453 134736 193660 134738
rect 190453 134680 190458 134736
rect 190514 134680 193660 134736
rect 190453 134678 193660 134680
rect 224940 134678 226380 134738
rect 190453 134675 190519 134678
rect 226374 134676 226380 134678
rect 226444 134738 226450 134740
rect 226701 134738 226767 134741
rect 226444 134736 226767 134738
rect 226444 134680 226706 134736
rect 226762 134680 226767 134736
rect 226444 134678 226767 134680
rect 226444 134676 226450 134678
rect 226701 134675 226767 134678
rect 137461 134466 137527 134469
rect 191741 134466 191807 134469
rect 192477 134466 192543 134469
rect 137461 134464 192543 134466
rect 137461 134408 137466 134464
rect 137522 134408 191746 134464
rect 191802 134408 192482 134464
rect 192538 134408 192543 134464
rect 137461 134406 192543 134408
rect 137461 134403 137527 134406
rect 191741 134403 191807 134406
rect 192477 134403 192543 134406
rect 134701 133922 134767 133925
rect 94668 133920 134767 133922
rect 94668 133864 134706 133920
rect 134762 133864 134767 133920
rect 94668 133862 134767 133864
rect 134701 133859 134767 133862
rect 189901 133922 189967 133925
rect 189901 133920 193660 133922
rect 189901 133864 189906 133920
rect 189962 133864 193660 133920
rect 189901 133862 193660 133864
rect 189901 133859 189967 133862
rect 66805 133650 66871 133653
rect 226701 133650 226767 133653
rect 66805 133648 68908 133650
rect 66805 133592 66810 133648
rect 66866 133592 68908 133648
rect 66805 133590 68908 133592
rect 224940 133648 226767 133650
rect 224940 133592 226706 133648
rect 226762 133592 226767 133648
rect 224940 133590 226767 133592
rect 66805 133587 66871 133590
rect 226701 133587 226767 133590
rect 224350 133316 224356 133380
rect 224420 133378 224426 133380
rect 226333 133378 226399 133381
rect 224420 133376 226399 133378
rect 224420 133320 226338 133376
rect 226394 133320 226399 133376
rect 224420 133318 226399 133320
rect 224420 133316 224426 133318
rect 96705 133106 96771 133109
rect 94668 133104 96771 133106
rect 94668 133048 96710 133104
rect 96766 133048 96771 133104
rect 94668 133046 96771 133048
rect 96705 133043 96771 133046
rect 67725 132834 67791 132837
rect 67725 132832 68908 132834
rect 67725 132776 67730 132832
rect 67786 132776 68908 132832
rect 224358 132804 224418 133316
rect 226333 133315 226399 133318
rect 67725 132774 68908 132776
rect 67725 132771 67791 132774
rect 189942 132500 189948 132564
rect 190012 132562 190018 132564
rect 193630 132562 193690 132804
rect 190012 132502 193690 132562
rect 190012 132500 190018 132502
rect 96705 132290 96771 132293
rect 94668 132288 96771 132290
rect 94668 132232 96710 132288
rect 96766 132232 96771 132288
rect 94668 132230 96771 132232
rect 96705 132227 96771 132230
rect 66805 132018 66871 132021
rect 193029 132018 193095 132021
rect 226333 132018 226399 132021
rect 66805 132016 68908 132018
rect 66805 131960 66810 132016
rect 66866 131960 68908 132016
rect 66805 131958 68908 131960
rect 193029 132016 193844 132018
rect 193029 131960 193034 132016
rect 193090 131988 193844 132016
rect 224940 132016 226399 132018
rect 193090 131960 193874 131988
rect 193029 131958 193874 131960
rect 224940 131960 226338 132016
rect 226394 131960 226399 132016
rect 224940 131958 226399 131960
rect 66805 131955 66871 131958
rect 193029 131955 193095 131958
rect 97349 131474 97415 131477
rect 193814 131476 193874 131958
rect 226333 131955 226399 131958
rect 94668 131472 97415 131474
rect 94668 131416 97354 131472
rect 97410 131416 97415 131472
rect 94668 131414 97415 131416
rect 97349 131411 97415 131414
rect 193806 131412 193812 131476
rect 193876 131412 193882 131476
rect 66253 131202 66319 131205
rect 191649 131202 191715 131205
rect 66253 131200 68908 131202
rect 66253 131144 66258 131200
rect 66314 131144 68908 131200
rect 66253 131142 68908 131144
rect 191649 131200 193660 131202
rect 191649 131144 191654 131200
rect 191710 131144 193660 131200
rect 191649 131142 193660 131144
rect 66253 131139 66319 131142
rect 191649 131139 191715 131142
rect 69422 131004 69428 131068
rect 69492 131004 69498 131068
rect 69430 130628 69490 131004
rect 96797 130930 96863 130933
rect 226701 130930 226767 130933
rect 94668 130928 96863 130930
rect 94668 130872 96802 130928
rect 96858 130872 96863 130928
rect 94668 130870 96863 130872
rect 224940 130928 226767 130930
rect 224940 130872 226706 130928
rect 226762 130872 226767 130928
rect 224940 130870 226767 130872
rect 96797 130867 96863 130870
rect 226701 130867 226767 130870
rect 96705 130114 96771 130117
rect 226793 130114 226859 130117
rect 94668 130112 96771 130114
rect 94668 130056 96710 130112
rect 96766 130056 96771 130112
rect 224940 130112 226859 130114
rect 94668 130054 96771 130056
rect 96705 130051 96771 130054
rect 67173 129842 67239 129845
rect 190269 129842 190335 129845
rect 193630 129842 193690 130084
rect 224940 130056 226798 130112
rect 226854 130056 226859 130112
rect 224940 130054 226859 130056
rect 226793 130051 226859 130054
rect 67173 129840 68908 129842
rect 67173 129784 67178 129840
rect 67234 129784 68908 129840
rect 67173 129782 68908 129784
rect 190269 129840 193690 129842
rect 190269 129784 190274 129840
rect 190330 129784 193690 129840
rect 190269 129782 193690 129784
rect 67173 129779 67239 129782
rect 190269 129779 190335 129782
rect 224350 129644 224356 129708
rect 224420 129706 224426 129708
rect 224420 129646 224970 129706
rect 224420 129644 224426 129646
rect 94630 129508 94636 129572
rect 94700 129508 94706 129572
rect 94638 129268 94698 129508
rect 191649 129298 191715 129301
rect 224910 129298 224970 129646
rect 227989 129298 228055 129301
rect 191649 129296 193660 129298
rect 191649 129240 191654 129296
rect 191710 129240 193660 129296
rect 224910 129296 228055 129298
rect 224910 129268 227994 129296
rect 191649 129238 193660 129240
rect 224940 129240 227994 129268
rect 228050 129240 228055 129296
rect 224940 129238 228055 129240
rect 191649 129235 191715 129238
rect 227989 129235 228055 129238
rect 67725 129026 67791 129029
rect 67725 129024 68908 129026
rect 67725 128968 67730 129024
rect 67786 128968 68908 129024
rect 67725 128966 68908 128968
rect 67725 128963 67791 128966
rect 103830 128482 103836 128484
rect 94668 128422 103836 128482
rect 103830 128420 103836 128422
rect 103900 128420 103906 128484
rect 191741 128482 191807 128485
rect 226701 128482 226767 128485
rect 191741 128480 193660 128482
rect 191741 128424 191746 128480
rect 191802 128424 193660 128480
rect 191741 128422 193660 128424
rect 224940 128480 226767 128482
rect 224940 128424 226706 128480
rect 226762 128424 226767 128480
rect 224940 128422 226767 128424
rect 191741 128419 191807 128422
rect 226701 128419 226767 128422
rect 66805 128210 66871 128213
rect 66805 128208 68908 128210
rect 66805 128152 66810 128208
rect 66866 128152 68908 128208
rect 66805 128150 68908 128152
rect 66805 128147 66871 128150
rect 67817 127666 67883 127669
rect 97441 127666 97507 127669
rect 67817 127664 68908 127666
rect 67817 127608 67822 127664
rect 67878 127608 68908 127664
rect 67817 127606 68908 127608
rect 94668 127664 97507 127666
rect 94668 127608 97446 127664
rect 97502 127608 97507 127664
rect 94668 127606 97507 127608
rect 67817 127603 67883 127606
rect 97441 127603 97507 127606
rect 129089 127666 129155 127669
rect 141509 127666 141575 127669
rect 129089 127664 141575 127666
rect 129089 127608 129094 127664
rect 129150 127608 141514 127664
rect 141570 127608 141575 127664
rect 129089 127606 141575 127608
rect 129089 127603 129155 127606
rect 141509 127603 141575 127606
rect 192293 127666 192359 127669
rect 192293 127664 193660 127666
rect 192293 127608 192298 127664
rect 192354 127608 193660 127664
rect 192293 127606 193660 127608
rect 192293 127603 192359 127606
rect 226701 127394 226767 127397
rect 224940 127392 226767 127394
rect 224940 127336 226706 127392
rect 226762 127336 226767 127392
rect 224940 127334 226767 127336
rect 226701 127331 226767 127334
rect 69238 127060 69244 127124
rect 69308 127060 69314 127124
rect 97625 127122 97691 127125
rect 94668 127120 97691 127122
rect 94668 127064 97630 127120
rect 97686 127064 97691 127120
rect 94668 127062 97691 127064
rect 69246 126820 69306 127060
rect 97625 127059 97691 127062
rect 192385 126578 192451 126581
rect 193029 126578 193095 126581
rect 226333 126578 226399 126581
rect 192385 126576 193660 126578
rect 192385 126520 192390 126576
rect 192446 126520 193034 126576
rect 193090 126520 193660 126576
rect 192385 126518 193660 126520
rect 224940 126576 226399 126578
rect 224940 126520 226338 126576
rect 226394 126520 226399 126576
rect 224940 126518 226399 126520
rect 192385 126515 192451 126518
rect 193029 126515 193095 126518
rect 226333 126515 226399 126518
rect 97257 126306 97323 126309
rect 94668 126304 97323 126306
rect 94668 126248 97262 126304
rect 97318 126248 97323 126304
rect 94668 126246 97323 126248
rect 97257 126243 97323 126246
rect 66161 126034 66227 126037
rect 582925 126034 582991 126037
rect 583520 126034 584960 126124
rect 66161 126032 68908 126034
rect 66161 125976 66166 126032
rect 66222 125976 68908 126032
rect 66161 125974 68908 125976
rect 582925 126032 584960 126034
rect 582925 125976 582930 126032
rect 582986 125976 584960 126032
rect 582925 125974 584960 125976
rect 66161 125971 66227 125974
rect 582925 125971 582991 125974
rect 583520 125884 584960 125974
rect 190453 125762 190519 125765
rect 227713 125762 227779 125765
rect 190453 125760 193660 125762
rect 190453 125704 190458 125760
rect 190514 125704 193660 125760
rect 190453 125702 193660 125704
rect 224940 125760 227779 125762
rect 224940 125704 227718 125760
rect 227774 125704 227779 125760
rect 224940 125702 227779 125704
rect 190453 125699 190519 125702
rect 227713 125699 227779 125702
rect 96613 125490 96679 125493
rect 94668 125488 96679 125490
rect 94668 125432 96618 125488
rect 96674 125432 96679 125488
rect 94668 125430 96679 125432
rect 96613 125427 96679 125430
rect 67909 125218 67975 125221
rect 67909 125216 68908 125218
rect 67909 125160 67914 125216
rect 67970 125160 68908 125216
rect 67909 125158 68908 125160
rect 67909 125155 67975 125158
rect 192937 124946 193003 124949
rect 192937 124944 193660 124946
rect 192937 124888 192942 124944
rect 192998 124888 193660 124944
rect 192937 124886 193660 124888
rect 192937 124883 193003 124886
rect 97533 124674 97599 124677
rect 226517 124674 226583 124677
rect 94668 124672 97599 124674
rect 94668 124616 97538 124672
rect 97594 124616 97599 124672
rect 94668 124614 97599 124616
rect 224940 124672 226583 124674
rect 224940 124616 226522 124672
rect 226578 124616 226583 124672
rect 224940 124614 226583 124616
rect 97533 124611 97599 124614
rect 226517 124611 226583 124614
rect 66897 124402 66963 124405
rect 66897 124400 68908 124402
rect 66897 124344 66902 124400
rect 66958 124344 68908 124400
rect 66897 124342 68908 124344
rect 66897 124339 66963 124342
rect 97901 124130 97967 124133
rect 94668 124128 97967 124130
rect 94668 124072 97906 124128
rect 97962 124072 97967 124128
rect 94668 124070 97967 124072
rect 97901 124067 97967 124070
rect 126605 124130 126671 124133
rect 193213 124130 193279 124133
rect 193438 124130 193444 124132
rect 126605 124128 193444 124130
rect 126605 124072 126610 124128
rect 126666 124072 193218 124128
rect 193274 124072 193444 124128
rect 126605 124070 193444 124072
rect 126605 124067 126671 124070
rect 193213 124067 193279 124070
rect 193438 124068 193444 124070
rect 193508 124068 193514 124132
rect 66805 123858 66871 123861
rect 66805 123856 68908 123858
rect -960 123572 480 123812
rect 66805 123800 66810 123856
rect 66866 123800 68908 123856
rect 66805 123798 68908 123800
rect 66805 123795 66871 123798
rect 192702 123796 192708 123860
rect 192772 123858 192778 123860
rect 225229 123858 225295 123861
rect 192772 123798 193660 123858
rect 224940 123856 225295 123858
rect 224940 123800 225234 123856
rect 225290 123800 225295 123856
rect 224940 123798 225295 123800
rect 192772 123796 192778 123798
rect 225229 123795 225295 123798
rect 97165 123314 97231 123317
rect 94668 123312 97231 123314
rect 94668 123256 97170 123312
rect 97226 123256 97231 123312
rect 94668 123254 97231 123256
rect 97165 123251 97231 123254
rect 66253 123042 66319 123045
rect 191741 123042 191807 123045
rect 226333 123042 226399 123045
rect 66253 123040 68908 123042
rect 66253 122984 66258 123040
rect 66314 122984 68908 123040
rect 66253 122982 68908 122984
rect 191741 123040 193660 123042
rect 191741 122984 191746 123040
rect 191802 122984 193660 123040
rect 191741 122982 193660 122984
rect 224940 123040 226399 123042
rect 224940 122984 226338 123040
rect 226394 122984 226399 123040
rect 224940 122982 226399 122984
rect 66253 122979 66319 122982
rect 191741 122979 191807 122982
rect 226333 122979 226399 122982
rect 97533 122498 97599 122501
rect 94668 122496 97599 122498
rect 94668 122440 97538 122496
rect 97594 122440 97599 122496
rect 94668 122438 97599 122440
rect 97533 122435 97599 122438
rect 66345 122226 66411 122229
rect 226333 122226 226399 122229
rect 66345 122224 68908 122226
rect 66345 122168 66350 122224
rect 66406 122168 68908 122224
rect 224940 122224 226399 122226
rect 66345 122166 68908 122168
rect 66345 122163 66411 122166
rect 138749 121682 138815 121685
rect 94668 121680 138815 121682
rect 94668 121624 138754 121680
rect 138810 121624 138815 121680
rect 94668 121622 138815 121624
rect 138749 121619 138815 121622
rect 190453 121682 190519 121685
rect 193630 121682 193690 122196
rect 224940 122168 226338 122224
rect 226394 122168 226399 122224
rect 224940 122166 226399 122168
rect 226333 122163 226399 122166
rect 190453 121680 193690 121682
rect 190453 121624 190458 121680
rect 190514 121624 193690 121680
rect 190453 121622 193690 121624
rect 190453 121619 190519 121622
rect 65977 121410 66043 121413
rect 191189 121410 191255 121413
rect 65977 121408 68908 121410
rect 65977 121352 65982 121408
rect 66038 121352 68908 121408
rect 65977 121350 68908 121352
rect 191189 121408 193660 121410
rect 191189 121352 191194 121408
rect 191250 121352 193660 121408
rect 191189 121350 193660 121352
rect 65977 121347 66043 121350
rect 191189 121347 191255 121350
rect 227662 121138 227668 121140
rect 224940 121078 227668 121138
rect 227662 121076 227668 121078
rect 227732 121076 227738 121140
rect 97717 120866 97783 120869
rect 94668 120864 97783 120866
rect 94668 120808 97722 120864
rect 97778 120808 97783 120864
rect 94668 120806 97783 120808
rect 97717 120803 97783 120806
rect 43989 120730 44055 120733
rect 66897 120730 66963 120733
rect 43989 120728 66963 120730
rect 43989 120672 43994 120728
rect 44050 120672 66902 120728
rect 66958 120672 66963 120728
rect 43989 120670 66963 120672
rect 43989 120667 44055 120670
rect 66897 120667 66963 120670
rect 127709 120730 127775 120733
rect 184054 120730 184060 120732
rect 127709 120728 184060 120730
rect 127709 120672 127714 120728
rect 127770 120672 184060 120728
rect 127709 120670 184060 120672
rect 127709 120667 127775 120670
rect 184054 120668 184060 120670
rect 184124 120730 184130 120732
rect 184749 120730 184815 120733
rect 184124 120728 184815 120730
rect 184124 120672 184754 120728
rect 184810 120672 184815 120728
rect 184124 120670 184815 120672
rect 184124 120668 184130 120670
rect 184749 120667 184815 120670
rect 66805 120594 66871 120597
rect 66805 120592 68908 120594
rect 66805 120536 66810 120592
rect 66866 120536 68908 120592
rect 66805 120534 68908 120536
rect 66805 120531 66871 120534
rect 95325 120322 95391 120325
rect 97533 120322 97599 120325
rect 94668 120320 97599 120322
rect 94668 120264 95330 120320
rect 95386 120264 97538 120320
rect 97594 120264 97599 120320
rect 94668 120262 97599 120264
rect 95325 120259 95391 120262
rect 97533 120259 97599 120262
rect 191741 120322 191807 120325
rect 226425 120322 226491 120325
rect 191741 120320 193660 120322
rect 191741 120264 191746 120320
rect 191802 120264 193660 120320
rect 191741 120262 193660 120264
rect 224940 120320 226491 120322
rect 224940 120264 226430 120320
rect 226486 120264 226491 120320
rect 224940 120262 226491 120264
rect 191741 120259 191807 120262
rect 226425 120259 226491 120262
rect 66805 120050 66871 120053
rect 66805 120048 68908 120050
rect 66805 119992 66810 120048
rect 66866 119992 68908 120048
rect 66805 119990 68908 119992
rect 66805 119987 66871 119990
rect 224902 119988 224908 120052
rect 224972 119988 224978 120052
rect 97717 119506 97783 119509
rect 94668 119504 97783 119506
rect 94668 119448 97722 119504
rect 97778 119448 97783 119504
rect 94668 119446 97783 119448
rect 97717 119443 97783 119446
rect 191741 119506 191807 119509
rect 191741 119504 193660 119506
rect 191741 119448 191746 119504
rect 191802 119448 193660 119504
rect 224910 119476 224970 119988
rect 191741 119446 193660 119448
rect 191741 119443 191807 119446
rect 66897 119234 66963 119237
rect 66897 119232 68908 119234
rect 66897 119176 66902 119232
rect 66958 119176 68908 119232
rect 66897 119174 68908 119176
rect 66897 119171 66963 119174
rect 97901 118690 97967 118693
rect 94668 118688 97967 118690
rect 94668 118632 97906 118688
rect 97962 118632 97967 118688
rect 94668 118630 97967 118632
rect 97901 118627 97967 118630
rect 191741 118690 191807 118693
rect 191741 118688 193660 118690
rect 191741 118632 191746 118688
rect 191802 118632 193660 118688
rect 191741 118630 193660 118632
rect 191741 118627 191807 118630
rect 66805 118418 66871 118421
rect 226517 118418 226583 118421
rect 66805 118416 68908 118418
rect 66805 118360 66810 118416
rect 66866 118360 68908 118416
rect 66805 118358 68908 118360
rect 224940 118416 226583 118418
rect 224940 118360 226522 118416
rect 226578 118360 226583 118416
rect 224940 118358 226583 118360
rect 66805 118355 66871 118358
rect 226517 118355 226583 118358
rect 102777 117874 102843 117877
rect 94668 117872 102843 117874
rect 94668 117816 102782 117872
rect 102838 117816 102843 117872
rect 94668 117814 102843 117816
rect 102777 117811 102843 117814
rect 66897 117602 66963 117605
rect 191097 117602 191163 117605
rect 226701 117602 226767 117605
rect 66897 117600 68908 117602
rect 66897 117544 66902 117600
rect 66958 117544 68908 117600
rect 66897 117542 68908 117544
rect 191097 117600 193660 117602
rect 191097 117544 191102 117600
rect 191158 117544 193660 117600
rect 191097 117542 193660 117544
rect 224940 117600 226767 117602
rect 224940 117544 226706 117600
rect 226762 117544 226767 117600
rect 224940 117542 226767 117544
rect 66897 117539 66963 117542
rect 191097 117539 191163 117542
rect 226701 117539 226767 117542
rect 233877 117194 233943 117197
rect 291285 117194 291351 117197
rect 291653 117194 291719 117197
rect 233877 117192 291719 117194
rect 233877 117136 233882 117192
rect 233938 117136 291290 117192
rect 291346 117136 291658 117192
rect 291714 117136 291719 117192
rect 233877 117134 291719 117136
rect 233877 117131 233943 117134
rect 291285 117131 291351 117134
rect 291653 117131 291719 117134
rect 66069 117058 66135 117061
rect 97349 117058 97415 117061
rect 66069 117056 68908 117058
rect 66069 117000 66074 117056
rect 66130 117000 68908 117056
rect 66069 116998 68908 117000
rect 94668 117056 97415 117058
rect 94668 117000 97354 117056
rect 97410 117000 97415 117056
rect 94668 116998 97415 117000
rect 66069 116995 66135 116998
rect 97349 116995 97415 116998
rect 191281 116786 191347 116789
rect 227897 116786 227963 116789
rect 191281 116784 193660 116786
rect 191281 116728 191286 116784
rect 191342 116728 193660 116784
rect 191281 116726 193660 116728
rect 224940 116784 227963 116786
rect 224940 116728 227902 116784
rect 227958 116728 227963 116784
rect 224940 116726 227963 116728
rect 191281 116723 191347 116726
rect 227897 116723 227963 116726
rect 97901 116514 97967 116517
rect 94668 116512 97967 116514
rect 94668 116456 97906 116512
rect 97962 116456 97967 116512
rect 94668 116454 97967 116456
rect 97901 116451 97967 116454
rect 66805 116242 66871 116245
rect 66805 116240 68908 116242
rect 66805 116184 66810 116240
rect 66866 116184 68908 116240
rect 66805 116182 68908 116184
rect 66805 116179 66871 116182
rect 191741 115970 191807 115973
rect 226701 115970 226767 115973
rect 191741 115968 193660 115970
rect 191741 115912 191746 115968
rect 191802 115912 193660 115968
rect 191741 115910 193660 115912
rect 224940 115968 226767 115970
rect 224940 115912 226706 115968
rect 226762 115912 226767 115968
rect 224940 115910 226767 115912
rect 191741 115907 191807 115910
rect 226701 115907 226767 115910
rect 97901 115698 97967 115701
rect 94668 115696 97967 115698
rect 94668 115640 97906 115696
rect 97962 115640 97967 115696
rect 94668 115638 97967 115640
rect 97901 115635 97967 115638
rect 66805 115426 66871 115429
rect 66805 115424 68908 115426
rect 66805 115368 66810 115424
rect 66866 115368 68908 115424
rect 66805 115366 68908 115368
rect 66805 115363 66871 115366
rect 191005 115154 191071 115157
rect 191005 115152 193660 115154
rect 191005 115096 191010 115152
rect 191066 115096 193660 115152
rect 191005 115094 193660 115096
rect 191005 115091 191071 115094
rect 97809 114882 97875 114885
rect 226333 114882 226399 114885
rect 94668 114880 97875 114882
rect 94668 114824 97814 114880
rect 97870 114824 97875 114880
rect 94668 114822 97875 114824
rect 224940 114880 226399 114882
rect 224940 114824 226338 114880
rect 226394 114824 226399 114880
rect 224940 114822 226399 114824
rect 97809 114819 97875 114822
rect 226333 114819 226399 114822
rect 66805 114610 66871 114613
rect 66805 114608 68908 114610
rect 66805 114552 66810 114608
rect 66866 114552 68908 114608
rect 66805 114550 68908 114552
rect 66805 114547 66871 114550
rect 252737 114474 252803 114477
rect 253013 114474 253079 114477
rect 224910 114472 253079 114474
rect 224910 114416 252742 114472
rect 252798 114416 253018 114472
rect 253074 114416 253079 114472
rect 224910 114414 253079 114416
rect 96705 114066 96771 114069
rect 94668 114064 96771 114066
rect 94668 114008 96710 114064
rect 96766 114008 96771 114064
rect 94668 114006 96771 114008
rect 96705 114003 96771 114006
rect 191741 114066 191807 114069
rect 191741 114064 193660 114066
rect 191741 114008 191746 114064
rect 191802 114008 193660 114064
rect 224910 114036 224970 114414
rect 252737 114411 252803 114414
rect 253013 114411 253079 114414
rect 191741 114006 193660 114008
rect 191741 114003 191807 114006
rect 66805 113794 66871 113797
rect 66805 113792 68908 113794
rect 66805 113736 66810 113792
rect 66866 113736 68908 113792
rect 66805 113734 68908 113736
rect 66805 113731 66871 113734
rect 101990 113732 101996 113796
rect 102060 113794 102066 113796
rect 150433 113794 150499 113797
rect 227621 113794 227687 113797
rect 102060 113792 150499 113794
rect 102060 113736 150438 113792
rect 150494 113736 150499 113792
rect 102060 113734 150499 113736
rect 102060 113732 102066 113734
rect 150433 113731 150499 113734
rect 224910 113792 227687 113794
rect 224910 113736 227626 113792
rect 227682 113736 227687 113792
rect 224910 113734 227687 113736
rect 97533 113522 97599 113525
rect 94668 113520 97599 113522
rect 94668 113464 97538 113520
rect 97594 113464 97599 113520
rect 94668 113462 97599 113464
rect 97533 113459 97599 113462
rect 65977 113250 66043 113253
rect 191189 113250 191255 113253
rect 65977 113248 68908 113250
rect 65977 113192 65982 113248
rect 66038 113192 68908 113248
rect 65977 113190 68908 113192
rect 191189 113248 193660 113250
rect 191189 113192 191194 113248
rect 191250 113192 193660 113248
rect 224910 113220 224970 113734
rect 227621 113731 227687 113734
rect 253013 113250 253079 113253
rect 258717 113250 258783 113253
rect 253013 113248 258783 113250
rect 191189 113190 193660 113192
rect 253013 113192 253018 113248
rect 253074 113192 258722 113248
rect 258778 113192 258783 113248
rect 253013 113190 258783 113192
rect 65977 113187 66043 113190
rect 191189 113187 191255 113190
rect 253013 113187 253079 113190
rect 258717 113187 258783 113190
rect 583109 112842 583175 112845
rect 583520 112842 584960 112932
rect 583109 112840 584960 112842
rect 583109 112784 583114 112840
rect 583170 112784 584960 112840
rect 583109 112782 584960 112784
rect 583109 112779 583175 112782
rect 97901 112706 97967 112709
rect 94668 112704 97967 112706
rect 94668 112648 97906 112704
rect 97962 112648 97967 112704
rect 583520 112692 584960 112782
rect 94668 112646 97967 112648
rect 97901 112643 97967 112646
rect 66805 112434 66871 112437
rect 66805 112432 68908 112434
rect 66805 112376 66810 112432
rect 66866 112376 68908 112432
rect 66805 112374 68908 112376
rect 66805 112371 66871 112374
rect 96889 111890 96955 111893
rect 94668 111888 96955 111890
rect 94668 111832 96894 111888
rect 96950 111832 96955 111888
rect 94668 111830 96955 111832
rect 96889 111827 96955 111830
rect 159357 111890 159423 111893
rect 193630 111890 193690 112404
rect 226701 112162 226767 112165
rect 224940 112160 226767 112162
rect 224940 112104 226706 112160
rect 226762 112104 226767 112160
rect 224940 112102 226767 112104
rect 226701 112099 226767 112102
rect 159357 111888 193690 111890
rect 159357 111832 159362 111888
rect 159418 111832 193690 111888
rect 159357 111830 193690 111832
rect 159357 111827 159423 111830
rect 66897 111618 66963 111621
rect 66897 111616 68908 111618
rect 66897 111560 66902 111616
rect 66958 111560 68908 111616
rect 66897 111558 68908 111560
rect 66897 111555 66963 111558
rect 226333 111346 226399 111349
rect 224940 111344 226399 111346
rect 97349 111074 97415 111077
rect 94668 111072 97415 111074
rect 94668 111016 97354 111072
rect 97410 111016 97415 111072
rect 94668 111014 97415 111016
rect 97349 111011 97415 111014
rect 66805 110802 66871 110805
rect 190269 110802 190335 110805
rect 193630 110802 193690 111316
rect 224940 111288 226338 111344
rect 226394 111288 226399 111344
rect 224940 111286 226399 111288
rect 226333 111283 226399 111286
rect 66805 110800 68908 110802
rect -960 110666 480 110756
rect 66805 110744 66810 110800
rect 66866 110744 68908 110800
rect 66805 110742 68908 110744
rect 190269 110800 193690 110802
rect 190269 110744 190274 110800
rect 190330 110744 193690 110800
rect 190269 110742 193690 110744
rect 66805 110739 66871 110742
rect 190269 110739 190335 110742
rect 2865 110666 2931 110669
rect -960 110664 2931 110666
rect -960 110608 2870 110664
rect 2926 110608 2931 110664
rect -960 110606 2931 110608
rect -960 110516 480 110606
rect 2865 110603 2931 110606
rect 191373 110530 191439 110533
rect 226517 110530 226583 110533
rect 191373 110528 193660 110530
rect 191373 110472 191378 110528
rect 191434 110472 193660 110528
rect 191373 110470 193660 110472
rect 224940 110528 226583 110530
rect 224940 110472 226522 110528
rect 226578 110472 226583 110528
rect 224940 110470 226583 110472
rect 191373 110467 191439 110470
rect 226517 110467 226583 110470
rect 66897 110258 66963 110261
rect 98085 110258 98151 110261
rect 66897 110256 68908 110258
rect 66897 110200 66902 110256
rect 66958 110200 68908 110256
rect 66897 110198 68908 110200
rect 94668 110256 98151 110258
rect 94668 110200 98090 110256
rect 98146 110200 98151 110256
rect 94668 110198 98151 110200
rect 66897 110195 66963 110198
rect 98085 110195 98151 110198
rect 97809 109714 97875 109717
rect 94668 109712 97875 109714
rect 94668 109656 97814 109712
rect 97870 109656 97875 109712
rect 94668 109654 97875 109656
rect 97809 109651 97875 109654
rect 191557 109714 191623 109717
rect 225137 109714 225203 109717
rect 191557 109712 193660 109714
rect 191557 109656 191562 109712
rect 191618 109656 193660 109712
rect 191557 109654 193660 109656
rect 224940 109712 225203 109714
rect 224940 109656 225142 109712
rect 225198 109656 225203 109712
rect 224940 109654 225203 109656
rect 191557 109651 191623 109654
rect 225137 109651 225203 109654
rect 97206 109516 97212 109580
rect 97276 109578 97282 109580
rect 111885 109578 111951 109581
rect 97276 109576 111951 109578
rect 97276 109520 111890 109576
rect 111946 109520 111951 109576
rect 97276 109518 111951 109520
rect 97276 109516 97282 109518
rect 111885 109515 111951 109518
rect 66805 109442 66871 109445
rect 66805 109440 68908 109442
rect 66805 109384 66810 109440
rect 66866 109384 68908 109440
rect 66805 109382 68908 109384
rect 66805 109379 66871 109382
rect 96286 108898 96292 108900
rect 94668 108838 96292 108898
rect 96286 108836 96292 108838
rect 96356 108836 96362 108900
rect 191189 108898 191255 108901
rect 191189 108896 193660 108898
rect 191189 108840 191194 108896
rect 191250 108840 193660 108896
rect 191189 108838 193660 108840
rect 191189 108835 191255 108838
rect 66437 108626 66503 108629
rect 227069 108626 227135 108629
rect 66437 108624 68908 108626
rect 66437 108568 66442 108624
rect 66498 108568 68908 108624
rect 66437 108566 68908 108568
rect 224940 108624 227135 108626
rect 224940 108568 227074 108624
rect 227130 108568 227135 108624
rect 224940 108566 227135 108568
rect 66437 108563 66503 108566
rect 227069 108563 227135 108566
rect 97901 108082 97967 108085
rect 94668 108080 97967 108082
rect 94668 108024 97906 108080
rect 97962 108024 97967 108080
rect 94668 108022 97967 108024
rect 97901 108019 97967 108022
rect 66713 107810 66779 107813
rect 191189 107810 191255 107813
rect 226374 107810 226380 107812
rect 66713 107808 68908 107810
rect 66713 107752 66718 107808
rect 66774 107752 68908 107808
rect 66713 107750 68908 107752
rect 191189 107808 193660 107810
rect 191189 107752 191194 107808
rect 191250 107752 193660 107808
rect 191189 107750 193660 107752
rect 224940 107750 226380 107810
rect 66713 107747 66779 107750
rect 191189 107747 191255 107750
rect 226374 107748 226380 107750
rect 226444 107810 226450 107812
rect 226517 107810 226583 107813
rect 226444 107808 226583 107810
rect 226444 107752 226522 107808
rect 226578 107752 226583 107808
rect 226444 107750 226583 107752
rect 226444 107748 226450 107750
rect 226517 107747 226583 107750
rect 96981 107266 97047 107269
rect 94668 107264 97047 107266
rect 94668 107208 96986 107264
rect 97042 107208 97047 107264
rect 94668 107206 97047 107208
rect 96981 107203 97047 107206
rect 66989 106994 67055 106997
rect 67357 106994 67423 106997
rect 191741 106994 191807 106997
rect 226701 106994 226767 106997
rect 66989 106992 68908 106994
rect 66989 106936 66994 106992
rect 67050 106936 67362 106992
rect 67418 106936 68908 106992
rect 66989 106934 68908 106936
rect 191741 106992 193660 106994
rect 191741 106936 191746 106992
rect 191802 106936 193660 106992
rect 191741 106934 193660 106936
rect 224940 106992 226767 106994
rect 224940 106936 226706 106992
rect 226762 106936 226767 106992
rect 224940 106934 226767 106936
rect 66989 106931 67055 106934
rect 67357 106931 67423 106934
rect 191741 106931 191807 106934
rect 226701 106931 226767 106934
rect 187049 106722 187115 106725
rect 94668 106720 187115 106722
rect 94668 106664 187054 106720
rect 187110 106664 187115 106720
rect 94668 106662 187115 106664
rect 187049 106659 187115 106662
rect 64638 106252 64644 106316
rect 64708 106314 64714 106316
rect 68878 106314 68938 106420
rect 64708 106254 68938 106314
rect 64708 106252 64714 106254
rect 191741 106178 191807 106181
rect 191741 106176 193660 106178
rect 191741 106120 191746 106176
rect 191802 106120 193660 106176
rect 191741 106118 193660 106120
rect 191741 106115 191807 106118
rect 97533 105906 97599 105909
rect 226701 105906 226767 105909
rect 94668 105904 97599 105906
rect 94668 105848 97538 105904
rect 97594 105848 97599 105904
rect 94668 105846 97599 105848
rect 224940 105904 226767 105906
rect 224940 105848 226706 105904
rect 226762 105848 226767 105904
rect 224940 105846 226767 105848
rect 97533 105843 97599 105846
rect 226701 105843 226767 105846
rect 66529 105634 66595 105637
rect 66529 105632 68908 105634
rect 66529 105576 66534 105632
rect 66590 105576 68908 105632
rect 66529 105574 68908 105576
rect 66529 105571 66595 105574
rect 96889 105090 96955 105093
rect 94668 105088 96955 105090
rect 94668 105032 96894 105088
rect 96950 105032 96955 105088
rect 94668 105030 96955 105032
rect 96889 105027 96955 105030
rect 191741 105090 191807 105093
rect 191741 105088 193660 105090
rect 191741 105032 191746 105088
rect 191802 105032 193660 105088
rect 191741 105030 193660 105032
rect 191741 105027 191807 105030
rect 224910 104954 224970 105060
rect 225045 104954 225111 104957
rect 224910 104952 225111 104954
rect 224910 104896 225050 104952
rect 225106 104896 225111 104952
rect 224910 104894 225111 104896
rect 225045 104891 225111 104894
rect 66345 104818 66411 104821
rect 66345 104816 68908 104818
rect 66345 104760 66350 104816
rect 66406 104760 68908 104816
rect 66345 104758 68908 104760
rect 66345 104755 66411 104758
rect 97717 104274 97783 104277
rect 94668 104272 97783 104274
rect 94668 104216 97722 104272
rect 97778 104216 97783 104272
rect 94668 104214 97783 104216
rect 97717 104211 97783 104214
rect 191741 104274 191807 104277
rect 193213 104274 193279 104277
rect 226517 104274 226583 104277
rect 191741 104272 193660 104274
rect 191741 104216 191746 104272
rect 191802 104216 193218 104272
rect 193274 104216 193660 104272
rect 191741 104214 193660 104216
rect 224940 104272 226583 104274
rect 224940 104216 226522 104272
rect 226578 104216 226583 104272
rect 224940 104214 226583 104216
rect 191741 104211 191807 104214
rect 193213 104211 193279 104214
rect 226517 104211 226583 104214
rect 98729 104138 98795 104141
rect 114737 104138 114803 104141
rect 98729 104136 114803 104138
rect 98729 104080 98734 104136
rect 98790 104080 114742 104136
rect 114798 104080 114803 104136
rect 98729 104078 114803 104080
rect 98729 104075 98795 104078
rect 114737 104075 114803 104078
rect 67265 104002 67331 104005
rect 67265 104000 68908 104002
rect 67265 103944 67270 104000
rect 67326 103944 68908 104000
rect 67265 103942 68908 103944
rect 67265 103939 67331 103942
rect 96521 103594 96587 103597
rect 96521 103592 96630 103594
rect 96521 103536 96526 103592
rect 96582 103536 96630 103592
rect 96521 103531 96630 103536
rect 96570 103458 96630 103531
rect 94668 103398 96630 103458
rect 191649 103458 191715 103461
rect 226701 103458 226767 103461
rect 191649 103456 193660 103458
rect 191649 103400 191654 103456
rect 191710 103400 193660 103456
rect 191649 103398 193660 103400
rect 224940 103456 226767 103458
rect 224940 103400 226706 103456
rect 226762 103400 226767 103456
rect 224940 103398 226767 103400
rect 191649 103395 191715 103398
rect 226701 103395 226767 103398
rect 66529 103186 66595 103189
rect 66529 103184 68908 103186
rect 66529 103128 66534 103184
rect 66590 103128 68908 103184
rect 66529 103126 68908 103128
rect 66529 103123 66595 103126
rect 97901 102914 97967 102917
rect 94668 102912 97967 102914
rect 94668 102856 97906 102912
rect 97962 102856 97967 102912
rect 94668 102854 97967 102856
rect 97901 102851 97967 102854
rect 66621 102642 66687 102645
rect 191097 102642 191163 102645
rect 66621 102640 68908 102642
rect 66621 102584 66626 102640
rect 66682 102584 68908 102640
rect 66621 102582 68908 102584
rect 191097 102640 193660 102642
rect 191097 102584 191102 102640
rect 191158 102584 193660 102640
rect 191097 102582 193660 102584
rect 66621 102579 66687 102582
rect 191097 102579 191163 102582
rect 226701 102370 226767 102373
rect 224940 102368 226767 102370
rect 224940 102312 226706 102368
rect 226762 102312 226767 102368
rect 224940 102310 226767 102312
rect 226701 102307 226767 102310
rect 97901 102098 97967 102101
rect 94668 102096 97967 102098
rect 94668 102040 97906 102096
rect 97962 102040 97967 102096
rect 94668 102038 97967 102040
rect 97901 102035 97967 102038
rect 66805 101826 66871 101829
rect 66805 101824 68908 101826
rect 66805 101768 66810 101824
rect 66866 101768 68908 101824
rect 66805 101766 68908 101768
rect 66805 101763 66871 101766
rect 191649 101554 191715 101557
rect 226333 101554 226399 101557
rect 191649 101552 193660 101554
rect 191649 101496 191654 101552
rect 191710 101496 193660 101552
rect 191649 101494 193660 101496
rect 224940 101552 226399 101554
rect 224940 101496 226338 101552
rect 226394 101496 226399 101552
rect 224940 101494 226399 101496
rect 191649 101491 191715 101494
rect 226333 101491 226399 101494
rect 97901 101282 97967 101285
rect 94668 101280 97967 101282
rect 94668 101224 97906 101280
rect 97962 101224 97967 101280
rect 94668 101222 97967 101224
rect 97901 101219 97967 101222
rect 67817 101010 67883 101013
rect 67817 101008 68908 101010
rect 67817 100952 67822 101008
rect 67878 100952 68908 101008
rect 67817 100950 68908 100952
rect 67817 100947 67883 100950
rect 191557 100738 191623 100741
rect 226333 100738 226399 100741
rect 191557 100736 193660 100738
rect 191557 100680 191562 100736
rect 191618 100680 193660 100736
rect 191557 100678 193660 100680
rect 224940 100736 226399 100738
rect 224940 100680 226338 100736
rect 226394 100680 226399 100736
rect 224940 100678 226399 100680
rect 191557 100675 191623 100678
rect 226333 100675 226399 100678
rect 97533 100466 97599 100469
rect 94668 100464 97599 100466
rect 94668 100408 97538 100464
rect 97594 100408 97599 100464
rect 94668 100406 97599 100408
rect 97533 100403 97599 100406
rect 67265 100194 67331 100197
rect 67265 100192 68908 100194
rect 67265 100136 67270 100192
rect 67326 100136 68908 100192
rect 67265 100134 68908 100136
rect 67265 100131 67331 100134
rect 190637 99922 190703 99925
rect 190637 99920 193660 99922
rect 190637 99864 190642 99920
rect 190698 99864 193660 99920
rect 190637 99862 193660 99864
rect 190637 99859 190703 99862
rect 66805 99650 66871 99653
rect 97901 99650 97967 99653
rect 226425 99650 226491 99653
rect 66805 99648 68908 99650
rect 66805 99592 66810 99648
rect 66866 99592 68908 99648
rect 66805 99590 68908 99592
rect 94668 99648 97967 99650
rect 94668 99592 97906 99648
rect 97962 99592 97967 99648
rect 94668 99590 97967 99592
rect 224940 99648 226491 99650
rect 224940 99592 226430 99648
rect 226486 99592 226491 99648
rect 224940 99590 226491 99592
rect 66805 99587 66871 99590
rect 97901 99587 97967 99590
rect 226425 99587 226491 99590
rect 98637 99514 98703 99517
rect 191557 99514 191623 99517
rect 98637 99512 191623 99514
rect 98637 99456 98642 99512
rect 98698 99456 191562 99512
rect 191618 99456 191623 99512
rect 98637 99454 191623 99456
rect 98637 99451 98703 99454
rect 191557 99451 191623 99454
rect 583017 99514 583083 99517
rect 583520 99514 584960 99604
rect 583017 99512 584960 99514
rect 583017 99456 583022 99512
rect 583078 99456 584960 99512
rect 583017 99454 584960 99456
rect 583017 99451 583083 99454
rect 583520 99364 584960 99454
rect 96889 99106 96955 99109
rect 94668 99104 96955 99106
rect 94668 99048 96894 99104
rect 96950 99048 96955 99104
rect 94668 99046 96955 99048
rect 96889 99043 96955 99046
rect 66805 98834 66871 98837
rect 226333 98834 226399 98837
rect 226977 98834 227043 98837
rect 66805 98832 68908 98834
rect 66805 98776 66810 98832
rect 66866 98776 68908 98832
rect 224940 98832 227043 98834
rect 66805 98774 68908 98776
rect 66805 98771 66871 98774
rect 97349 98290 97415 98293
rect 94668 98288 97415 98290
rect 94668 98232 97354 98288
rect 97410 98232 97415 98288
rect 94668 98230 97415 98232
rect 97349 98227 97415 98230
rect 151169 98290 151235 98293
rect 193630 98290 193690 98804
rect 224940 98776 226338 98832
rect 226394 98776 226982 98832
rect 227038 98776 227043 98832
rect 224940 98774 227043 98776
rect 226333 98771 226399 98774
rect 226977 98771 227043 98774
rect 227897 98698 227963 98701
rect 237373 98698 237439 98701
rect 227897 98696 237439 98698
rect 227897 98640 227902 98696
rect 227958 98640 237378 98696
rect 237434 98640 237439 98696
rect 227897 98638 237439 98640
rect 227897 98635 227963 98638
rect 237373 98635 237439 98638
rect 151169 98288 193690 98290
rect 151169 98232 151174 98288
rect 151230 98232 193690 98288
rect 151169 98230 193690 98232
rect 151169 98227 151235 98230
rect 66662 97956 66668 98020
rect 66732 98018 66738 98020
rect 67541 98018 67607 98021
rect 191649 98018 191715 98021
rect 227897 98018 227963 98021
rect 66732 98016 68908 98018
rect 66732 97960 67546 98016
rect 67602 97960 68908 98016
rect 66732 97958 68908 97960
rect 191649 98016 193660 98018
rect 191649 97960 191654 98016
rect 191710 97960 193660 98016
rect 191649 97958 193660 97960
rect 224940 98016 227963 98018
rect 224940 97960 227902 98016
rect 227958 97960 227963 98016
rect 224940 97958 227963 97960
rect 66732 97956 66738 97958
rect 67541 97955 67607 97958
rect 191649 97955 191715 97958
rect 227897 97955 227963 97958
rect -960 97610 480 97700
rect 3049 97610 3115 97613
rect -960 97608 3115 97610
rect -960 97552 3054 97608
rect 3110 97552 3115 97608
rect -960 97550 3115 97552
rect -960 97460 480 97550
rect 3049 97547 3115 97550
rect 97901 97474 97967 97477
rect 94668 97472 97967 97474
rect 94668 97416 97906 97472
rect 97962 97416 97967 97472
rect 94668 97414 97967 97416
rect 97901 97411 97967 97414
rect 224718 97412 224724 97476
rect 224788 97474 224794 97476
rect 270493 97474 270559 97477
rect 224788 97472 270559 97474
rect 224788 97416 270498 97472
rect 270554 97416 270559 97472
rect 224788 97414 270559 97416
rect 224788 97412 224794 97414
rect 270493 97411 270559 97414
rect 67449 97202 67515 97205
rect 190637 97202 190703 97205
rect 225137 97202 225203 97205
rect 67449 97200 68908 97202
rect 67449 97144 67454 97200
rect 67510 97144 68908 97200
rect 67449 97142 68908 97144
rect 190637 97200 193660 97202
rect 190637 97144 190642 97200
rect 190698 97144 193660 97200
rect 190637 97142 193660 97144
rect 224940 97200 225203 97202
rect 224940 97144 225142 97200
rect 225198 97144 225203 97200
rect 224940 97142 225203 97144
rect 67449 97139 67515 97142
rect 190637 97139 190703 97142
rect 225137 97139 225203 97142
rect 96889 96658 96955 96661
rect 94668 96656 96955 96658
rect 94668 96600 96894 96656
rect 96950 96600 96955 96656
rect 94668 96598 96955 96600
rect 96889 96595 96955 96598
rect 178861 96658 178927 96661
rect 179229 96658 179295 96661
rect 188286 96658 188292 96660
rect 178861 96656 188292 96658
rect 178861 96600 178866 96656
rect 178922 96600 179234 96656
rect 179290 96600 188292 96656
rect 178861 96598 188292 96600
rect 178861 96595 178927 96598
rect 179229 96595 179295 96598
rect 188286 96596 188292 96598
rect 188356 96596 188362 96660
rect 66110 96324 66116 96388
rect 66180 96386 66186 96388
rect 193121 96386 193187 96389
rect 66180 96326 68908 96386
rect 193121 96384 193660 96386
rect 193121 96328 193126 96384
rect 193182 96328 193660 96384
rect 193121 96326 193660 96328
rect 66180 96324 66186 96326
rect 193121 96323 193187 96326
rect 188470 96114 188476 96116
rect 94668 96054 188476 96114
rect 188470 96052 188476 96054
rect 188540 96052 188546 96116
rect 226517 96114 226583 96117
rect 224940 96112 226583 96114
rect 224940 96056 226522 96112
rect 226578 96056 226583 96112
rect 224940 96054 226583 96056
rect 226517 96051 226583 96054
rect 68553 95842 68619 95845
rect 68553 95840 68908 95842
rect 68553 95784 68558 95840
rect 68614 95784 68908 95840
rect 68553 95782 68908 95784
rect 68553 95779 68619 95782
rect 224350 95780 224356 95844
rect 224420 95842 224426 95844
rect 256693 95842 256759 95845
rect 224420 95840 256759 95842
rect 224420 95784 256698 95840
rect 256754 95784 256759 95840
rect 224420 95782 256759 95784
rect 224420 95780 224426 95782
rect 256693 95779 256759 95782
rect 97257 95298 97323 95301
rect 94668 95296 97323 95298
rect 94668 95240 97262 95296
rect 97318 95240 97323 95296
rect 94668 95238 97323 95240
rect 97257 95235 97323 95238
rect 189717 95298 189783 95301
rect 226517 95298 226583 95301
rect 189717 95296 193660 95298
rect 189717 95240 189722 95296
rect 189778 95240 193660 95296
rect 189717 95238 193660 95240
rect 224940 95296 226583 95298
rect 224940 95240 226522 95296
rect 226578 95240 226583 95296
rect 224940 95238 226583 95240
rect 189717 95235 189783 95238
rect 226517 95235 226583 95238
rect 66805 95026 66871 95029
rect 66805 95024 68908 95026
rect 66805 94968 66810 95024
rect 66866 94968 68908 95024
rect 66805 94966 68908 94968
rect 66805 94963 66871 94966
rect 59169 94482 59235 94485
rect 69013 94482 69079 94485
rect 96981 94482 97047 94485
rect 59169 94480 69079 94482
rect 59169 94424 59174 94480
rect 59230 94424 69018 94480
rect 69074 94424 69079 94480
rect 59169 94422 69079 94424
rect 94668 94480 97047 94482
rect 94668 94424 96986 94480
rect 97042 94424 97047 94480
rect 94668 94422 97047 94424
rect 59169 94419 59235 94422
rect 69013 94419 69079 94422
rect 96981 94419 97047 94422
rect 191649 94482 191715 94485
rect 226609 94482 226675 94485
rect 191649 94480 193660 94482
rect 191649 94424 191654 94480
rect 191710 94424 193660 94480
rect 191649 94422 193660 94424
rect 224940 94480 226675 94482
rect 224940 94424 226614 94480
rect 226670 94424 226675 94480
rect 224940 94422 226675 94424
rect 191649 94419 191715 94422
rect 226609 94419 226675 94422
rect 66662 94148 66668 94212
rect 66732 94210 66738 94212
rect 66732 94150 68908 94210
rect 66732 94148 66738 94150
rect 94814 93876 94820 93940
rect 94884 93938 94890 93940
rect 191097 93938 191163 93941
rect 94884 93936 191163 93938
rect 94884 93880 191102 93936
rect 191158 93880 191163 93936
rect 94884 93878 191163 93880
rect 94884 93876 94890 93878
rect 191097 93875 191163 93878
rect 97901 93666 97967 93669
rect 94668 93664 97967 93666
rect 94668 93608 97906 93664
rect 97962 93608 97967 93664
rect 94668 93606 97967 93608
rect 97901 93603 97967 93606
rect 191741 93666 191807 93669
rect 227621 93666 227687 93669
rect 191741 93664 193660 93666
rect 191741 93608 191746 93664
rect 191802 93608 193660 93664
rect 191741 93606 193660 93608
rect 224940 93664 227687 93666
rect 224940 93608 227626 93664
rect 227682 93608 227687 93664
rect 224940 93606 227687 93608
rect 191741 93603 191807 93606
rect 227621 93603 227687 93606
rect 68001 93394 68067 93397
rect 199101 93394 199167 93397
rect 200614 93394 200620 93396
rect 68001 93392 68908 93394
rect 68001 93336 68006 93392
rect 68062 93336 68908 93392
rect 68001 93334 68908 93336
rect 199101 93392 200620 93394
rect 199101 93336 199106 93392
rect 199162 93336 200620 93392
rect 199101 93334 200620 93336
rect 68001 93331 68067 93334
rect 199101 93331 199167 93334
rect 200614 93332 200620 93334
rect 200684 93332 200690 93396
rect 205582 93332 205588 93396
rect 205652 93394 205658 93396
rect 205725 93394 205791 93397
rect 205652 93392 205791 93394
rect 205652 93336 205730 93392
rect 205786 93336 205791 93392
rect 205652 93334 205791 93336
rect 205652 93332 205658 93334
rect 205725 93331 205791 93334
rect 208945 93394 209011 93397
rect 211705 93396 211771 93397
rect 224769 93396 224835 93397
rect 209998 93394 210004 93396
rect 208945 93392 210004 93394
rect 208945 93336 208950 93392
rect 209006 93336 210004 93392
rect 208945 93334 210004 93336
rect 208945 93331 209011 93334
rect 209998 93332 210004 93334
rect 210068 93332 210074 93396
rect 211654 93332 211660 93396
rect 211724 93394 211771 93396
rect 211724 93392 211816 93394
rect 211766 93336 211816 93392
rect 211724 93334 211816 93336
rect 211724 93332 211771 93334
rect 224718 93332 224724 93396
rect 224788 93394 224835 93396
rect 224788 93392 224880 93394
rect 224830 93336 224880 93392
rect 224788 93334 224880 93336
rect 224788 93332 224835 93334
rect 211705 93331 211771 93332
rect 224769 93331 224835 93332
rect 100017 93122 100083 93125
rect 185117 93122 185183 93125
rect 100017 93120 185183 93122
rect 100017 93064 100022 93120
rect 100078 93064 185122 93120
rect 185178 93064 185183 93120
rect 100017 93062 185183 93064
rect 100017 93059 100083 93062
rect 185117 93059 185183 93062
rect 212441 92986 212507 92989
rect 213126 92986 213132 92988
rect 212441 92984 213132 92986
rect 212441 92928 212446 92984
rect 212502 92928 213132 92984
rect 212441 92926 213132 92928
rect 212441 92923 212507 92926
rect 213126 92924 213132 92926
rect 213196 92924 213202 92988
rect 219390 92926 229110 92986
rect 97206 92850 97212 92852
rect 94668 92790 97212 92850
rect 97206 92788 97212 92790
rect 97276 92788 97282 92852
rect 172329 92850 172395 92853
rect 200389 92850 200455 92853
rect 172329 92848 200455 92850
rect 172329 92792 172334 92848
rect 172390 92792 200394 92848
rect 200450 92792 200455 92848
rect 172329 92790 200455 92792
rect 172329 92787 172395 92790
rect 200389 92787 200455 92790
rect 203333 92850 203399 92853
rect 219390 92850 219450 92926
rect 203333 92848 219450 92850
rect 203333 92792 203338 92848
rect 203394 92792 219450 92848
rect 203333 92790 219450 92792
rect 224033 92850 224099 92853
rect 224350 92850 224356 92852
rect 224033 92848 224356 92850
rect 224033 92792 224038 92848
rect 224094 92792 224356 92848
rect 224033 92790 224356 92792
rect 203333 92787 203399 92790
rect 224033 92787 224099 92790
rect 224350 92788 224356 92790
rect 224420 92788 224426 92852
rect 229050 92850 229110 92926
rect 231853 92850 231919 92853
rect 229050 92848 231919 92850
rect 229050 92792 231858 92848
rect 231914 92792 231919 92848
rect 229050 92790 231919 92792
rect 231853 92787 231919 92790
rect 73470 92652 73476 92716
rect 73540 92714 73546 92716
rect 74303 92714 74369 92717
rect 73540 92712 74369 92714
rect 73540 92656 74308 92712
rect 74364 92656 74369 92712
rect 73540 92654 74369 92656
rect 73540 92652 73546 92654
rect 74303 92651 74369 92654
rect 74855 92714 74921 92717
rect 75310 92714 75316 92716
rect 74855 92712 75316 92714
rect 74855 92656 74860 92712
rect 74916 92656 75316 92712
rect 74855 92654 75316 92656
rect 74855 92651 74921 92654
rect 75310 92652 75316 92654
rect 75380 92652 75386 92716
rect 76879 92714 76945 92717
rect 77150 92714 77156 92716
rect 76879 92712 77156 92714
rect 76879 92656 76884 92712
rect 76940 92656 77156 92712
rect 76879 92654 77156 92656
rect 76879 92651 76945 92654
rect 77150 92652 77156 92654
rect 77220 92652 77226 92716
rect 89621 92714 89687 92717
rect 92606 92714 92612 92716
rect 89621 92712 92612 92714
rect 89621 92656 89626 92712
rect 89682 92656 92612 92712
rect 89621 92654 92612 92656
rect 89621 92651 89687 92654
rect 92606 92652 92612 92654
rect 92676 92652 92682 92716
rect 184841 92714 184907 92717
rect 196525 92714 196591 92717
rect 184841 92712 196591 92714
rect 184841 92656 184846 92712
rect 184902 92656 196530 92712
rect 196586 92656 196591 92712
rect 184841 92654 196591 92656
rect 184841 92651 184907 92654
rect 196525 92651 196591 92654
rect 75126 92516 75132 92580
rect 75196 92578 75202 92580
rect 75361 92578 75427 92581
rect 75196 92576 75427 92578
rect 75196 92520 75366 92576
rect 75422 92520 75427 92576
rect 75196 92518 75427 92520
rect 75196 92516 75202 92518
rect 75361 92515 75427 92518
rect 71630 92380 71636 92444
rect 71700 92442 71706 92444
rect 71773 92442 71839 92445
rect 71700 92440 71839 92442
rect 71700 92384 71778 92440
rect 71834 92384 71839 92440
rect 71700 92382 71839 92384
rect 71700 92380 71706 92382
rect 71773 92379 71839 92382
rect 72918 92380 72924 92444
rect 72988 92442 72994 92444
rect 73337 92442 73403 92445
rect 72988 92440 73403 92442
rect 72988 92384 73342 92440
rect 73398 92384 73403 92440
rect 72988 92382 73403 92384
rect 72988 92380 72994 92382
rect 73337 92379 73403 92382
rect 76966 92380 76972 92444
rect 77036 92442 77042 92444
rect 81433 92442 81499 92445
rect 77036 92440 81499 92442
rect 77036 92384 81438 92440
rect 81494 92384 81499 92440
rect 77036 92382 81499 92384
rect 77036 92380 77042 92382
rect 81433 92379 81499 92382
rect 83549 92442 83615 92445
rect 178861 92442 178927 92445
rect 83549 92440 178927 92442
rect 83549 92384 83554 92440
rect 83610 92384 178866 92440
rect 178922 92384 178927 92440
rect 83549 92382 178927 92384
rect 83549 92379 83615 92382
rect 178861 92379 178927 92382
rect 200205 92442 200271 92445
rect 200941 92442 201007 92445
rect 250437 92442 250503 92445
rect 200205 92440 250503 92442
rect 200205 92384 200210 92440
rect 200266 92384 200946 92440
rect 201002 92384 250442 92440
rect 250498 92384 250503 92440
rect 200205 92382 250503 92384
rect 200205 92379 200271 92382
rect 200941 92379 201007 92382
rect 250437 92379 250503 92382
rect 68870 92244 68876 92308
rect 68940 92306 68946 92308
rect 76281 92306 76347 92309
rect 68940 92304 76347 92306
rect 68940 92248 76286 92304
rect 76342 92248 76347 92304
rect 68940 92246 76347 92248
rect 68940 92244 68946 92246
rect 76281 92243 76347 92246
rect 92749 92306 92815 92309
rect 107653 92306 107719 92309
rect 92749 92304 107719 92306
rect 92749 92248 92754 92304
rect 92810 92248 107658 92304
rect 107714 92248 107719 92304
rect 92749 92246 107719 92248
rect 92749 92243 92815 92246
rect 107653 92243 107719 92246
rect 188429 92306 188495 92309
rect 209814 92306 209820 92308
rect 188429 92304 209820 92306
rect 188429 92248 188434 92304
rect 188490 92248 209820 92304
rect 188429 92246 209820 92248
rect 188429 92243 188495 92246
rect 209814 92244 209820 92246
rect 209884 92306 209890 92308
rect 225137 92306 225203 92309
rect 209884 92304 225203 92306
rect 209884 92248 225142 92304
rect 225198 92248 225203 92304
rect 209884 92246 225203 92248
rect 209884 92244 209890 92246
rect 225137 92243 225203 92246
rect 177389 92170 177455 92173
rect 202597 92170 202663 92173
rect 177389 92168 202663 92170
rect 177389 92112 177394 92168
rect 177450 92112 202602 92168
rect 202658 92112 202663 92168
rect 177389 92110 202663 92112
rect 177389 92107 177455 92110
rect 202597 92107 202663 92110
rect 67817 92034 67883 92037
rect 94814 92034 94820 92036
rect 67817 92032 94820 92034
rect 67817 91976 67822 92032
rect 67878 91976 94820 92032
rect 67817 91974 94820 91976
rect 67817 91971 67883 91974
rect 94814 91972 94820 91974
rect 94884 91972 94890 92036
rect 188521 91220 188587 91221
rect 188470 91218 188476 91220
rect 188430 91158 188476 91218
rect 188540 91216 188587 91220
rect 188582 91160 188587 91216
rect 188470 91156 188476 91158
rect 188540 91156 188587 91160
rect 188521 91155 188587 91156
rect 68686 91020 68692 91084
rect 68756 91082 68762 91084
rect 69841 91082 69907 91085
rect 68756 91080 69907 91082
rect 68756 91024 69846 91080
rect 69902 91024 69907 91080
rect 68756 91022 69907 91024
rect 68756 91020 68762 91022
rect 69841 91019 69907 91022
rect 78949 91082 79015 91085
rect 105077 91082 105143 91085
rect 205081 91082 205147 91085
rect 78949 91080 205147 91082
rect 78949 91024 78954 91080
rect 79010 91024 105082 91080
rect 105138 91024 205086 91080
rect 205142 91024 205147 91080
rect 78949 91022 205147 91024
rect 78949 91019 79015 91022
rect 105077 91019 105143 91022
rect 205081 91019 205147 91022
rect 218789 90946 218855 90949
rect 225597 90946 225663 90949
rect 218789 90944 225663 90946
rect 218789 90888 218794 90944
rect 218850 90888 225602 90944
rect 225658 90888 225663 90944
rect 218789 90886 225663 90888
rect 218789 90883 218855 90886
rect 225597 90883 225663 90886
rect 224309 90674 224375 90677
rect 240869 90674 240935 90677
rect 224309 90672 240935 90674
rect 224309 90616 224314 90672
rect 224370 90616 240874 90672
rect 240930 90616 240935 90672
rect 224309 90614 240935 90616
rect 224309 90611 224375 90614
rect 240869 90611 240935 90614
rect 106038 90476 106044 90540
rect 106108 90538 106114 90540
rect 203701 90538 203767 90541
rect 106108 90536 203767 90538
rect 106108 90480 203706 90536
rect 203762 90480 203767 90536
rect 106108 90478 203767 90480
rect 106108 90476 106114 90478
rect 203701 90475 203767 90478
rect 94078 90340 94084 90404
rect 94148 90402 94154 90404
rect 94497 90402 94563 90405
rect 94148 90400 94563 90402
rect 94148 90344 94502 90400
rect 94558 90344 94563 90400
rect 94148 90342 94563 90344
rect 94148 90340 94154 90342
rect 94497 90339 94563 90342
rect 104157 90402 104223 90405
rect 104525 90402 104591 90405
rect 204437 90402 204503 90405
rect 104157 90400 204503 90402
rect 104157 90344 104162 90400
rect 104218 90344 104530 90400
rect 104586 90344 204442 90400
rect 204498 90344 204503 90400
rect 104157 90342 204503 90344
rect 104157 90339 104223 90342
rect 104525 90339 104591 90342
rect 204437 90339 204503 90342
rect 215293 90268 215359 90269
rect 215293 90266 215340 90268
rect 215212 90264 215340 90266
rect 215404 90266 215410 90268
rect 216397 90266 216463 90269
rect 215404 90264 216463 90266
rect 215212 90208 215298 90264
rect 215404 90208 216402 90264
rect 216458 90208 216463 90264
rect 215212 90206 215340 90208
rect 215293 90204 215340 90206
rect 215404 90206 216463 90208
rect 215404 90204 215410 90206
rect 215293 90203 215359 90204
rect 216397 90203 216463 90206
rect 105629 89858 105695 89861
rect 106038 89858 106044 89860
rect 105629 89856 106044 89858
rect 105629 89800 105634 89856
rect 105690 89800 106044 89856
rect 105629 89798 106044 89800
rect 105629 89795 105695 89798
rect 106038 89796 106044 89798
rect 106108 89796 106114 89860
rect 78397 89722 78463 89725
rect 111149 89722 111215 89725
rect 204989 89722 205055 89725
rect 78397 89720 205055 89722
rect 78397 89664 78402 89720
rect 78458 89664 111154 89720
rect 111210 89664 204994 89720
rect 205050 89664 205055 89720
rect 78397 89662 205055 89664
rect 78397 89659 78463 89662
rect 111149 89659 111215 89662
rect 204989 89659 205055 89662
rect 68369 89586 68435 89589
rect 95417 89586 95483 89589
rect 68369 89584 95483 89586
rect 68369 89528 68374 89584
rect 68430 89528 95422 89584
rect 95478 89528 95483 89584
rect 68369 89526 95483 89528
rect 68369 89523 68435 89526
rect 95417 89523 95483 89526
rect 189809 89586 189875 89589
rect 227897 89586 227963 89589
rect 189809 89584 227963 89586
rect 189809 89528 189814 89584
rect 189870 89528 227902 89584
rect 227958 89528 227963 89584
rect 189809 89526 227963 89528
rect 189809 89523 189875 89526
rect 227897 89523 227963 89526
rect 78029 89450 78095 89453
rect 104525 89450 104591 89453
rect 78029 89448 104591 89450
rect 78029 89392 78034 89448
rect 78090 89392 104530 89448
rect 104586 89392 104591 89448
rect 78029 89390 104591 89392
rect 78029 89387 78095 89390
rect 104525 89387 104591 89390
rect 188286 89388 188292 89452
rect 188356 89450 188362 89452
rect 210509 89450 210575 89453
rect 211061 89450 211127 89453
rect 188356 89448 211127 89450
rect 188356 89392 210514 89448
rect 210570 89392 211066 89448
rect 211122 89392 211127 89448
rect 188356 89390 211127 89392
rect 188356 89388 188362 89390
rect 210509 89387 210575 89390
rect 211061 89387 211127 89390
rect 196065 88226 196131 88229
rect 226517 88226 226583 88229
rect 196065 88224 226583 88226
rect 196065 88168 196070 88224
rect 196126 88168 226522 88224
rect 226578 88168 226583 88224
rect 196065 88166 226583 88168
rect 196065 88163 196131 88166
rect 226517 88163 226583 88166
rect 82077 88090 82143 88093
rect 109033 88090 109099 88093
rect 209221 88090 209287 88093
rect 82077 88088 209287 88090
rect 82077 88032 82082 88088
rect 82138 88032 109038 88088
rect 109094 88032 209226 88088
rect 209282 88032 209287 88088
rect 82077 88030 209287 88032
rect 82077 88027 82143 88030
rect 109033 88027 109099 88030
rect 209221 88027 209287 88030
rect 71773 87954 71839 87957
rect 197077 87954 197143 87957
rect 71773 87952 197143 87954
rect 71773 87896 71778 87952
rect 71834 87896 197082 87952
rect 197138 87896 197143 87952
rect 71773 87894 197143 87896
rect 71773 87891 71839 87894
rect 197077 87891 197143 87894
rect 192702 87484 192708 87548
rect 192772 87546 192778 87548
rect 338113 87546 338179 87549
rect 192772 87544 338179 87546
rect 192772 87488 338118 87544
rect 338174 87488 338179 87544
rect 192772 87486 338179 87488
rect 192772 87484 192778 87486
rect 338113 87483 338179 87486
rect 82997 86866 83063 86869
rect 180057 86866 180123 86869
rect 204437 86866 204503 86869
rect 277393 86866 277459 86869
rect 278681 86866 278747 86869
rect 82997 86864 180810 86866
rect 82997 86808 83002 86864
rect 83058 86808 180062 86864
rect 180118 86808 180810 86864
rect 82997 86806 180810 86808
rect 82997 86803 83063 86806
rect 180057 86803 180123 86806
rect 67541 86730 67607 86733
rect 151169 86730 151235 86733
rect 67541 86728 151235 86730
rect 67541 86672 67546 86728
rect 67602 86672 151174 86728
rect 151230 86672 151235 86728
rect 67541 86670 151235 86672
rect 180750 86730 180810 86806
rect 204437 86864 278747 86866
rect 204437 86808 204442 86864
rect 204498 86808 277398 86864
rect 277454 86808 278686 86864
rect 278742 86808 278747 86864
rect 204437 86806 278747 86808
rect 204437 86803 204503 86806
rect 277393 86803 277459 86806
rect 278681 86803 278747 86806
rect 210325 86730 210391 86733
rect 180750 86728 210391 86730
rect 180750 86672 210330 86728
rect 210386 86672 210391 86728
rect 180750 86670 210391 86672
rect 67541 86667 67607 86670
rect 151169 86667 151235 86670
rect 210325 86667 210391 86670
rect 70853 86594 70919 86597
rect 100109 86594 100175 86597
rect 70853 86592 100175 86594
rect 70853 86536 70858 86592
rect 70914 86536 100114 86592
rect 100170 86536 100175 86592
rect 70853 86534 100175 86536
rect 70853 86531 70919 86534
rect 100109 86531 100175 86534
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 278681 85642 278747 85645
rect 583526 85642 583586 85990
rect 278681 85640 583586 85642
rect 278681 85584 278686 85640
rect 278742 85584 583586 85640
rect 278681 85582 583586 85584
rect 278681 85579 278747 85582
rect 194685 85506 194751 85509
rect 195881 85506 195947 85509
rect 237649 85506 237715 85509
rect 238477 85506 238543 85509
rect 180750 85504 195947 85506
rect 180750 85448 194690 85504
rect 194746 85448 195886 85504
rect 195942 85448 195947 85504
rect 180750 85446 195947 85448
rect 69841 85370 69907 85373
rect 180750 85370 180810 85446
rect 194685 85443 194751 85446
rect 195881 85443 195947 85446
rect 200070 85504 238543 85506
rect 200070 85448 237654 85504
rect 237710 85448 238482 85504
rect 238538 85448 238543 85504
rect 200070 85446 238543 85448
rect 69841 85368 180810 85370
rect 69841 85312 69846 85368
rect 69902 85312 180810 85368
rect 69841 85310 180810 85312
rect 191097 85370 191163 85373
rect 200070 85370 200130 85446
rect 237649 85443 237715 85446
rect 238477 85443 238543 85446
rect 191097 85368 200130 85370
rect 191097 85312 191102 85368
rect 191158 85312 200130 85368
rect 191097 85310 200130 85312
rect 210233 85370 210299 85373
rect 231301 85370 231367 85373
rect 210233 85368 231367 85370
rect 210233 85312 210238 85368
rect 210294 85312 231306 85368
rect 231362 85312 231367 85368
rect 210233 85310 231367 85312
rect 69841 85307 69907 85310
rect 191097 85307 191163 85310
rect 210233 85307 210299 85310
rect 231301 85307 231367 85310
rect 90357 84826 90423 84829
rect 96797 84826 96863 84829
rect 90357 84824 96863 84826
rect -960 84690 480 84780
rect 90357 84768 90362 84824
rect 90418 84768 96802 84824
rect 96858 84768 96863 84824
rect 90357 84766 96863 84768
rect 90357 84763 90423 84766
rect 96797 84763 96863 84766
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 187049 84146 187115 84149
rect 226374 84146 226380 84148
rect 187049 84144 226380 84146
rect 187049 84088 187054 84144
rect 187110 84088 226380 84144
rect 187049 84086 226380 84088
rect 187049 84083 187115 84086
rect 226374 84084 226380 84086
rect 226444 84084 226450 84148
rect 85665 84010 85731 84013
rect 116025 84010 116091 84013
rect 85665 84008 116091 84010
rect 85665 83952 85670 84008
rect 85726 83952 116030 84008
rect 116086 83952 116091 84008
rect 85665 83950 116091 83952
rect 85665 83947 85731 83950
rect 116025 83947 116091 83950
rect 91461 83874 91527 83877
rect 104985 83874 105051 83877
rect 91461 83872 105051 83874
rect 91461 83816 91466 83872
rect 91522 83816 104990 83872
rect 105046 83816 105051 83872
rect 91461 83814 105051 83816
rect 91461 83811 91527 83814
rect 104985 83811 105051 83814
rect 64781 83738 64847 83741
rect 189073 83738 189139 83741
rect 64781 83736 189139 83738
rect 64781 83680 64786 83736
rect 64842 83680 189078 83736
rect 189134 83680 189139 83736
rect 64781 83678 189139 83680
rect 64781 83675 64847 83678
rect 189073 83675 189139 83678
rect 191557 83466 191623 83469
rect 228357 83466 228423 83469
rect 191557 83464 228423 83466
rect 191557 83408 191562 83464
rect 191618 83408 228362 83464
rect 228418 83408 228423 83464
rect 191557 83406 228423 83408
rect 191557 83403 191623 83406
rect 228357 83403 228423 83406
rect 189073 82922 189139 82925
rect 189717 82922 189783 82925
rect 189073 82920 189783 82922
rect 189073 82864 189078 82920
rect 189134 82864 189722 82920
rect 189778 82864 189783 82920
rect 189073 82862 189783 82864
rect 189073 82859 189139 82862
rect 189717 82859 189783 82862
rect 63401 82786 63467 82789
rect 98637 82786 98703 82789
rect 63401 82784 98703 82786
rect 63401 82728 63406 82784
rect 63462 82728 98642 82784
rect 98698 82728 98703 82784
rect 63401 82726 98703 82728
rect 63401 82723 63467 82726
rect 98637 82723 98703 82726
rect 98913 82786 98979 82789
rect 226333 82786 226399 82789
rect 98913 82784 226399 82786
rect 98913 82728 98918 82784
rect 98974 82728 226338 82784
rect 226394 82728 226399 82784
rect 98913 82726 226399 82728
rect 98913 82723 98979 82726
rect 226333 82723 226399 82726
rect 69013 82106 69079 82109
rect 182766 82106 182772 82108
rect 69013 82104 182772 82106
rect 69013 82048 69018 82104
rect 69074 82048 182772 82104
rect 69013 82046 182772 82048
rect 69013 82043 69079 82046
rect 182766 82044 182772 82046
rect 182836 82044 182842 82108
rect 212441 82106 212507 82109
rect 353293 82106 353359 82109
rect 212441 82104 353359 82106
rect 212441 82048 212446 82104
rect 212502 82048 353298 82104
rect 353354 82048 353359 82104
rect 212441 82046 353359 82048
rect 212441 82043 212507 82046
rect 353293 82043 353359 82046
rect 91093 81426 91159 81429
rect 187550 81426 187556 81428
rect 91093 81424 187556 81426
rect 91093 81368 91098 81424
rect 91154 81368 187556 81424
rect 91093 81366 187556 81368
rect 91093 81363 91159 81366
rect 187550 81364 187556 81366
rect 187620 81426 187626 81428
rect 219617 81426 219683 81429
rect 187620 81424 219683 81426
rect 187620 81368 219622 81424
rect 219678 81368 219683 81424
rect 187620 81366 219683 81368
rect 187620 81364 187626 81366
rect 219617 81363 219683 81366
rect 193806 80684 193812 80748
rect 193876 80746 193882 80748
rect 273253 80746 273319 80749
rect 193876 80744 273319 80746
rect 193876 80688 273258 80744
rect 273314 80688 273319 80744
rect 193876 80686 273319 80688
rect 193876 80684 193882 80686
rect 273253 80683 273319 80686
rect 77293 80066 77359 80069
rect 105629 80066 105695 80069
rect 77293 80064 105695 80066
rect 77293 80008 77298 80064
rect 77354 80008 105634 80064
rect 105690 80008 105695 80064
rect 77293 80006 105695 80008
rect 77293 80003 77359 80006
rect 105629 80003 105695 80006
rect 196566 79460 196572 79524
rect 196636 79522 196642 79524
rect 262213 79522 262279 79525
rect 196636 79520 262279 79522
rect 196636 79464 262218 79520
rect 262274 79464 262279 79520
rect 196636 79462 262279 79464
rect 196636 79460 196642 79462
rect 262213 79459 262279 79462
rect 205541 79386 205607 79389
rect 288433 79386 288499 79389
rect 205541 79384 288499 79386
rect 205541 79328 205546 79384
rect 205602 79328 288438 79384
rect 288494 79328 288499 79384
rect 205541 79326 288499 79328
rect 205541 79323 205607 79326
rect 288433 79323 288499 79326
rect 185577 78706 185643 78709
rect 186221 78706 186287 78709
rect 205541 78706 205607 78709
rect 185577 78704 205607 78706
rect 185577 78648 185582 78704
rect 185638 78648 186226 78704
rect 186282 78648 205546 78704
rect 205602 78648 205607 78704
rect 185577 78646 205607 78648
rect 185577 78643 185643 78646
rect 186221 78643 186287 78646
rect 205541 78643 205607 78646
rect 195881 78570 195947 78573
rect 287145 78570 287211 78573
rect 288341 78570 288407 78573
rect 195881 78568 288407 78570
rect 195881 78512 195886 78568
rect 195942 78512 287150 78568
rect 287206 78512 288346 78568
rect 288402 78512 288407 78568
rect 195881 78510 288407 78512
rect 195881 78507 195947 78510
rect 287145 78507 287211 78510
rect 288341 78507 288407 78510
rect 52545 77890 52611 77893
rect 181437 77890 181503 77893
rect 52545 77888 181503 77890
rect 52545 77832 52550 77888
rect 52606 77832 181442 77888
rect 181498 77832 181503 77888
rect 52545 77830 181503 77832
rect 52545 77827 52611 77830
rect 181437 77827 181503 77830
rect 191097 77210 191163 77213
rect 191649 77210 191715 77213
rect 278773 77210 278839 77213
rect 280061 77210 280127 77213
rect 191097 77208 280127 77210
rect 191097 77152 191102 77208
rect 191158 77152 191654 77208
rect 191710 77152 278778 77208
rect 278834 77152 280066 77208
rect 280122 77152 280127 77208
rect 191097 77150 280127 77152
rect 191097 77147 191163 77150
rect 191649 77147 191715 77150
rect 278773 77147 278839 77150
rect 280061 77147 280127 77150
rect 70393 76530 70459 76533
rect 176653 76530 176719 76533
rect 70393 76528 176719 76530
rect 70393 76472 70398 76528
rect 70454 76472 176658 76528
rect 176714 76472 176719 76528
rect 70393 76470 176719 76472
rect 70393 76467 70459 76470
rect 176653 76467 176719 76470
rect 89897 75850 89963 75853
rect 220077 75850 220143 75853
rect 89897 75848 220143 75850
rect 89897 75792 89902 75848
rect 89958 75792 220082 75848
rect 220138 75792 220143 75848
rect 89897 75790 220143 75792
rect 89897 75787 89963 75790
rect 220077 75787 220143 75790
rect 184054 74428 184060 74492
rect 184124 74490 184130 74492
rect 284937 74490 285003 74493
rect 184124 74488 285003 74490
rect 184124 74432 284942 74488
rect 284998 74432 285003 74488
rect 184124 74430 285003 74432
rect 184124 74428 184130 74430
rect 284937 74427 285003 74430
rect 284293 73266 284359 73269
rect 284937 73266 285003 73269
rect 284293 73264 285003 73266
rect 284293 73208 284298 73264
rect 284354 73208 284942 73264
rect 284998 73208 285003 73264
rect 284293 73206 285003 73208
rect 284293 73203 284359 73206
rect 284937 73203 285003 73206
rect 580257 72994 580323 72997
rect 583520 72994 584960 73084
rect 580257 72992 584960 72994
rect 580257 72936 580262 72992
rect 580318 72936 584960 72992
rect 580257 72934 584960 72936
rect 580257 72931 580323 72934
rect 583520 72844 584960 72934
rect 74441 71770 74507 71773
rect 200757 71770 200823 71773
rect 74441 71768 200823 71770
rect -960 71634 480 71724
rect 74441 71712 74446 71768
rect 74502 71712 200762 71768
rect 200818 71712 200823 71768
rect 74441 71710 200823 71712
rect 74441 71707 74507 71710
rect 200757 71707 200823 71710
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 176561 65514 176627 65517
rect 335353 65514 335419 65517
rect 176561 65512 335419 65514
rect 176561 65456 176566 65512
rect 176622 65456 335358 65512
rect 335414 65456 335419 65512
rect 176561 65454 335419 65456
rect 176561 65451 176627 65454
rect 335353 65451 335419 65454
rect 121545 62794 121611 62797
rect 215201 62794 215267 62797
rect 121545 62792 215267 62794
rect 121545 62736 121550 62792
rect 121606 62736 215206 62792
rect 215262 62736 215267 62792
rect 121545 62734 215267 62736
rect 121545 62731 121611 62734
rect 215201 62731 215267 62734
rect 66662 62052 66668 62116
rect 66732 62114 66738 62116
rect 191097 62114 191163 62117
rect 66732 62112 191163 62114
rect 66732 62056 191102 62112
rect 191158 62056 191163 62112
rect 66732 62054 191163 62056
rect 66732 62052 66738 62054
rect 191097 62051 191163 62054
rect 68001 60618 68067 60621
rect 183553 60618 183619 60621
rect 184289 60618 184355 60621
rect 68001 60616 184355 60618
rect 68001 60560 68006 60616
rect 68062 60560 183558 60616
rect 183614 60560 184294 60616
rect 184350 60560 184355 60616
rect 68001 60558 184355 60560
rect 68001 60555 68067 60558
rect 183553 60555 183619 60558
rect 184289 60555 184355 60558
rect 582741 59666 582807 59669
rect 583520 59666 584960 59756
rect 582741 59664 584960 59666
rect 582741 59608 582746 59664
rect 582802 59608 584960 59664
rect 582741 59606 584960 59608
rect 582741 59603 582807 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 60733 46202 60799 46205
rect 173934 46202 173940 46204
rect 60733 46200 173940 46202
rect 60733 46144 60738 46200
rect 60794 46144 173940 46200
rect 60733 46142 173940 46144
rect 60733 46139 60799 46142
rect 173934 46140 173940 46142
rect 174004 46140 174010 46204
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 56593 40626 56659 40629
rect 175774 40626 175780 40628
rect 56593 40624 175780 40626
rect 56593 40568 56598 40624
rect 56654 40568 175780 40624
rect 56593 40566 175780 40568
rect 56593 40563 56659 40566
rect 175774 40564 175780 40566
rect 175844 40564 175850 40628
rect 208158 39204 208164 39268
rect 208228 39266 208234 39268
rect 299565 39266 299631 39269
rect 208228 39264 299631 39266
rect 208228 39208 299570 39264
rect 299626 39208 299631 39264
rect 208228 39206 299631 39208
rect 208228 39204 208234 39206
rect 299565 39203 299631 39206
rect 582925 33146 582991 33149
rect 583520 33146 584960 33236
rect 582925 33144 584960 33146
rect 582925 33088 582930 33144
rect 582986 33088 584960 33144
rect 582925 33086 584960 33088
rect 582925 33083 582991 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 103513 30970 103579 30973
rect 141366 30970 141372 30972
rect 103513 30968 141372 30970
rect 103513 30912 103518 30968
rect 103574 30912 141372 30968
rect 103513 30910 141372 30912
rect 103513 30907 103579 30910
rect 141366 30908 141372 30910
rect 141436 30908 141442 30972
rect 197854 26828 197860 26892
rect 197924 26890 197930 26892
rect 300853 26890 300919 26893
rect 197924 26888 300919 26890
rect 197924 26832 300858 26888
rect 300914 26832 300919 26888
rect 197924 26830 300919 26832
rect 197924 26828 197930 26830
rect 300853 26827 300919 26830
rect 11145 25530 11211 25533
rect 159214 25530 159220 25532
rect 11145 25528 159220 25530
rect 11145 25472 11150 25528
rect 11206 25472 159220 25528
rect 11145 25470 159220 25472
rect 11145 25467 11211 25470
rect 159214 25468 159220 25470
rect 159284 25468 159290 25532
rect 203190 21252 203196 21316
rect 203260 21314 203266 21316
rect 302969 21314 303035 21317
rect 203260 21312 303035 21314
rect 203260 21256 302974 21312
rect 303030 21256 303035 21312
rect 203260 21254 303035 21256
rect 203260 21252 203266 21254
rect 302969 21251 303035 21254
rect 582649 19818 582715 19821
rect 583520 19818 584960 19908
rect 582649 19816 584960 19818
rect 582649 19760 582654 19816
rect 582710 19760 584960 19816
rect 582649 19758 584960 19760
rect 582649 19755 582715 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 582833 6626 582899 6629
rect 583520 6626 584960 6716
rect 582833 6624 584960 6626
rect -960 6490 480 6580
rect 582833 6568 582838 6624
rect 582894 6568 584960 6624
rect 582833 6566 584960 6568
rect 582833 6563 582899 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 304257 4042 304323 4045
rect 307937 4042 308003 4045
rect 304257 4040 308003 4042
rect 304257 3984 304262 4040
rect 304318 3984 307942 4040
rect 307998 3984 308003 4040
rect 304257 3982 308003 3984
rect 304257 3979 304323 3982
rect 307937 3979 308003 3982
rect 101029 3498 101095 3501
rect 101990 3498 101996 3500
rect 101029 3496 101996 3498
rect 101029 3440 101034 3496
rect 101090 3440 101996 3496
rect 101029 3438 101996 3440
rect 101029 3435 101095 3438
rect 101990 3436 101996 3438
rect 102060 3436 102066 3500
rect 147121 3498 147187 3501
rect 147438 3498 147444 3500
rect 147121 3496 147444 3498
rect 147121 3440 147126 3496
rect 147182 3440 147444 3496
rect 147121 3438 147444 3440
rect 147121 3435 147187 3438
rect 147438 3436 147444 3438
rect 147508 3436 147514 3500
rect 269021 3498 269087 3501
rect 274817 3498 274883 3501
rect 269021 3496 274883 3498
rect 269021 3440 269026 3496
rect 269082 3440 274822 3496
rect 274878 3440 274883 3496
rect 269021 3438 274883 3440
rect 269021 3435 269087 3438
rect 274817 3435 274883 3438
rect 341517 3362 341583 3365
rect 350441 3362 350507 3365
rect 341517 3360 350507 3362
rect 341517 3304 341522 3360
rect 341578 3304 350446 3360
rect 350502 3304 350507 3360
rect 341517 3302 350507 3304
rect 341517 3299 341583 3302
rect 350441 3299 350507 3302
<< via3 >>
rect 259500 606052 259564 606116
rect 188292 604556 188356 604620
rect 155724 603196 155788 603260
rect 211660 600748 211724 600812
rect 246252 600748 246316 600812
rect 258396 600612 258460 600676
rect 219940 600476 220004 600540
rect 229692 600476 229756 600540
rect 237972 600476 238036 600540
rect 192340 600340 192404 600404
rect 215340 600400 215404 600404
rect 215340 600344 215354 600400
rect 215354 600344 215404 600400
rect 215340 600340 215404 600344
rect 226932 600340 226996 600404
rect 239260 600340 239324 600404
rect 222700 599116 222764 599180
rect 223804 599116 223868 599180
rect 197124 599040 197188 599044
rect 197124 598984 197174 599040
rect 197174 598984 197188 599040
rect 197124 598980 197188 598984
rect 203196 598980 203260 599044
rect 207060 599040 207124 599044
rect 207060 598984 207110 599040
rect 207110 598984 207124 599040
rect 207060 598980 207124 598984
rect 210372 599040 210436 599044
rect 210372 598984 210422 599040
rect 210422 598984 210436 599040
rect 210372 598980 210436 598984
rect 216444 598980 216508 599044
rect 216628 599040 216692 599044
rect 216628 598984 216678 599040
rect 216678 598984 216692 599040
rect 216628 598980 216692 598984
rect 218652 599040 218716 599044
rect 218652 598984 218702 599040
rect 218702 598984 218716 599040
rect 218652 598980 218716 598984
rect 220860 599040 220924 599044
rect 220860 598984 220910 599040
rect 220910 598984 220924 599040
rect 220860 598980 220924 598984
rect 223988 599040 224052 599044
rect 223988 598984 224038 599040
rect 224038 598984 224052 599040
rect 223988 598980 224052 598984
rect 226196 598980 226260 599044
rect 226380 598980 226444 599044
rect 228220 598980 228284 599044
rect 233004 598980 233068 599044
rect 233188 599040 233252 599044
rect 233188 598984 233238 599040
rect 233238 598984 233252 599040
rect 233188 598980 233252 598984
rect 234660 599040 234724 599044
rect 234660 598984 234710 599040
rect 234710 598984 234724 599040
rect 234660 598980 234724 598984
rect 236500 598980 236564 599044
rect 240732 599040 240796 599044
rect 240732 598984 240746 599040
rect 240746 598984 240796 599040
rect 240732 598980 240796 598984
rect 247724 599040 247788 599044
rect 247724 598984 247774 599040
rect 247774 598984 247788 599040
rect 247724 598980 247788 598984
rect 251036 598980 251100 599044
rect 252508 598980 252572 599044
rect 193260 598436 193324 598500
rect 170996 596804 171060 596868
rect 254532 595172 254596 595236
rect 266308 594900 266372 594964
rect 179276 592724 179340 592788
rect 191604 590684 191668 590748
rect 193260 589868 193324 589932
rect 262260 589324 262324 589388
rect 168236 588100 168300 588164
rect 162716 587964 162780 588028
rect 256740 586468 256804 586532
rect 280292 584020 280356 584084
rect 79916 581224 79980 581228
rect 79916 581168 79966 581224
rect 79966 581168 79980 581224
rect 75684 581028 75748 581092
rect 79916 581164 79980 581168
rect 71636 580756 71700 580820
rect 81020 580756 81084 580820
rect 83964 580756 84028 580820
rect 89300 580816 89364 580820
rect 89300 580760 89314 580816
rect 89314 580760 89364 580816
rect 89300 580756 89364 580760
rect 263548 580212 263612 580276
rect 267780 578308 267844 578372
rect 191604 575452 191668 575516
rect 193444 575452 193508 575516
rect 192340 570692 192404 570756
rect 159956 565796 160020 565860
rect 267964 563348 268028 563412
rect 161244 558996 161308 559060
rect 269068 558996 269132 559060
rect 96660 553420 96724 553484
rect 104940 551924 105004 551988
rect 69244 550836 69308 550900
rect 96660 551244 96724 551308
rect 67772 549476 67836 549540
rect 100708 549340 100772 549404
rect 96844 547028 96908 547092
rect 151676 547028 151740 547092
rect 270540 542676 270604 542740
rect 69428 542132 69492 542196
rect 276244 539684 276308 539748
rect 67772 538732 67836 538796
rect 82860 538732 82924 538796
rect 262444 536012 262508 536076
rect 206140 535468 206204 535532
rect 242940 535468 243004 535532
rect 104204 534652 104268 534716
rect 66116 533292 66180 533356
rect 111748 533292 111812 533356
rect 244412 531932 244476 531996
rect 249012 531252 249076 531316
rect 106780 530708 106844 530772
rect 69796 530572 69860 530636
rect 88932 530572 88996 530636
rect 177804 530572 177868 530636
rect 233004 529076 233068 529140
rect 249748 529076 249812 529140
rect 97028 527716 97092 527780
rect 81020 526764 81084 526828
rect 81020 525812 81084 525876
rect 77156 523636 77220 523700
rect 226196 523636 226260 523700
rect 245700 523636 245764 523700
rect 219940 522276 220004 522340
rect 72740 520916 72804 520980
rect 96844 519420 96908 519484
rect 222700 518060 222764 518124
rect 69612 516700 69676 516764
rect 249012 516700 249076 516764
rect 169340 513300 169404 513364
rect 218652 512620 218716 512684
rect 163636 511260 163700 511324
rect 216628 509764 216692 509828
rect 203196 508404 203260 508468
rect 254716 508404 254780 508468
rect 254532 507860 254596 507924
rect 159772 502964 159836 503028
rect 244780 500108 244844 500172
rect 229692 498748 229756 498812
rect 252508 496028 252572 496092
rect 216444 493444 216508 493508
rect 197124 493308 197188 493372
rect 252508 493308 252572 493372
rect 210372 492764 210436 492828
rect 251036 492628 251100 492692
rect 226932 491812 226996 491876
rect 237972 491132 238036 491196
rect 223804 490588 223868 490652
rect 169524 490452 169588 490516
rect 226380 489228 226444 489292
rect 158484 489092 158548 489156
rect 172100 489092 172164 489156
rect 180196 485828 180260 485892
rect 239260 485012 239324 485076
rect 89300 484332 89364 484396
rect 156644 483652 156708 483716
rect 215340 483652 215404 483716
rect 75684 482156 75748 482220
rect 206140 482156 206204 482220
rect 236500 482156 236564 482220
rect 240732 481536 240796 481540
rect 240732 481480 240782 481536
rect 240782 481480 240796 481536
rect 240732 481476 240796 481480
rect 249012 481476 249076 481540
rect 166212 480796 166276 480860
rect 162532 479436 162596 479500
rect 234660 478076 234724 478140
rect 176516 476716 176580 476780
rect 207060 475356 207124 475420
rect 181484 473996 181548 474060
rect 220860 473996 220924 474060
rect 287100 472092 287164 472156
rect 91324 469780 91388 469844
rect 165476 469780 165540 469844
rect 173756 468556 173820 468620
rect 180012 467740 180076 467804
rect 186820 467196 186884 467260
rect 174676 467060 174740 467124
rect 256556 466652 256620 466716
rect 285628 466576 285692 466580
rect 285628 466520 285678 466576
rect 285678 466520 285692 466576
rect 285628 466516 285692 466520
rect 246252 465972 246316 466036
rect 273484 465020 273548 465084
rect 169340 464340 169404 464404
rect 82676 463524 82740 463588
rect 83964 463524 84028 463588
rect 211660 462844 211724 462908
rect 170812 461484 170876 461548
rect 223988 460260 224052 460324
rect 233188 458900 233252 458964
rect 113220 458764 113284 458828
rect 228220 458764 228284 458828
rect 184796 458220 184860 458284
rect 148916 458084 148980 458148
rect 96844 457404 96908 457468
rect 284340 457404 284404 457468
rect 150940 456860 151004 456924
rect 168972 456180 169036 456244
rect 106780 456044 106844 456108
rect 247724 456044 247788 456108
rect 179092 454684 179156 454748
rect 113036 454064 113100 454068
rect 113036 454008 113050 454064
rect 113050 454008 113100 454064
rect 113036 454004 113100 454008
rect 147444 454004 147508 454068
rect 241652 453868 241716 453932
rect 277164 452644 277228 452708
rect 253980 452100 254044 452164
rect 245884 450256 245948 450260
rect 245884 450200 245934 450256
rect 245934 450200 245948 450256
rect 245884 450196 245948 450200
rect 245700 449652 245764 449716
rect 247724 449652 247788 449716
rect 192708 448624 192772 448628
rect 192708 448568 192758 448624
rect 192758 448568 192772 448624
rect 192708 448564 192772 448568
rect 271092 447748 271156 447812
rect 188844 447340 188908 447404
rect 188292 446388 188356 446452
rect 253980 446116 254044 446180
rect 66668 444892 66732 444956
rect 69428 440812 69492 440876
rect 254532 440404 254596 440468
rect 68140 439452 68204 439516
rect 70716 438908 70780 438972
rect 71636 438908 71700 438972
rect 256556 437548 256620 437612
rect 73476 436324 73540 436388
rect 78260 436188 78324 436252
rect 102732 436188 102796 436252
rect 79732 436052 79796 436116
rect 84700 436052 84764 436116
rect 94452 436052 94516 436116
rect 67404 434556 67468 434620
rect 83044 434420 83108 434484
rect 69060 434284 69124 434348
rect 80100 434284 80164 434348
rect 84516 434344 84580 434348
rect 84516 434288 84566 434344
rect 84566 434288 84580 434344
rect 84516 434284 84580 434288
rect 85804 434344 85868 434348
rect 85804 434288 85854 434344
rect 85854 434288 85868 434344
rect 85804 434284 85868 434288
rect 95188 434284 95252 434348
rect 100156 434344 100220 434348
rect 100156 434288 100206 434344
rect 100206 434288 100220 434344
rect 100156 434284 100220 434288
rect 92612 434208 92676 434212
rect 92612 434152 92662 434208
rect 92662 434152 92676 434208
rect 92612 434148 92676 434152
rect 67404 433876 67468 433940
rect 74948 433740 75012 433804
rect 98500 433740 98564 433804
rect 70716 433664 70780 433668
rect 70716 433608 70730 433664
rect 70730 433608 70780 433664
rect 70716 433604 70780 433608
rect 73660 433604 73724 433668
rect 74764 433664 74828 433668
rect 74764 433608 74814 433664
rect 74814 433608 74828 433664
rect 74764 433604 74828 433608
rect 76052 433604 76116 433668
rect 78444 433604 78508 433668
rect 86724 433604 86788 433668
rect 87092 433604 87156 433668
rect 87460 433604 87524 433668
rect 89668 433664 89732 433668
rect 89668 433608 89682 433664
rect 89682 433608 89732 433664
rect 89668 433604 89732 433608
rect 90036 433664 90100 433668
rect 90036 433608 90086 433664
rect 90086 433608 90100 433664
rect 90036 433604 90100 433608
rect 91508 433664 91572 433668
rect 91508 433608 91558 433664
rect 91558 433608 91572 433664
rect 91508 433604 91572 433608
rect 92796 433604 92860 433668
rect 97948 433604 98012 433668
rect 99972 433604 100036 433668
rect 100892 433664 100956 433668
rect 100892 433608 100942 433664
rect 100942 433608 100956 433664
rect 100892 433604 100956 433608
rect 105124 433664 105188 433668
rect 105124 433608 105174 433664
rect 105174 433608 105188 433664
rect 105124 433604 105188 433608
rect 106412 433604 106476 433668
rect 109540 433664 109604 433668
rect 109540 433608 109554 433664
rect 109554 433608 109604 433664
rect 109540 433604 109604 433608
rect 111012 433604 111076 433668
rect 180196 430612 180260 430676
rect 114508 430068 114572 430132
rect 68140 429388 68204 429452
rect 161060 428436 161124 428500
rect 69428 427620 69492 427684
rect 67404 425172 67468 425236
rect 159772 418780 159836 418844
rect 166396 418780 166460 418844
rect 150940 418236 151004 418300
rect 180564 417480 180628 417484
rect 180564 417424 180578 417480
rect 180578 417424 180628 417480
rect 180564 417420 180628 417424
rect 281580 416604 281644 416668
rect 159772 414564 159836 414628
rect 114692 413748 114756 413812
rect 179276 413204 179340 413268
rect 252876 404772 252940 404836
rect 112116 402596 112180 402660
rect 112116 398924 112180 398988
rect 113036 398924 113100 398988
rect 177804 398788 177868 398852
rect 66668 397428 66732 397492
rect 253060 397292 253124 397356
rect 253980 396884 254044 396948
rect 113220 396340 113284 396404
rect 66668 395252 66732 395316
rect 254532 394572 254596 394636
rect 69428 393892 69492 393956
rect 254716 392532 254780 392596
rect 253980 392048 254044 392052
rect 253980 391992 254030 392048
rect 254030 391992 254044 392048
rect 253980 391988 254044 391992
rect 82308 391852 82372 391916
rect 82676 391852 82740 391916
rect 82308 390900 82372 390964
rect 84516 390900 84580 390964
rect 114692 391444 114756 391508
rect 107516 390900 107580 390964
rect 91324 390764 91388 390828
rect 96844 390824 96908 390828
rect 96844 390768 96858 390824
rect 96858 390768 96908 390824
rect 96844 390764 96908 390768
rect 97028 390824 97092 390828
rect 97028 390768 97078 390824
rect 97078 390768 97092 390824
rect 97028 390764 97092 390768
rect 82860 390628 82924 390692
rect 88932 390628 88996 390692
rect 249012 390900 249076 390964
rect 111748 390492 111812 390556
rect 72740 390356 72804 390420
rect 77156 390416 77220 390420
rect 77156 390360 77206 390416
rect 77206 390360 77220 390416
rect 77156 390356 77220 390360
rect 100708 390416 100772 390420
rect 100708 390360 100722 390416
rect 100722 390360 100772 390416
rect 100708 390356 100772 390360
rect 104204 390416 104268 390420
rect 104204 390360 104254 390416
rect 104254 390360 104268 390416
rect 104204 390356 104268 390360
rect 104940 390356 105004 390420
rect 79916 390084 79980 390148
rect 73660 389268 73724 389332
rect 244228 388996 244292 389060
rect 78444 388452 78508 388516
rect 251036 388452 251100 388516
rect 254716 388044 254780 388108
rect 100156 387908 100220 387972
rect 84700 387500 84764 387564
rect 78260 386956 78324 387020
rect 87460 386820 87524 386884
rect 170996 386140 171060 386204
rect 100892 385868 100956 385932
rect 66668 385596 66732 385660
rect 271092 385596 271156 385660
rect 85804 385052 85868 385116
rect 187556 384372 187620 384436
rect 80100 382876 80164 382940
rect 94452 382876 94516 382940
rect 114508 382876 114572 382940
rect 102732 382332 102796 382396
rect 180012 382332 180076 382396
rect 187556 382196 187620 382260
rect 248460 381652 248524 381716
rect 280292 380700 280356 380764
rect 273300 378932 273364 378996
rect 192708 378660 192772 378724
rect 288388 377980 288452 378044
rect 69612 377436 69676 377500
rect 241652 377300 241716 377364
rect 276428 376620 276492 376684
rect 111012 370500 111076 370564
rect 181484 370500 181548 370564
rect 77156 369200 77220 369204
rect 77156 369144 77206 369200
rect 77206 369144 77220 369200
rect 77156 369140 77220 369144
rect 252692 366964 252756 367028
rect 258396 366284 258460 366348
rect 247724 364924 247788 364988
rect 270724 364924 270788 364988
rect 262260 363564 262324 363628
rect 71636 362204 71700 362268
rect 256740 362204 256804 362268
rect 245884 359076 245948 359140
rect 273484 356764 273548 356828
rect 259500 356628 259564 356692
rect 280108 355268 280172 355332
rect 162532 351868 162596 351932
rect 169708 351868 169772 351932
rect 263732 351732 263796 351796
rect 179092 351188 179156 351252
rect 244228 351052 244292 351116
rect 262444 349692 262508 349756
rect 267964 345748 268028 345812
rect 254532 345612 254596 345676
rect 269068 344252 269132 344316
rect 173572 341532 173636 341596
rect 163636 341396 163700 341460
rect 268332 341396 268396 341460
rect 160692 339492 160756 339556
rect 161244 339492 161308 339556
rect 173756 337316 173820 337380
rect 245700 337316 245764 337380
rect 156644 336228 156708 336292
rect 141372 336092 141436 336156
rect 156644 335956 156708 336020
rect 158484 334596 158548 334660
rect 242940 334596 243004 334660
rect 267964 334596 268028 334660
rect 267780 334112 267844 334116
rect 267780 334056 267794 334112
rect 267794 334056 267844 334112
rect 267780 334052 267844 334056
rect 159772 333372 159836 333436
rect 258580 333236 258644 333300
rect 263916 330652 263980 330716
rect 166212 330576 166276 330580
rect 166212 330520 166262 330576
rect 166262 330520 166276 330576
rect 166212 330516 166276 330520
rect 252508 330516 252572 330580
rect 172100 330380 172164 330444
rect 263548 330380 263612 330444
rect 260972 329156 261036 329220
rect 259500 327252 259564 327316
rect 265756 325756 265820 325820
rect 155172 325076 155236 325140
rect 258580 324940 258644 325004
rect 162716 323580 162780 323644
rect 155724 320724 155788 320788
rect 97764 320180 97828 320244
rect 170812 319364 170876 319428
rect 269068 319364 269132 319428
rect 169524 318820 169588 318884
rect 109540 318004 109604 318068
rect 79732 317460 79796 317524
rect 256740 317324 256804 317388
rect 276244 316644 276308 316708
rect 86724 315964 86788 316028
rect 105124 315284 105188 315348
rect 95188 313924 95252 313988
rect 270540 313924 270604 313988
rect 166764 313380 166828 313444
rect 92796 312428 92860 312492
rect 109540 312428 109604 312492
rect 160692 312020 160756 312084
rect 266308 312020 266372 312084
rect 266492 311340 266556 311404
rect 90036 311068 90100 311132
rect 98500 311068 98564 311132
rect 106412 309708 106476 309772
rect 83044 309028 83108 309092
rect 92612 308348 92676 308412
rect 194732 308076 194796 308140
rect 76052 307804 76116 307868
rect 84516 307668 84580 307732
rect 259684 307124 259748 307188
rect 97948 306988 98012 307052
rect 86724 306444 86788 306508
rect 91508 305764 91572 305828
rect 185348 304948 185412 305012
rect 186820 304948 186884 305012
rect 159220 304268 159284 304332
rect 89668 304132 89732 304196
rect 101260 304132 101324 304196
rect 182772 304132 182836 304196
rect 262444 304132 262508 304196
rect 249748 303724 249812 303788
rect 262260 303588 262324 303652
rect 151676 302772 151740 302836
rect 178540 302500 178604 302564
rect 186268 302560 186332 302564
rect 186268 302504 186282 302560
rect 186282 302504 186332 302560
rect 186268 302500 186332 302504
rect 166948 302364 167012 302428
rect 168236 302364 168300 302428
rect 86540 301548 86604 301612
rect 166948 301548 167012 301612
rect 169156 301412 169220 301476
rect 252692 301548 252756 301612
rect 244780 301004 244844 301068
rect 248460 300732 248524 300796
rect 194732 300052 194796 300116
rect 256740 298692 256804 298756
rect 273116 298148 273180 298212
rect 186820 296924 186884 296988
rect 259684 296652 259748 296716
rect 148916 295156 148980 295220
rect 81940 294612 82004 294676
rect 148916 294476 148980 294540
rect 87092 293116 87156 293180
rect 185348 291892 185412 291956
rect 260972 291620 261036 291684
rect 260972 291212 261036 291276
rect 68876 291076 68940 291140
rect 78444 291076 78508 291140
rect 80652 291076 80716 291140
rect 91508 289988 91572 290052
rect 258580 289988 258644 290052
rect 88012 289580 88076 289644
rect 259500 288764 259564 288828
rect 79180 288628 79244 288692
rect 74764 288492 74828 288556
rect 99972 287812 100036 287876
rect 74948 287132 75012 287196
rect 268332 286044 268396 286108
rect 83412 285636 83476 285700
rect 86724 285636 86788 285700
rect 166764 285636 166828 285700
rect 268332 285772 268396 285836
rect 276244 285772 276308 285836
rect 186268 284956 186332 285020
rect 73476 284140 73540 284204
rect 75684 284140 75748 284204
rect 78260 284140 78324 284204
rect 91140 284140 91204 284204
rect 71820 283460 71884 283524
rect 73292 283520 73356 283524
rect 73292 283464 73306 283520
rect 73306 283464 73356 283520
rect 73292 283460 73356 283464
rect 75316 283460 75380 283524
rect 76972 283460 77036 283524
rect 89852 283520 89916 283524
rect 89852 283464 89866 283520
rect 89866 283464 89916 283520
rect 89852 283460 89916 283464
rect 93348 283460 93412 283524
rect 67588 283324 67652 283388
rect 69060 283188 69124 283252
rect 94084 283324 94148 283388
rect 97764 283324 97828 283388
rect 281764 283596 281828 283660
rect 79916 283052 79980 283116
rect 84700 283052 84764 283116
rect 70164 282916 70228 282980
rect 82676 282976 82740 282980
rect 82676 282920 82690 282976
rect 82690 282920 82740 282976
rect 82676 282916 82740 282920
rect 83412 282976 83476 282980
rect 83412 282920 83462 282976
rect 83462 282920 83476 282976
rect 83412 282916 83476 282920
rect 86724 282916 86788 282980
rect 88748 282916 88812 282980
rect 65932 280468 65996 280532
rect 99972 280196 100036 280260
rect 101260 278564 101324 278628
rect 67588 278080 67652 278084
rect 67588 278024 67602 278080
rect 67602 278024 67652 278080
rect 67588 278020 67652 278024
rect 193812 275300 193876 275364
rect 103836 275164 103900 275228
rect 185348 274620 185412 274684
rect 155172 272444 155236 272508
rect 176516 270404 176580 270468
rect 263732 270404 263796 270468
rect 165476 269724 165540 269788
rect 260972 267004 261036 267068
rect 288388 267004 288452 267068
rect 252876 265916 252940 265980
rect 262444 265508 262508 265572
rect 262444 265100 262508 265164
rect 281580 262788 281644 262852
rect 263916 262712 263980 262716
rect 263916 262656 263930 262712
rect 263930 262656 263980 262712
rect 263916 262652 263980 262656
rect 270724 262380 270788 262444
rect 273668 262108 273732 262172
rect 263548 261428 263612 261492
rect 284340 261428 284404 261492
rect 273668 261156 273732 261220
rect 263548 261020 263612 261084
rect 168972 260476 169036 260540
rect 260972 260476 261036 260540
rect 273300 260204 273364 260268
rect 159956 260068 160020 260132
rect 263732 259932 263796 259996
rect 271092 259388 271156 259452
rect 276428 259388 276492 259452
rect 258396 258844 258460 258908
rect 271092 258300 271156 258364
rect 285628 258164 285692 258228
rect 262444 257212 262508 257276
rect 173940 255988 174004 256052
rect 100708 255716 100772 255780
rect 64644 255308 64708 255372
rect 188844 254084 188908 254148
rect 175780 253948 175844 254012
rect 178540 253948 178604 254012
rect 173572 253812 173636 253876
rect 287100 253812 287164 253876
rect 256740 253676 256804 253740
rect 101260 252452 101324 252516
rect 265940 252452 266004 252516
rect 265756 252044 265820 252108
rect 98132 251228 98196 251292
rect 273116 251092 273180 251156
rect 186820 250412 186884 250476
rect 267964 250064 268028 250068
rect 267964 250008 267978 250064
rect 267978 250008 268028 250064
rect 267964 250004 268028 250008
rect 191788 249052 191852 249116
rect 188292 248508 188356 248572
rect 266492 247692 266556 247756
rect 192340 247420 192404 247484
rect 66668 247012 66732 247076
rect 193444 245788 193508 245852
rect 184796 245652 184860 245716
rect 259500 246332 259564 246396
rect 280292 246332 280356 246396
rect 254532 245652 254596 245716
rect 256740 245652 256804 245716
rect 66852 245516 66916 245580
rect 66116 245380 66180 245444
rect 69428 244292 69492 244356
rect 267780 244156 267844 244220
rect 269620 244156 269684 244220
rect 277164 244156 277228 244220
rect 193260 243476 193324 243540
rect 256740 243340 256804 243404
rect 66852 242932 66916 242996
rect 253612 243204 253676 243268
rect 191788 242856 191852 242860
rect 191788 242800 191838 242856
rect 191838 242800 191852 242856
rect 191788 242796 191852 242800
rect 180564 242116 180628 242180
rect 269068 242252 269132 242316
rect 193260 241980 193324 242044
rect 251036 241980 251100 242044
rect 251772 241980 251836 242044
rect 71636 241708 71700 241772
rect 75684 241708 75748 241772
rect 77156 241708 77220 241772
rect 78076 241708 78140 241772
rect 78444 241768 78508 241772
rect 78444 241712 78458 241768
rect 78458 241712 78508 241768
rect 78444 241708 78508 241712
rect 80652 241708 80716 241772
rect 81940 241768 82004 241772
rect 81940 241712 81990 241768
rect 81990 241712 82004 241768
rect 81940 241708 82004 241712
rect 84516 241708 84580 241772
rect 86540 241768 86604 241772
rect 86540 241712 86590 241768
rect 86590 241712 86604 241768
rect 86540 241708 86604 241712
rect 91140 241708 91204 241772
rect 88012 241572 88076 241636
rect 91508 241572 91572 241636
rect 68876 241436 68940 241500
rect 187556 241436 187620 241500
rect 258396 241436 258460 241500
rect 253612 240892 253676 240956
rect 71636 240076 71700 240140
rect 73476 240076 73540 240140
rect 75132 240076 75196 240140
rect 88012 240076 88076 240140
rect 91140 240136 91204 240140
rect 91140 240080 91154 240136
rect 91154 240080 91204 240136
rect 91140 240076 91204 240080
rect 72924 239940 72988 240004
rect 254532 239668 254596 239732
rect 68876 238852 68940 238916
rect 77156 238580 77220 238644
rect 169708 237280 169772 237284
rect 169708 237224 169758 237280
rect 169758 237224 169772 237280
rect 169708 237220 169772 237224
rect 256740 237220 256804 237284
rect 266308 236676 266372 236740
rect 106044 236540 106108 236604
rect 93900 236404 93964 236468
rect 69612 235724 69676 235788
rect 262260 235180 262324 235244
rect 273484 235180 273548 235244
rect 160140 234500 160204 234564
rect 161060 234500 161124 234564
rect 265756 234500 265820 234564
rect 160140 233820 160204 233884
rect 267964 231780 268028 231844
rect 260972 231100 261036 231164
rect 93900 230420 93964 230484
rect 193812 230420 193876 230484
rect 251772 230012 251836 230076
rect 213132 229876 213196 229940
rect 252692 229876 252756 229940
rect 263732 229740 263796 229804
rect 66668 226204 66732 226268
rect 215340 224164 215404 224228
rect 97948 223484 98012 223548
rect 262444 222124 262508 222188
rect 271092 222124 271156 222188
rect 192340 221988 192404 222052
rect 266492 219268 266556 219332
rect 259500 217228 259564 217292
rect 101260 216684 101324 216748
rect 94084 211788 94148 211852
rect 68876 210972 68940 211036
rect 269620 210836 269684 210900
rect 71636 209612 71700 209676
rect 185348 204988 185412 205052
rect 66116 204852 66180 204916
rect 273668 203492 273732 203556
rect 188292 202132 188356 202196
rect 65932 192476 65996 192540
rect 223620 192476 223684 192540
rect 263548 189620 263612 189684
rect 226380 182820 226444 182884
rect 83412 177244 83476 177308
rect 82676 176700 82740 176764
rect 76972 176564 77036 176628
rect 76972 176156 77036 176220
rect 189948 174524 190012 174588
rect 86724 172348 86788 172412
rect 188292 168948 188356 169012
rect 189948 164324 190012 164388
rect 211660 163372 211724 163436
rect 281764 159292 281828 159356
rect 205588 158068 205652 158132
rect 200620 157932 200684 157996
rect 276244 156572 276308 156636
rect 209820 155892 209884 155956
rect 193996 153852 194060 153916
rect 227668 150996 227732 151060
rect 96292 149228 96356 149292
rect 100708 149228 100772 149292
rect 192340 149092 192404 149156
rect 194548 148276 194612 148340
rect 192340 146236 192404 146300
rect 89852 144740 89916 144804
rect 92612 144740 92676 144804
rect 99972 144740 100036 144804
rect 188292 144800 188356 144804
rect 188292 144744 188342 144800
rect 188342 144744 188356 144800
rect 188292 144740 188356 144744
rect 224356 143652 224420 143716
rect 88748 143516 88812 143580
rect 223620 143516 223684 143580
rect 68692 143380 68756 143444
rect 70164 143244 70228 143308
rect 70164 142972 70228 143036
rect 193260 142896 193324 142900
rect 193260 142840 193310 142896
rect 193310 142840 193324 142896
rect 193260 142836 193324 142840
rect 73292 142292 73356 142356
rect 197860 142156 197924 142220
rect 84700 142020 84764 142084
rect 224908 141068 224972 141132
rect 76972 140796 77036 140860
rect 93348 140796 93412 140860
rect 210004 140524 210068 140588
rect 196572 140388 196636 140452
rect 203196 140388 203260 140452
rect 208164 140448 208228 140452
rect 208164 140392 208214 140448
rect 208214 140392 208228 140448
rect 208164 140388 208228 140392
rect 71820 139572 71884 139636
rect 75316 139300 75380 139364
rect 69428 138620 69492 138684
rect 193260 138620 193324 138684
rect 194180 138756 194244 138820
rect 73292 138212 73356 138276
rect 79916 137260 79980 137324
rect 69244 135084 69308 135148
rect 73476 134812 73540 134876
rect 75316 134676 75380 134740
rect 93716 134676 93780 134740
rect 94084 134676 94148 134740
rect 226380 134676 226444 134740
rect 224356 133316 224420 133380
rect 189948 132500 190012 132564
rect 193812 131412 193876 131476
rect 69428 131004 69492 131068
rect 224356 129644 224420 129708
rect 94636 129508 94700 129572
rect 103836 128420 103900 128484
rect 69244 127060 69308 127124
rect 193444 124068 193508 124132
rect 192708 123796 192772 123860
rect 227668 121076 227732 121140
rect 184060 120668 184124 120732
rect 224908 119988 224972 120052
rect 101996 113732 102060 113796
rect 97212 109516 97276 109580
rect 96292 108836 96356 108900
rect 226380 107748 226444 107812
rect 64644 106252 64708 106316
rect 66668 97956 66732 98020
rect 224724 97412 224788 97476
rect 188292 96596 188356 96660
rect 66116 96324 66180 96388
rect 188476 96052 188540 96116
rect 224356 95780 224420 95844
rect 66668 94148 66732 94212
rect 94820 93876 94884 93940
rect 200620 93332 200684 93396
rect 205588 93332 205652 93396
rect 210004 93332 210068 93396
rect 211660 93392 211724 93396
rect 211660 93336 211710 93392
rect 211710 93336 211724 93392
rect 211660 93332 211724 93336
rect 224724 93392 224788 93396
rect 224724 93336 224774 93392
rect 224774 93336 224788 93392
rect 224724 93332 224788 93336
rect 213132 92924 213196 92988
rect 97212 92788 97276 92852
rect 224356 92788 224420 92852
rect 73476 92652 73540 92716
rect 75316 92652 75380 92716
rect 77156 92652 77220 92716
rect 92612 92652 92676 92716
rect 75132 92516 75196 92580
rect 71636 92380 71700 92444
rect 72924 92380 72988 92444
rect 76972 92380 77036 92444
rect 68876 92244 68940 92308
rect 209820 92244 209884 92308
rect 94820 91972 94884 92036
rect 188476 91216 188540 91220
rect 188476 91160 188526 91216
rect 188526 91160 188540 91216
rect 188476 91156 188540 91160
rect 68692 91020 68756 91084
rect 106044 90476 106108 90540
rect 94084 90340 94148 90404
rect 215340 90264 215404 90268
rect 215340 90208 215354 90264
rect 215354 90208 215404 90264
rect 215340 90204 215404 90208
rect 106044 89796 106108 89860
rect 188292 89388 188356 89452
rect 192708 87484 192772 87548
rect 226380 84084 226444 84148
rect 182772 82044 182836 82108
rect 187556 81364 187620 81428
rect 193812 80684 193876 80748
rect 196572 79460 196636 79524
rect 184060 74428 184124 74492
rect 66668 62052 66732 62116
rect 173940 46140 174004 46204
rect 175780 40564 175844 40628
rect 208164 39204 208228 39268
rect 141372 30908 141436 30972
rect 197860 26828 197924 26892
rect 159220 25468 159284 25532
rect 203196 21252 203260 21316
rect 101996 3436 102060 3500
rect 147444 3436 147508 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 583166 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 583166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 583166 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 583166 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 583166 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 583166 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 79915 581228 79981 581229
rect 79915 581164 79916 581228
rect 79980 581164 79981 581228
rect 79915 581163 79981 581164
rect 75683 581092 75749 581093
rect 75683 581028 75684 581092
rect 75748 581028 75749 581092
rect 75683 581027 75749 581028
rect 71635 580820 71701 580821
rect 71635 580756 71636 580820
rect 71700 580756 71701 580820
rect 71635 580755 71701 580756
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 69243 550900 69309 550901
rect 69243 550836 69244 550900
rect 69308 550836 69309 550900
rect 69243 550835 69309 550836
rect 67771 549540 67837 549541
rect 67771 549476 67772 549540
rect 67836 549476 67837 549540
rect 67771 549475 67837 549476
rect 67774 538797 67834 549475
rect 67771 538796 67837 538797
rect 67771 538732 67772 538796
rect 67836 538732 67837 538796
rect 67771 538731 67837 538732
rect 69246 538250 69306 550835
rect 69427 542196 69493 542197
rect 69427 542132 69428 542196
rect 69492 542132 69493 542196
rect 69427 542131 69493 542132
rect 69430 540970 69490 542131
rect 69430 540910 69858 540970
rect 69246 538190 69674 538250
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66115 533356 66181 533357
rect 66115 533292 66116 533356
rect 66180 533292 66181 533356
rect 66115 533291 66181 533292
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66118 395450 66178 533291
rect 66954 500614 67574 536058
rect 69614 516765 69674 538190
rect 69798 530637 69858 540910
rect 69795 530636 69861 530637
rect 69795 530572 69796 530636
rect 69860 530572 69861 530636
rect 69795 530571 69861 530572
rect 69611 516764 69677 516765
rect 69611 516700 69612 516764
rect 69676 516700 69677 516764
rect 69611 516699 69677 516700
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66667 444956 66733 444957
rect 66667 444892 66668 444956
rect 66732 444892 66733 444956
rect 66667 444891 66733 444892
rect 66670 397493 66730 444891
rect 66954 436356 67574 464058
rect 69427 440876 69493 440877
rect 69427 440812 69428 440876
rect 69492 440812 69493 440876
rect 69427 440811 69493 440812
rect 68139 439516 68205 439517
rect 68139 439452 68140 439516
rect 68204 439452 68205 439516
rect 68139 439451 68205 439452
rect 67403 434620 67469 434621
rect 67403 434556 67404 434620
rect 67468 434556 67469 434620
rect 67403 434555 67469 434556
rect 67406 433941 67466 434555
rect 67403 433940 67469 433941
rect 67403 433876 67404 433940
rect 67468 433876 67469 433940
rect 67403 433875 67469 433876
rect 67406 425237 67466 433875
rect 68142 429453 68202 439451
rect 69059 434348 69125 434349
rect 69059 434284 69060 434348
rect 69124 434284 69125 434348
rect 69059 434283 69125 434284
rect 68139 429452 68205 429453
rect 68139 429388 68140 429452
rect 68204 429388 68205 429452
rect 68139 429387 68205 429388
rect 67403 425236 67469 425237
rect 67403 425172 67404 425236
rect 67468 425172 67469 425236
rect 67403 425171 67469 425172
rect 66667 397492 66733 397493
rect 66667 397428 66668 397492
rect 66732 397428 66733 397492
rect 66667 397427 66733 397428
rect 66118 395390 66730 395450
rect 66670 395317 66730 395390
rect 66667 395316 66733 395317
rect 66667 395252 66668 395316
rect 66732 395252 66733 395316
rect 66667 395251 66733 395252
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 66670 385661 66730 395251
rect 66667 385660 66733 385661
rect 66667 385596 66668 385660
rect 66732 385596 66733 385660
rect 66667 385595 66733 385596
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 66954 356614 67574 388356
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 285592 67574 320058
rect 68875 291140 68941 291141
rect 68875 291076 68876 291140
rect 68940 291076 68941 291140
rect 68875 291075 68941 291076
rect 67587 283388 67653 283389
rect 67587 283324 67588 283388
rect 67652 283324 67653 283388
rect 67587 283323 67653 283324
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 65931 280532 65997 280533
rect 65931 280468 65932 280532
rect 65996 280468 65997 280532
rect 65931 280467 65997 280468
rect 63234 244894 63854 280338
rect 64643 255372 64709 255373
rect 64643 255308 64644 255372
rect 64708 255308 64709 255372
rect 64643 255307 64709 255308
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 64646 106317 64706 255307
rect 65934 192541 65994 280467
rect 67590 278085 67650 283323
rect 67587 278084 67653 278085
rect 67587 278020 67588 278084
rect 67652 278020 67653 278084
rect 67587 278019 67653 278020
rect 66667 247076 66733 247077
rect 66667 247012 66668 247076
rect 66732 247012 66733 247076
rect 66667 247011 66733 247012
rect 66115 245444 66181 245445
rect 66115 245380 66116 245444
rect 66180 245380 66181 245444
rect 66115 245379 66181 245380
rect 66118 204917 66178 245379
rect 66670 226269 66730 247011
rect 66851 245580 66917 245581
rect 66851 245516 66852 245580
rect 66916 245516 66917 245580
rect 66851 245515 66917 245516
rect 66854 242997 66914 245515
rect 66851 242996 66917 242997
rect 66851 242932 66852 242996
rect 66916 242932 66917 242996
rect 66851 242931 66917 242932
rect 68878 241501 68938 291075
rect 69062 283253 69122 434283
rect 69430 427685 69490 440811
rect 71638 438973 71698 580755
rect 73679 543454 73999 543486
rect 73679 543218 73721 543454
rect 73957 543218 73999 543454
rect 73679 543134 73999 543218
rect 73679 542898 73721 543134
rect 73957 542898 73999 543134
rect 73679 542866 73999 542898
rect 72739 520980 72805 520981
rect 72739 520916 72740 520980
rect 72804 520916 72805 520980
rect 72739 520915 72805 520916
rect 70715 438972 70781 438973
rect 70715 438908 70716 438972
rect 70780 438908 70781 438972
rect 70715 438907 70781 438908
rect 71635 438972 71701 438973
rect 71635 438908 71636 438972
rect 71700 438908 71701 438972
rect 71635 438907 71701 438908
rect 70718 433669 70778 438907
rect 70715 433668 70781 433669
rect 70715 433604 70716 433668
rect 70780 433604 70781 433668
rect 70715 433603 70781 433604
rect 69427 427684 69493 427685
rect 69427 427620 69428 427684
rect 69492 427620 69493 427684
rect 69427 427619 69493 427620
rect 69427 393956 69493 393957
rect 69427 393892 69428 393956
rect 69492 393892 69493 393956
rect 69427 393891 69493 393892
rect 69430 393330 69490 393891
rect 69430 393270 69674 393330
rect 69614 377501 69674 393270
rect 72742 390421 72802 520915
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 75686 482221 75746 581027
rect 77644 561454 77964 561486
rect 77644 561218 77686 561454
rect 77922 561218 77964 561454
rect 77644 561134 77964 561218
rect 77644 560898 77686 561134
rect 77922 560898 77964 561134
rect 77644 560866 77964 560898
rect 77155 523700 77221 523701
rect 77155 523636 77156 523700
rect 77220 523636 77221 523700
rect 77155 523635 77221 523636
rect 75683 482220 75749 482221
rect 75683 482156 75684 482220
rect 75748 482156 75749 482220
rect 75683 482155 75749 482156
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73475 436388 73541 436389
rect 73475 436324 73476 436388
rect 73540 436324 73541 436388
rect 73794 436356 74414 470898
rect 73475 436323 73541 436324
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 72739 390420 72805 390421
rect 72739 390356 72740 390420
rect 72804 390356 72805 390420
rect 72739 390355 72805 390356
rect 69611 377500 69677 377501
rect 69611 377436 69612 377500
rect 69676 377436 69677 377500
rect 69611 377435 69677 377436
rect 71635 362268 71701 362269
rect 71635 362204 71636 362268
rect 71700 362204 71701 362268
rect 71635 362203 71701 362204
rect 69059 283252 69125 283253
rect 69059 283188 69060 283252
rect 69124 283188 69125 283252
rect 69059 283187 69125 283188
rect 70163 282980 70229 282981
rect 70163 282916 70164 282980
rect 70228 282916 70229 282980
rect 70163 282915 70229 282916
rect 69427 244356 69493 244357
rect 69427 244292 69428 244356
rect 69492 244292 69493 244356
rect 69427 244291 69493 244292
rect 68875 241500 68941 241501
rect 68875 241436 68876 241500
rect 68940 241436 68941 241500
rect 68875 241435 68941 241436
rect 66667 226268 66733 226269
rect 66667 226204 66668 226268
rect 66732 226204 66733 226268
rect 66667 226203 66733 226204
rect 66115 204916 66181 204917
rect 66115 204852 66116 204916
rect 66180 204852 66181 204916
rect 66115 204851 66181 204852
rect 65931 192540 65997 192541
rect 65931 192476 65932 192540
rect 65996 192476 65997 192540
rect 65931 192475 65997 192476
rect 64643 106316 64709 106317
rect 64643 106252 64644 106316
rect 64708 106252 64709 106316
rect 64643 106251 64709 106252
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 66118 96389 66178 204851
rect 66670 98021 66730 226203
rect 66954 212614 67574 239592
rect 68875 238916 68941 238917
rect 68875 238852 68876 238916
rect 68940 238852 68941 238916
rect 68875 238851 68941 238852
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 68878 211037 68938 238851
rect 69430 238770 69490 244291
rect 69430 238710 69674 238770
rect 69614 235789 69674 238710
rect 69611 235788 69677 235789
rect 69611 235724 69612 235788
rect 69676 235724 69677 235788
rect 69611 235723 69677 235724
rect 68875 211036 68941 211037
rect 68875 210972 68876 211036
rect 68940 210972 68941 211036
rect 68875 210971 68941 210972
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 68691 143444 68757 143445
rect 68691 143380 68692 143444
rect 68756 143380 68757 143444
rect 68691 143379 68757 143380
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 136782 67574 140058
rect 66667 98020 66733 98021
rect 66667 97956 66668 98020
rect 66732 97956 66733 98020
rect 66667 97955 66733 97956
rect 66115 96388 66181 96389
rect 66115 96324 66116 96388
rect 66180 96324 66181 96388
rect 66115 96323 66181 96324
rect 66667 94212 66733 94213
rect 66667 94148 66668 94212
rect 66732 94148 66733 94212
rect 66667 94147 66733 94148
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 66670 62117 66730 94147
rect 68694 91085 68754 143379
rect 68878 92309 68938 210971
rect 70166 143309 70226 282915
rect 71638 241773 71698 362203
rect 73478 292590 73538 436323
rect 74947 433804 75013 433805
rect 74947 433740 74948 433804
rect 75012 433740 75013 433804
rect 74947 433739 75013 433740
rect 73659 433668 73725 433669
rect 73659 433604 73660 433668
rect 73724 433604 73725 433668
rect 73659 433603 73725 433604
rect 74763 433668 74829 433669
rect 74763 433604 74764 433668
rect 74828 433604 74829 433668
rect 74763 433603 74829 433604
rect 73662 389333 73722 433603
rect 73659 389332 73725 389333
rect 73659 389268 73660 389332
rect 73724 389268 73725 389332
rect 73659 389267 73725 389268
rect 73294 292530 73538 292590
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73294 283525 73354 292530
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 285592 74414 290898
rect 74766 288557 74826 433603
rect 74763 288556 74829 288557
rect 74763 288492 74764 288556
rect 74828 288492 74829 288556
rect 74763 288491 74829 288492
rect 74950 287197 75010 433739
rect 76051 433668 76117 433669
rect 76051 433604 76052 433668
rect 76116 433604 76117 433668
rect 76051 433603 76117 433604
rect 76054 307869 76114 433603
rect 77158 390421 77218 523635
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 436356 78134 438618
rect 78259 436252 78325 436253
rect 78259 436188 78260 436252
rect 78324 436188 78325 436252
rect 78259 436187 78325 436188
rect 77155 390420 77221 390421
rect 77155 390356 77156 390420
rect 77220 390356 77221 390420
rect 77155 390355 77221 390356
rect 77155 369204 77221 369205
rect 77155 369140 77156 369204
rect 77220 369140 77221 369204
rect 77155 369139 77221 369140
rect 76051 307868 76117 307869
rect 76051 307804 76052 307868
rect 76116 307804 76117 307868
rect 76051 307803 76117 307804
rect 74947 287196 75013 287197
rect 74947 287132 74948 287196
rect 75012 287132 75013 287196
rect 74947 287131 75013 287132
rect 73475 284204 73541 284205
rect 73475 284140 73476 284204
rect 73540 284140 73541 284204
rect 73475 284139 73541 284140
rect 75683 284204 75749 284205
rect 75683 284140 75684 284204
rect 75748 284140 75749 284204
rect 75683 284139 75749 284140
rect 71819 283524 71885 283525
rect 71819 283460 71820 283524
rect 71884 283460 71885 283524
rect 71819 283459 71885 283460
rect 73291 283524 73357 283525
rect 73291 283460 73292 283524
rect 73356 283460 73357 283524
rect 73291 283459 73357 283460
rect 71635 241772 71701 241773
rect 71635 241708 71636 241772
rect 71700 241708 71701 241772
rect 71635 241707 71701 241708
rect 71635 240140 71701 240141
rect 71635 240076 71636 240140
rect 71700 240076 71701 240140
rect 71635 240075 71701 240076
rect 71638 209677 71698 240075
rect 71635 209676 71701 209677
rect 71635 209612 71636 209676
rect 71700 209612 71701 209676
rect 71635 209611 71701 209612
rect 70163 143308 70229 143309
rect 70163 143244 70164 143308
rect 70228 143244 70229 143308
rect 70163 143243 70229 143244
rect 70166 143037 70226 143243
rect 70163 143036 70229 143037
rect 70163 142972 70164 143036
rect 70228 142972 70229 143036
rect 70163 142971 70229 142972
rect 69427 138684 69493 138685
rect 69427 138620 69428 138684
rect 69492 138620 69493 138684
rect 69427 138619 69493 138620
rect 69243 135148 69309 135149
rect 69243 135084 69244 135148
rect 69308 135084 69309 135148
rect 69243 135083 69309 135084
rect 69246 127125 69306 135083
rect 69430 131069 69490 138619
rect 69427 131068 69493 131069
rect 69427 131004 69428 131068
rect 69492 131004 69493 131068
rect 69427 131003 69493 131004
rect 69243 127124 69309 127125
rect 69243 127060 69244 127124
rect 69308 127060 69309 127124
rect 69243 127059 69309 127060
rect 71638 92445 71698 209611
rect 71822 139637 71882 283459
rect 72923 240004 72989 240005
rect 72923 239940 72924 240004
rect 72988 239940 72989 240004
rect 72923 239939 72989 239940
rect 71819 139636 71885 139637
rect 71819 139572 71820 139636
rect 71884 139572 71885 139636
rect 71819 139571 71885 139572
rect 72926 92445 72986 239939
rect 73294 142357 73354 283459
rect 73478 240141 73538 284139
rect 75315 283524 75381 283525
rect 75315 283460 75316 283524
rect 75380 283460 75381 283524
rect 75315 283459 75381 283460
rect 74345 255454 74665 255486
rect 74345 255218 74387 255454
rect 74623 255218 74665 255454
rect 74345 255134 74665 255218
rect 74345 254898 74387 255134
rect 74623 254898 74665 255134
rect 74345 254866 74665 254898
rect 73475 240140 73541 240141
rect 73475 240076 73476 240140
rect 73540 240076 73541 240140
rect 73475 240075 73541 240076
rect 75131 240140 75197 240141
rect 75131 240076 75132 240140
rect 75196 240076 75197 240140
rect 75131 240075 75197 240076
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73291 142356 73357 142357
rect 73291 142292 73292 142356
rect 73356 142292 73357 142356
rect 73291 142291 73357 142292
rect 73294 138277 73354 142291
rect 73291 138276 73357 138277
rect 73291 138212 73292 138276
rect 73356 138212 73357 138276
rect 73291 138211 73357 138212
rect 73794 136782 74414 146898
rect 73475 134876 73541 134877
rect 73475 134812 73476 134876
rect 73540 134812 73541 134876
rect 73475 134811 73541 134812
rect 73478 92717 73538 134811
rect 73679 111454 73999 111486
rect 73679 111218 73721 111454
rect 73957 111218 73999 111454
rect 73679 111134 73999 111218
rect 73679 110898 73721 111134
rect 73957 110898 73999 111134
rect 73679 110866 73999 110898
rect 73475 92716 73541 92717
rect 73475 92652 73476 92716
rect 73540 92652 73541 92716
rect 73475 92651 73541 92652
rect 75134 92581 75194 240075
rect 75318 139365 75378 283459
rect 75686 241773 75746 284139
rect 76971 283524 77037 283525
rect 76971 283460 76972 283524
rect 77036 283460 77037 283524
rect 76971 283459 77037 283460
rect 75683 241772 75749 241773
rect 75683 241708 75684 241772
rect 75748 241708 75749 241772
rect 75683 241707 75749 241708
rect 76974 176629 77034 283459
rect 77158 241773 77218 369139
rect 77514 367174 78134 388356
rect 78262 387021 78322 436187
rect 79731 436116 79797 436117
rect 79731 436052 79732 436116
rect 79796 436052 79797 436116
rect 79731 436051 79797 436052
rect 78443 433668 78509 433669
rect 78443 433604 78444 433668
rect 78508 433604 78509 433668
rect 78443 433603 78509 433604
rect 78446 388517 78506 433603
rect 78443 388516 78509 388517
rect 78443 388452 78444 388516
rect 78508 388452 78509 388516
rect 78443 388451 78509 388452
rect 78259 387020 78325 387021
rect 78259 386956 78260 387020
rect 78324 386956 78325 387020
rect 78259 386955 78325 386956
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 79734 317525 79794 436051
rect 79918 390149 79978 581163
rect 81019 580820 81085 580821
rect 81019 580756 81020 580820
rect 81084 580756 81085 580820
rect 81019 580755 81085 580756
rect 83963 580820 84029 580821
rect 83963 580756 83964 580820
rect 84028 580756 84029 580820
rect 83963 580755 84029 580756
rect 89299 580820 89365 580821
rect 89299 580756 89300 580820
rect 89364 580756 89365 580820
rect 89299 580755 89365 580756
rect 81022 526829 81082 580755
rect 81609 543454 81929 543486
rect 81609 543218 81651 543454
rect 81887 543218 81929 543454
rect 81609 543134 81929 543218
rect 81609 542898 81651 543134
rect 81887 542898 81929 543134
rect 81609 542866 81929 542898
rect 82859 538796 82925 538797
rect 82859 538732 82860 538796
rect 82924 538732 82925 538796
rect 82859 538731 82925 538732
rect 81019 526828 81085 526829
rect 81019 526764 81020 526828
rect 81084 526764 81085 526828
rect 81019 526763 81085 526764
rect 81022 525877 81082 526763
rect 81019 525876 81085 525877
rect 81019 525812 81020 525876
rect 81084 525812 81085 525876
rect 81019 525811 81085 525812
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 82675 463588 82741 463589
rect 82675 463524 82676 463588
rect 82740 463524 82741 463588
rect 82675 463523 82741 463524
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 436356 81854 442338
rect 80099 434348 80165 434349
rect 80099 434284 80100 434348
rect 80164 434284 80165 434348
rect 80099 434283 80165 434284
rect 79915 390148 79981 390149
rect 79915 390084 79916 390148
rect 79980 390084 79981 390148
rect 79915 390083 79981 390084
rect 80102 382941 80162 434283
rect 82678 391917 82738 463523
rect 82307 391916 82373 391917
rect 82307 391852 82308 391916
rect 82372 391852 82373 391916
rect 82307 391851 82373 391852
rect 82675 391916 82741 391917
rect 82675 391852 82676 391916
rect 82740 391852 82741 391916
rect 82675 391851 82741 391852
rect 82310 390965 82370 391851
rect 82307 390964 82373 390965
rect 82307 390900 82308 390964
rect 82372 390900 82373 390964
rect 82307 390899 82373 390900
rect 82862 390693 82922 538731
rect 83966 463589 84026 580755
rect 85575 561454 85895 561486
rect 85575 561218 85617 561454
rect 85853 561218 85895 561454
rect 85575 561134 85895 561218
rect 85575 560898 85617 561134
rect 85853 560898 85895 561134
rect 85575 560866 85895 560898
rect 84954 518614 85574 537166
rect 88931 530636 88997 530637
rect 88931 530572 88932 530636
rect 88996 530572 88997 530636
rect 88931 530571 88997 530572
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 83963 463588 84029 463589
rect 83963 463524 83964 463588
rect 84028 463524 84029 463588
rect 83963 463523 84029 463524
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 436356 85574 446058
rect 84699 436116 84765 436117
rect 84699 436052 84700 436116
rect 84764 436052 84765 436116
rect 84699 436051 84765 436052
rect 83043 434484 83109 434485
rect 83043 434420 83044 434484
rect 83108 434420 83109 434484
rect 83043 434419 83109 434420
rect 82859 390692 82925 390693
rect 82859 390628 82860 390692
rect 82924 390628 82925 390692
rect 82859 390627 82925 390628
rect 80099 382940 80165 382941
rect 80099 382876 80100 382940
rect 80164 382876 80165 382940
rect 80099 382875 80165 382876
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 79731 317524 79797 317525
rect 79731 317460 79732 317524
rect 79796 317460 79797 317524
rect 79731 317459 79797 317460
rect 79734 316050 79794 317459
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285592 78134 294618
rect 79182 315990 79794 316050
rect 78443 291140 78509 291141
rect 78443 291076 78444 291140
rect 78508 291076 78509 291140
rect 78443 291075 78509 291076
rect 78259 284204 78325 284205
rect 78259 284140 78260 284204
rect 78324 284140 78325 284204
rect 78259 284139 78325 284140
rect 78262 248430 78322 284139
rect 78078 248370 78322 248430
rect 78078 241773 78138 248370
rect 78446 241773 78506 291075
rect 79182 288693 79242 315990
rect 81234 298894 81854 334338
rect 83046 309093 83106 434419
rect 84515 434348 84581 434349
rect 84515 434284 84516 434348
rect 84580 434284 84581 434348
rect 84515 434283 84581 434284
rect 84518 390965 84578 434283
rect 84515 390964 84581 390965
rect 84515 390900 84516 390964
rect 84580 390900 84581 390964
rect 84515 390899 84581 390900
rect 84702 387565 84762 436051
rect 85803 434348 85869 434349
rect 85803 434284 85804 434348
rect 85868 434284 85869 434348
rect 85803 434283 85869 434284
rect 84699 387564 84765 387565
rect 84699 387500 84700 387564
rect 84764 387500 84765 387564
rect 84699 387499 84765 387500
rect 84954 374614 85574 388356
rect 85806 385117 85866 434283
rect 86723 433668 86789 433669
rect 86723 433604 86724 433668
rect 86788 433604 86789 433668
rect 86723 433603 86789 433604
rect 87091 433668 87157 433669
rect 87091 433604 87092 433668
rect 87156 433604 87157 433668
rect 87091 433603 87157 433604
rect 87459 433668 87525 433669
rect 87459 433604 87460 433668
rect 87524 433604 87525 433668
rect 87459 433603 87525 433604
rect 85803 385116 85869 385117
rect 85803 385052 85804 385116
rect 85868 385052 85869 385116
rect 85803 385051 85869 385052
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 83043 309092 83109 309093
rect 83043 309028 83044 309092
rect 83108 309028 83109 309092
rect 83043 309027 83109 309028
rect 84515 307732 84581 307733
rect 84515 307668 84516 307732
rect 84580 307668 84581 307732
rect 84515 307667 84581 307668
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 80651 291140 80717 291141
rect 80651 291076 80652 291140
rect 80716 291076 80717 291140
rect 80651 291075 80717 291076
rect 79179 288692 79245 288693
rect 79179 288628 79180 288692
rect 79244 288628 79245 288692
rect 79179 288627 79245 288628
rect 79915 283116 79981 283117
rect 79915 283052 79916 283116
rect 79980 283052 79981 283116
rect 79915 283051 79981 283052
rect 78977 273454 79297 273486
rect 78977 273218 79019 273454
rect 79255 273218 79297 273454
rect 78977 273134 79297 273218
rect 78977 272898 79019 273134
rect 79255 272898 79297 273134
rect 78977 272866 79297 272898
rect 77155 241772 77221 241773
rect 77155 241708 77156 241772
rect 77220 241708 77221 241772
rect 77155 241707 77221 241708
rect 78075 241772 78141 241773
rect 78075 241708 78076 241772
rect 78140 241708 78141 241772
rect 78075 241707 78141 241708
rect 78443 241772 78509 241773
rect 78443 241708 78444 241772
rect 78508 241708 78509 241772
rect 78443 241707 78509 241708
rect 77155 238644 77221 238645
rect 77155 238580 77156 238644
rect 77220 238580 77221 238644
rect 77155 238579 77221 238580
rect 76971 176628 77037 176629
rect 76971 176564 76972 176628
rect 77036 176564 77037 176628
rect 76971 176563 77037 176564
rect 76974 176221 77034 176563
rect 76971 176220 77037 176221
rect 76971 176156 76972 176220
rect 77036 176156 77037 176220
rect 76971 176155 77037 176156
rect 76971 140860 77037 140861
rect 76971 140796 76972 140860
rect 77036 140796 77037 140860
rect 76971 140795 77037 140796
rect 75315 139364 75381 139365
rect 75315 139300 75316 139364
rect 75380 139300 75381 139364
rect 75315 139299 75381 139300
rect 75315 134740 75381 134741
rect 75315 134676 75316 134740
rect 75380 134676 75381 134740
rect 75315 134675 75381 134676
rect 75318 92717 75378 134675
rect 75315 92716 75381 92717
rect 75315 92652 75316 92716
rect 75380 92652 75381 92716
rect 75315 92651 75381 92652
rect 75131 92580 75197 92581
rect 75131 92516 75132 92580
rect 75196 92516 75197 92580
rect 75131 92515 75197 92516
rect 76974 92445 77034 140795
rect 77158 92717 77218 238579
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 136782 78134 150618
rect 79918 137325 79978 283051
rect 80654 241773 80714 291075
rect 81234 285592 81854 298338
rect 81939 294676 82005 294677
rect 81939 294612 81940 294676
rect 82004 294612 82005 294676
rect 81939 294611 82005 294612
rect 81942 241773 82002 294611
rect 83411 285700 83477 285701
rect 83411 285636 83412 285700
rect 83476 285636 83477 285700
rect 83411 285635 83477 285636
rect 83414 282981 83474 285635
rect 82675 282980 82741 282981
rect 82675 282916 82676 282980
rect 82740 282916 82741 282980
rect 82675 282915 82741 282916
rect 83411 282980 83477 282981
rect 83411 282916 83412 282980
rect 83476 282916 83477 282980
rect 83411 282915 83477 282916
rect 80651 241772 80717 241773
rect 80651 241708 80652 241772
rect 80716 241708 80717 241772
rect 80651 241707 80717 241708
rect 81939 241772 82005 241773
rect 81939 241708 81940 241772
rect 82004 241708 82005 241772
rect 81939 241707 82005 241708
rect 81234 226894 81854 239592
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 82678 176765 82738 282915
rect 83414 177309 83474 282915
rect 83609 255454 83929 255486
rect 83609 255218 83651 255454
rect 83887 255218 83929 255454
rect 83609 255134 83929 255218
rect 83609 254898 83651 255134
rect 83887 254898 83929 255134
rect 83609 254866 83929 254898
rect 84518 241773 84578 307667
rect 84954 302614 85574 338058
rect 86726 316029 86786 433603
rect 86723 316028 86789 316029
rect 86723 315964 86724 316028
rect 86788 315964 86789 316028
rect 86723 315963 86789 315964
rect 86726 306509 86786 315963
rect 86723 306508 86789 306509
rect 86723 306444 86724 306508
rect 86788 306444 86789 306508
rect 86723 306443 86789 306444
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 285592 85574 302058
rect 86539 301612 86605 301613
rect 86539 301548 86540 301612
rect 86604 301548 86605 301612
rect 86539 301547 86605 301548
rect 84699 283116 84765 283117
rect 84699 283052 84700 283116
rect 84764 283052 84765 283116
rect 84699 283051 84765 283052
rect 84515 241772 84581 241773
rect 84515 241708 84516 241772
rect 84580 241708 84581 241772
rect 84515 241707 84581 241708
rect 83411 177308 83477 177309
rect 83411 177244 83412 177308
rect 83476 177244 83477 177308
rect 83411 177243 83477 177244
rect 82675 176764 82741 176765
rect 82675 176700 82676 176764
rect 82740 176700 82741 176764
rect 82675 176699 82741 176700
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 79915 137324 79981 137325
rect 79915 137260 79916 137324
rect 79980 137260 79981 137324
rect 79915 137259 79981 137260
rect 81234 136782 81854 154338
rect 84702 142085 84762 283051
rect 86542 241773 86602 301547
rect 87094 293181 87154 433603
rect 87462 386885 87522 433603
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 88934 390693 88994 530571
rect 89302 484397 89362 580755
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 96659 553484 96725 553485
rect 96659 553420 96660 553484
rect 96724 553420 96725 553484
rect 96659 553419 96725 553420
rect 96662 551309 96722 553419
rect 96659 551308 96725 551309
rect 96659 551244 96660 551308
rect 96724 551244 96725 551308
rect 96659 551243 96725 551244
rect 96843 547092 96909 547093
rect 96843 547028 96844 547092
rect 96908 547028 96909 547092
rect 96843 547027 96909 547028
rect 89540 543454 89860 543486
rect 89540 543218 89582 543454
rect 89818 543218 89860 543454
rect 89540 543134 89860 543218
rect 89540 542898 89582 543134
rect 89818 542898 89860 543134
rect 89540 542866 89860 542898
rect 91794 525454 92414 537166
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 89299 484396 89365 484397
rect 89299 484332 89300 484396
rect 89364 484332 89365 484396
rect 89299 484331 89365 484332
rect 91323 469844 91389 469845
rect 91323 469780 91324 469844
rect 91388 469780 91389 469844
rect 91323 469779 91389 469780
rect 89667 433668 89733 433669
rect 89667 433604 89668 433668
rect 89732 433604 89733 433668
rect 89667 433603 89733 433604
rect 90035 433668 90101 433669
rect 90035 433604 90036 433668
rect 90100 433604 90101 433668
rect 90035 433603 90101 433604
rect 89670 398850 89730 433603
rect 89670 398790 89914 398850
rect 88931 390692 88997 390693
rect 88931 390628 88932 390692
rect 88996 390628 88997 390692
rect 88931 390627 88997 390628
rect 89854 389190 89914 398790
rect 89670 389130 89914 389190
rect 87459 386884 87525 386885
rect 87459 386820 87460 386884
rect 87524 386820 87525 386884
rect 87459 386819 87525 386820
rect 89670 304197 89730 389130
rect 90038 311133 90098 433603
rect 91326 390829 91386 469779
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 436356 92414 452898
rect 95514 529174 96134 537166
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 96846 519485 96906 547027
rect 99234 532894 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 100707 549404 100773 549405
rect 100707 549340 100708 549404
rect 100772 549340 100773 549404
rect 100707 549339 100773 549340
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 97027 527780 97093 527781
rect 97027 527716 97028 527780
rect 97092 527716 97093 527780
rect 97027 527715 97093 527716
rect 96843 519484 96909 519485
rect 96843 519420 96844 519484
rect 96908 519420 96909 519484
rect 96843 519419 96909 519420
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 96843 457468 96909 457469
rect 96843 457404 96844 457468
rect 96908 457404 96909 457468
rect 96843 457403 96909 457404
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 436356 96134 456618
rect 94451 436116 94517 436117
rect 94451 436052 94452 436116
rect 94516 436052 94517 436116
rect 94451 436051 94517 436052
rect 92611 434212 92677 434213
rect 92611 434148 92612 434212
rect 92676 434148 92677 434212
rect 92611 434147 92677 434148
rect 91507 433668 91573 433669
rect 91507 433604 91508 433668
rect 91572 433604 91573 433668
rect 91507 433603 91573 433604
rect 91323 390828 91389 390829
rect 91323 390764 91324 390828
rect 91388 390764 91389 390828
rect 91323 390763 91389 390764
rect 90035 311132 90101 311133
rect 90035 311068 90036 311132
rect 90100 311068 90101 311132
rect 90035 311067 90101 311068
rect 91510 305829 91570 433603
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91507 305828 91573 305829
rect 91507 305764 91508 305828
rect 91572 305764 91573 305828
rect 91507 305763 91573 305764
rect 89667 304196 89733 304197
rect 89667 304132 89668 304196
rect 89732 304132 89733 304196
rect 89667 304131 89733 304132
rect 87091 293180 87157 293181
rect 87091 293116 87092 293180
rect 87156 293116 87157 293180
rect 87091 293115 87157 293116
rect 91507 290052 91573 290053
rect 91507 289988 91508 290052
rect 91572 289988 91573 290052
rect 91507 289987 91573 289988
rect 88011 289644 88077 289645
rect 88011 289580 88012 289644
rect 88076 289580 88077 289644
rect 88011 289579 88077 289580
rect 86723 285700 86789 285701
rect 86723 285636 86724 285700
rect 86788 285636 86789 285700
rect 86723 285635 86789 285636
rect 86726 282981 86786 285635
rect 86723 282980 86789 282981
rect 86723 282916 86724 282980
rect 86788 282916 86789 282980
rect 86723 282915 86789 282916
rect 86539 241772 86605 241773
rect 86539 241708 86540 241772
rect 86604 241708 86605 241772
rect 86539 241707 86605 241708
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 86726 172413 86786 282915
rect 88014 241637 88074 289579
rect 91139 284204 91205 284205
rect 91139 284140 91140 284204
rect 91204 284140 91205 284204
rect 91139 284139 91205 284140
rect 89851 283524 89917 283525
rect 89851 283460 89852 283524
rect 89916 283460 89917 283524
rect 89851 283459 89917 283460
rect 88747 282980 88813 282981
rect 88747 282916 88748 282980
rect 88812 282916 88813 282980
rect 88747 282915 88813 282916
rect 88241 273454 88561 273486
rect 88241 273218 88283 273454
rect 88519 273218 88561 273454
rect 88241 273134 88561 273218
rect 88241 272898 88283 273134
rect 88519 272898 88561 273134
rect 88241 272866 88561 272898
rect 88011 241636 88077 241637
rect 88011 241572 88012 241636
rect 88076 241572 88077 241636
rect 88011 241571 88077 241572
rect 88014 240141 88074 241571
rect 88011 240140 88077 240141
rect 88011 240076 88012 240140
rect 88076 240076 88077 240140
rect 88011 240075 88077 240076
rect 86723 172412 86789 172413
rect 86723 172348 86724 172412
rect 86788 172348 86789 172412
rect 86723 172347 86789 172348
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84699 142084 84765 142085
rect 84699 142020 84700 142084
rect 84764 142020 84765 142084
rect 84699 142019 84765 142020
rect 84954 136782 85574 158058
rect 88750 143581 88810 282915
rect 89854 144805 89914 283459
rect 91142 241773 91202 284139
rect 91139 241772 91205 241773
rect 91139 241708 91140 241772
rect 91204 241708 91205 241772
rect 91139 241707 91205 241708
rect 91142 240141 91202 241707
rect 91510 241637 91570 289987
rect 91794 285592 92414 308898
rect 92614 308413 92674 434147
rect 92795 433668 92861 433669
rect 92795 433604 92796 433668
rect 92860 433604 92861 433668
rect 92795 433603 92861 433604
rect 92798 312493 92858 433603
rect 94454 382941 94514 436051
rect 95187 434348 95253 434349
rect 95187 434284 95188 434348
rect 95252 434284 95253 434348
rect 95187 434283 95253 434284
rect 94451 382940 94517 382941
rect 94451 382876 94452 382940
rect 94516 382876 94517 382940
rect 94451 382875 94517 382876
rect 95190 313989 95250 434283
rect 96846 390829 96906 457403
rect 97030 390829 97090 527715
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 436356 99854 460338
rect 100155 434348 100221 434349
rect 100155 434284 100156 434348
rect 100220 434284 100221 434348
rect 100155 434283 100221 434284
rect 98499 433804 98565 433805
rect 98499 433740 98500 433804
rect 98564 433740 98565 433804
rect 98499 433739 98565 433740
rect 97947 433668 98013 433669
rect 97947 433604 97948 433668
rect 98012 433604 98013 433668
rect 97947 433603 98013 433604
rect 96843 390828 96909 390829
rect 96843 390764 96844 390828
rect 96908 390764 96909 390828
rect 96843 390763 96909 390764
rect 97027 390828 97093 390829
rect 97027 390764 97028 390828
rect 97092 390764 97093 390828
rect 97027 390763 97093 390764
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95187 313988 95253 313989
rect 95187 313924 95188 313988
rect 95252 313924 95253 313988
rect 95187 313923 95253 313924
rect 95514 313174 96134 348618
rect 97763 320244 97829 320245
rect 97763 320180 97764 320244
rect 97828 320180 97829 320244
rect 97763 320179 97829 320180
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 92795 312492 92861 312493
rect 92795 312428 92796 312492
rect 92860 312428 92861 312492
rect 92795 312427 92861 312428
rect 92611 308412 92677 308413
rect 92611 308348 92612 308412
rect 92676 308348 92677 308412
rect 92611 308347 92677 308348
rect 95514 285592 96134 312618
rect 93347 283524 93413 283525
rect 93347 283460 93348 283524
rect 93412 283460 93413 283524
rect 93347 283459 93413 283460
rect 92873 255454 93193 255486
rect 92873 255218 92915 255454
rect 93151 255218 93193 255454
rect 92873 255134 93193 255218
rect 92873 254898 92915 255134
rect 93151 254898 93193 255134
rect 92873 254866 93193 254898
rect 91507 241636 91573 241637
rect 91507 241572 91508 241636
rect 91572 241572 91573 241636
rect 91507 241571 91573 241572
rect 91139 240140 91205 240141
rect 91139 240076 91140 240140
rect 91204 240076 91205 240140
rect 91139 240075 91205 240076
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 89851 144804 89917 144805
rect 89851 144740 89852 144804
rect 89916 144740 89917 144804
rect 89851 144739 89917 144740
rect 88747 143580 88813 143581
rect 88747 143516 88748 143580
rect 88812 143516 88813 143580
rect 88747 143515 88813 143516
rect 91794 136782 92414 164898
rect 92611 144804 92677 144805
rect 92611 144740 92612 144804
rect 92676 144740 92677 144804
rect 92611 144739 92677 144740
rect 77644 129454 77964 129486
rect 77644 129218 77686 129454
rect 77922 129218 77964 129454
rect 77644 129134 77964 129218
rect 77644 128898 77686 129134
rect 77922 128898 77964 129134
rect 77644 128866 77964 128898
rect 85575 129454 85895 129486
rect 85575 129218 85617 129454
rect 85853 129218 85895 129454
rect 85575 129134 85895 129218
rect 85575 128898 85617 129134
rect 85853 128898 85895 129134
rect 85575 128866 85895 128898
rect 81609 111454 81929 111486
rect 81609 111218 81651 111454
rect 81887 111218 81929 111454
rect 81609 111134 81929 111218
rect 81609 110898 81651 111134
rect 81887 110898 81929 111134
rect 81609 110866 81929 110898
rect 89540 111454 89860 111486
rect 89540 111218 89582 111454
rect 89818 111218 89860 111454
rect 89540 111134 89860 111218
rect 89540 110898 89582 111134
rect 89818 110898 89860 111134
rect 89540 110866 89860 110898
rect 92614 92717 92674 144739
rect 93350 140861 93410 283459
rect 97766 283389 97826 320179
rect 97950 307053 98010 433603
rect 98502 311133 98562 433739
rect 99971 433668 100037 433669
rect 99971 433604 99972 433668
rect 100036 433604 100037 433668
rect 99971 433603 100037 433604
rect 99234 352894 99854 388356
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 98499 311132 98565 311133
rect 98499 311068 98500 311132
rect 98564 311068 98565 311132
rect 98499 311067 98565 311068
rect 97947 307052 98013 307053
rect 97947 306988 97948 307052
rect 98012 306988 98013 307052
rect 97947 306987 98013 306988
rect 99234 285592 99854 316338
rect 99974 287877 100034 433603
rect 100158 387973 100218 434283
rect 100710 390421 100770 549339
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 104939 551988 105005 551989
rect 104939 551924 104940 551988
rect 105004 551924 105005 551988
rect 104939 551923 105005 551924
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 104203 534716 104269 534717
rect 104203 534652 104204 534716
rect 104268 534652 104269 534716
rect 104203 534651 104269 534652
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 436356 103574 464058
rect 102731 436252 102797 436253
rect 102731 436188 102732 436252
rect 102796 436188 102797 436252
rect 102731 436187 102797 436188
rect 100891 433668 100957 433669
rect 100891 433604 100892 433668
rect 100956 433604 100957 433668
rect 100891 433603 100957 433604
rect 100707 390420 100773 390421
rect 100707 390356 100708 390420
rect 100772 390356 100773 390420
rect 100707 390355 100773 390356
rect 100155 387972 100221 387973
rect 100155 387908 100156 387972
rect 100220 387908 100221 387972
rect 100155 387907 100221 387908
rect 100894 385933 100954 433603
rect 100891 385932 100957 385933
rect 100891 385868 100892 385932
rect 100956 385868 100957 385932
rect 100891 385867 100957 385868
rect 102734 382397 102794 436187
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 104206 390421 104266 534651
rect 104942 390421 105002 551923
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 106779 530772 106845 530773
rect 106779 530708 106780 530772
rect 106844 530708 106845 530772
rect 106779 530707 106845 530708
rect 106782 456109 106842 530707
rect 109794 507454 110414 542898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 111747 533356 111813 533357
rect 111747 533292 111748 533356
rect 111812 533292 111813 533356
rect 111747 533291 111813 533292
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 106779 456108 106845 456109
rect 106779 456044 106780 456108
rect 106844 456044 106845 456108
rect 106779 456043 106845 456044
rect 106782 451290 106842 456043
rect 106782 451230 107578 451290
rect 105123 433668 105189 433669
rect 105123 433604 105124 433668
rect 105188 433604 105189 433668
rect 105123 433603 105189 433604
rect 106411 433668 106477 433669
rect 106411 433604 106412 433668
rect 106476 433604 106477 433668
rect 106411 433603 106477 433604
rect 104203 390420 104269 390421
rect 104203 390356 104204 390420
rect 104268 390356 104269 390420
rect 104203 390355 104269 390356
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 102731 382396 102797 382397
rect 102731 382332 102732 382396
rect 102796 382332 102797 382396
rect 102731 382331 102797 382332
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 101259 304196 101325 304197
rect 101259 304132 101260 304196
rect 101324 304132 101325 304196
rect 101259 304131 101325 304132
rect 99971 287876 100037 287877
rect 99971 287812 99972 287876
rect 100036 287812 100037 287876
rect 99971 287811 100037 287812
rect 94083 283388 94149 283389
rect 94083 283324 94084 283388
rect 94148 283324 94149 283388
rect 94083 283323 94149 283324
rect 97763 283388 97829 283389
rect 97763 283324 97764 283388
rect 97828 283324 97829 283388
rect 97763 283323 97829 283324
rect 94086 277410 94146 283323
rect 99971 280260 100037 280261
rect 99971 280196 99972 280260
rect 100036 280196 100037 280260
rect 99971 280195 100037 280196
rect 93902 277350 94146 277410
rect 93902 236469 93962 277350
rect 98131 251292 98197 251293
rect 98131 251228 98132 251292
rect 98196 251228 98197 251292
rect 98131 251227 98197 251228
rect 93899 236468 93965 236469
rect 93899 236404 93900 236468
rect 93964 236404 93965 236468
rect 93899 236403 93965 236404
rect 93899 230484 93965 230485
rect 93899 230420 93900 230484
rect 93964 230420 93965 230484
rect 93899 230419 93965 230420
rect 93347 140860 93413 140861
rect 93347 140796 93348 140860
rect 93412 140796 93413 140860
rect 93347 140795 93413 140796
rect 93715 134740 93781 134741
rect 93715 134676 93716 134740
rect 93780 134676 93781 134740
rect 93715 134675 93781 134676
rect 93718 125610 93778 134675
rect 93902 129570 93962 230419
rect 94083 211852 94149 211853
rect 94083 211788 94084 211852
rect 94148 211788 94149 211852
rect 94083 211787 94149 211788
rect 94086 134741 94146 211787
rect 95514 205174 96134 239592
rect 98134 238770 98194 251227
rect 97950 238710 98194 238770
rect 97950 223549 98010 238710
rect 97947 223548 98013 223549
rect 97947 223484 97948 223548
rect 98012 223484 98013 223548
rect 97947 223483 98013 223484
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 136782 96134 168618
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 96291 149292 96357 149293
rect 96291 149228 96292 149292
rect 96356 149228 96357 149292
rect 96291 149227 96357 149228
rect 94083 134740 94149 134741
rect 94083 134676 94084 134740
rect 94148 134676 94149 134740
rect 94083 134675 94149 134676
rect 94635 129572 94701 129573
rect 94635 129570 94636 129572
rect 93902 129510 94636 129570
rect 94635 129508 94636 129510
rect 94700 129508 94701 129572
rect 94635 129507 94701 129508
rect 93718 125550 94146 125610
rect 77155 92716 77221 92717
rect 77155 92652 77156 92716
rect 77220 92652 77221 92716
rect 77155 92651 77221 92652
rect 92611 92716 92677 92717
rect 92611 92652 92612 92716
rect 92676 92652 92677 92716
rect 92611 92651 92677 92652
rect 71635 92444 71701 92445
rect 71635 92380 71636 92444
rect 71700 92380 71701 92444
rect 71635 92379 71701 92380
rect 72923 92444 72989 92445
rect 72923 92380 72924 92444
rect 72988 92380 72989 92444
rect 72923 92379 72989 92380
rect 76971 92444 77037 92445
rect 76971 92380 76972 92444
rect 77036 92380 77037 92444
rect 76971 92379 77037 92380
rect 68875 92308 68941 92309
rect 68875 92244 68876 92308
rect 68940 92244 68941 92308
rect 68875 92243 68941 92244
rect 68691 91084 68757 91085
rect 68691 91020 68692 91084
rect 68756 91020 68757 91084
rect 68691 91019 68757 91020
rect 66954 68614 67574 90782
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66667 62116 66733 62117
rect 66667 62052 66668 62116
rect 66732 62052 66733 62116
rect 66667 62051 66733 62052
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 90782
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 90782
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 90782
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 90782
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 90782
rect 94086 90405 94146 125550
rect 96294 108901 96354 149227
rect 99234 136894 99854 172338
rect 99974 144805 100034 280195
rect 101262 278629 101322 304131
rect 102954 284614 103574 320058
rect 105126 315349 105186 433603
rect 105123 315348 105189 315349
rect 105123 315284 105124 315348
rect 105188 315284 105189 315348
rect 105123 315283 105189 315284
rect 106414 309773 106474 433603
rect 107518 390965 107578 451230
rect 109794 436356 110414 470898
rect 109539 433668 109605 433669
rect 109539 433604 109540 433668
rect 109604 433604 109605 433668
rect 109539 433603 109605 433604
rect 111011 433668 111077 433669
rect 111011 433604 111012 433668
rect 111076 433604 111077 433668
rect 111011 433603 111077 433604
rect 107515 390964 107581 390965
rect 107515 390900 107516 390964
rect 107580 390900 107581 390964
rect 107515 390899 107581 390900
rect 109542 318069 109602 433603
rect 109794 363454 110414 388356
rect 111014 370565 111074 433603
rect 111750 422310 111810 533291
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113219 458828 113285 458829
rect 113219 458764 113220 458828
rect 113284 458764 113285 458828
rect 113219 458763 113285 458764
rect 113035 454068 113101 454069
rect 113035 454004 113036 454068
rect 113100 454004 113101 454068
rect 113035 454003 113101 454004
rect 111750 422250 112178 422310
rect 112118 402661 112178 422250
rect 112115 402660 112181 402661
rect 112115 402596 112116 402660
rect 112180 402596 112181 402660
rect 112115 402595 112181 402596
rect 113038 398989 113098 454003
rect 112115 398988 112181 398989
rect 112115 398924 112116 398988
rect 112180 398924 112181 398988
rect 112115 398923 112181 398924
rect 113035 398988 113101 398989
rect 113035 398924 113036 398988
rect 113100 398924 113101 398988
rect 113035 398923 113101 398924
rect 112118 393330 112178 398923
rect 113222 396405 113282 458763
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 436356 114134 438618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 114507 430132 114573 430133
rect 114507 430068 114508 430132
rect 114572 430068 114573 430132
rect 114507 430067 114573 430068
rect 113219 396404 113285 396405
rect 113219 396340 113220 396404
rect 113284 396340 113285 396404
rect 113219 396339 113285 396340
rect 111750 393270 112178 393330
rect 111750 390557 111810 393270
rect 111747 390556 111813 390557
rect 111747 390492 111748 390556
rect 111812 390492 111813 390556
rect 111747 390491 111813 390492
rect 111011 370564 111077 370565
rect 111011 370500 111012 370564
rect 111076 370500 111077 370564
rect 111011 370499 111077 370500
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109539 318068 109605 318069
rect 109539 318004 109540 318068
rect 109604 318004 109605 318068
rect 109539 318003 109605 318004
rect 109542 312493 109602 318003
rect 109539 312492 109605 312493
rect 109539 312428 109540 312492
rect 109604 312428 109605 312492
rect 109539 312427 109605 312428
rect 106411 309772 106477 309773
rect 106411 309708 106412 309772
rect 106476 309708 106477 309772
rect 106411 309707 106477 309708
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 101259 278628 101325 278629
rect 101259 278564 101260 278628
rect 101324 278564 101325 278628
rect 101259 278563 101325 278564
rect 100707 255780 100773 255781
rect 100707 255716 100708 255780
rect 100772 255716 100773 255780
rect 100707 255715 100773 255716
rect 100710 149293 100770 255715
rect 101259 252516 101325 252517
rect 101259 252452 101260 252516
rect 101324 252452 101325 252516
rect 101259 252451 101325 252452
rect 101262 216749 101322 252451
rect 102954 248614 103574 284058
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 103835 275228 103901 275229
rect 103835 275164 103836 275228
rect 103900 275164 103901 275228
rect 103835 275163 103901 275164
rect 103838 258090 103898 275163
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 101259 216748 101325 216749
rect 101259 216684 101260 216748
rect 101324 216684 101325 216748
rect 101259 216683 101325 216684
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 100707 149292 100773 149293
rect 100707 149228 100708 149292
rect 100772 149228 100773 149292
rect 100707 149227 100773 149228
rect 99971 144804 100037 144805
rect 99971 144740 99972 144804
rect 100036 144740 100037 144804
rect 99971 144739 100037 144740
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 97211 109580 97277 109581
rect 97211 109516 97212 109580
rect 97276 109516 97277 109580
rect 97211 109515 97277 109516
rect 96291 108900 96357 108901
rect 96291 108836 96292 108900
rect 96356 108836 96357 108900
rect 96291 108835 96357 108836
rect 94819 93940 94885 93941
rect 94819 93876 94820 93940
rect 94884 93876 94885 93940
rect 94819 93875 94885 93876
rect 94822 92037 94882 93875
rect 97214 92853 97274 109515
rect 99234 100894 99854 136338
rect 102954 140614 103574 176058
rect 103654 258030 103898 258090
rect 103654 151830 103714 258030
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 106043 236604 106109 236605
rect 106043 236540 106044 236604
rect 106108 236540 106109 236604
rect 106043 236539 106109 236540
rect 103654 151770 103898 151830
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 101995 113796 102061 113797
rect 101995 113732 101996 113796
rect 102060 113732 102061 113796
rect 101995 113731 102061 113732
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 97211 92852 97277 92853
rect 97211 92788 97212 92852
rect 97276 92788 97277 92852
rect 97211 92787 97277 92788
rect 94819 92036 94885 92037
rect 94819 91972 94820 92036
rect 94884 91972 94885 92036
rect 94819 91971 94885 91972
rect 94083 90404 94149 90405
rect 94083 90340 94084 90404
rect 94148 90340 94149 90404
rect 94083 90339 94149 90340
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 90782
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 101998 3501 102058 113731
rect 102954 104614 103574 140058
rect 103838 128485 103898 151770
rect 103835 128484 103901 128485
rect 103835 128420 103836 128484
rect 103900 128420 103901 128484
rect 103835 128419 103901 128420
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 106046 90541 106106 236539
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 106043 90540 106109 90541
rect 106043 90476 106044 90540
rect 106108 90476 106109 90540
rect 106043 90475 106109 90476
rect 106046 89861 106106 90475
rect 106043 89860 106109 89861
rect 106043 89796 106044 89860
rect 106108 89796 106109 89860
rect 106043 89795 106109 89796
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 101995 3500 102061 3501
rect 101995 3436 101996 3500
rect 102060 3436 102061 3500
rect 101995 3435 102061 3436
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 367174 114134 388356
rect 114510 382941 114570 430067
rect 114691 413812 114757 413813
rect 114691 413748 114692 413812
rect 114756 413748 114757 413812
rect 114691 413747 114757 413748
rect 114694 391509 114754 413747
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 114691 391508 114757 391509
rect 114691 391444 114692 391508
rect 114756 391444 114757 391508
rect 114691 391443 114757 391444
rect 114507 382940 114573 382941
rect 114507 382876 114508 382940
rect 114572 382876 114573 382940
rect 114507 382875 114573 382876
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 155723 603260 155789 603261
rect 155723 603196 155724 603260
rect 155788 603196 155789 603260
rect 155723 603195 155789 603196
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 151675 547092 151741 547093
rect 151675 547028 151676 547092
rect 151740 547028 151741 547092
rect 151675 547027 151741 547028
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 148915 458148 148981 458149
rect 148915 458084 148916 458148
rect 148980 458084 148981 458148
rect 148915 458083 148981 458084
rect 147443 454068 147509 454069
rect 147443 454004 147444 454068
rect 147508 454004 147509 454068
rect 147443 454003 147509 454004
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 141371 336156 141437 336157
rect 141371 336092 141372 336156
rect 141436 336092 141437 336156
rect 141371 336091 141437 336092
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 141374 30973 141434 336091
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 141371 30972 141437 30973
rect 141371 30908 141372 30972
rect 141436 30908 141437 30972
rect 141371 30907 141437 30908
rect 145794 3454 146414 38898
rect 147446 3501 147506 454003
rect 148918 295221 148978 458083
rect 149514 439174 150134 474618
rect 150939 456924 151005 456925
rect 150939 456860 150940 456924
rect 151004 456860 151005 456924
rect 150939 456859 151005 456860
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 150942 418301 151002 456859
rect 150939 418300 151005 418301
rect 150939 418236 150940 418300
rect 151004 418236 151005 418300
rect 150939 418235 151005 418236
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 148915 295220 148981 295221
rect 148915 295156 148916 295220
rect 148980 295156 148981 295220
rect 148915 295155 148981 295156
rect 149514 295174 150134 330618
rect 151678 302837 151738 547027
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 151675 302836 151741 302837
rect 151675 302772 151676 302836
rect 151740 302772 151741 302836
rect 151675 302771 151741 302772
rect 148918 294541 148978 295155
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 148915 294540 148981 294541
rect 148915 294476 148916 294540
rect 148980 294476 148981 294540
rect 148915 294475 148981 294476
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 147443 3500 147509 3501
rect 147443 3436 147444 3500
rect 147508 3436 147509 3500
rect 147443 3435 147509 3436
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 298894 153854 334338
rect 155171 325140 155237 325141
rect 155171 325076 155172 325140
rect 155236 325076 155237 325140
rect 155171 325075 155237 325076
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 155174 272509 155234 325075
rect 155726 320789 155786 603195
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 162715 588028 162781 588029
rect 162715 587964 162716 588028
rect 162780 587964 162781 588028
rect 162715 587963 162781 587964
rect 159955 565860 160021 565861
rect 159955 565796 159956 565860
rect 160020 565796 160021 565860
rect 159955 565795 160021 565796
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156643 483716 156709 483717
rect 156643 483652 156644 483716
rect 156708 483652 156709 483716
rect 156643 483651 156709 483652
rect 156646 336293 156706 483651
rect 156954 482614 157574 518058
rect 159771 503028 159837 503029
rect 159771 502964 159772 503028
rect 159836 502964 159837 503028
rect 159771 502963 159837 502964
rect 158483 489156 158549 489157
rect 158483 489092 158484 489156
rect 158548 489092 158549 489156
rect 158483 489091 158549 489092
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156643 336292 156709 336293
rect 156643 336228 156644 336292
rect 156708 336228 156709 336292
rect 156643 336227 156709 336228
rect 156646 336021 156706 336227
rect 156643 336020 156709 336021
rect 156643 335956 156644 336020
rect 156708 335956 156709 336020
rect 156643 335955 156709 335956
rect 155723 320788 155789 320789
rect 155723 320724 155724 320788
rect 155788 320724 155789 320788
rect 155723 320723 155789 320724
rect 156954 302614 157574 338058
rect 158486 334661 158546 489091
rect 159774 418845 159834 502963
rect 159771 418844 159837 418845
rect 159771 418780 159772 418844
rect 159836 418780 159837 418844
rect 159771 418779 159837 418780
rect 159771 414628 159837 414629
rect 159771 414564 159772 414628
rect 159836 414564 159837 414628
rect 159771 414563 159837 414564
rect 158483 334660 158549 334661
rect 158483 334596 158484 334660
rect 158548 334596 158549 334660
rect 158483 334595 158549 334596
rect 159774 333437 159834 414563
rect 159771 333436 159837 333437
rect 159771 333372 159772 333436
rect 159836 333372 159837 333436
rect 159771 333371 159837 333372
rect 159219 304332 159285 304333
rect 159219 304268 159220 304332
rect 159284 304268 159285 304332
rect 159219 304267 159285 304268
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 155171 272508 155237 272509
rect 155171 272444 155172 272508
rect 155236 272444 155237 272508
rect 155171 272443 155237 272444
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 159222 25533 159282 304267
rect 159958 260133 160018 565795
rect 161243 559060 161309 559061
rect 161243 558996 161244 559060
rect 161308 558996 161309 559060
rect 161243 558995 161309 558996
rect 161059 428500 161125 428501
rect 161059 428436 161060 428500
rect 161124 428436 161125 428500
rect 161059 428435 161125 428436
rect 160691 339556 160757 339557
rect 160691 339492 160692 339556
rect 160756 339492 160757 339556
rect 160691 339491 160757 339492
rect 160694 312085 160754 339491
rect 160691 312084 160757 312085
rect 160691 312020 160692 312084
rect 160756 312020 160757 312084
rect 160691 312019 160757 312020
rect 159955 260132 160021 260133
rect 159955 260068 159956 260132
rect 160020 260068 160021 260132
rect 159955 260067 160021 260068
rect 161062 234565 161122 428435
rect 161246 339557 161306 558995
rect 162531 479500 162597 479501
rect 162531 479436 162532 479500
rect 162596 479436 162597 479500
rect 162531 479435 162597 479436
rect 162534 351933 162594 479435
rect 162531 351932 162597 351933
rect 162531 351868 162532 351932
rect 162596 351868 162597 351932
rect 162531 351867 162597 351868
rect 161243 339556 161309 339557
rect 161243 339492 161244 339556
rect 161308 339492 161309 339556
rect 161243 339491 161309 339492
rect 162718 323645 162778 587963
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163635 511324 163701 511325
rect 163635 511260 163636 511324
rect 163700 511260 163701 511324
rect 163635 511259 163701 511260
rect 163638 341461 163698 511259
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 170995 596868 171061 596869
rect 170995 596804 170996 596868
rect 171060 596804 171061 596868
rect 170995 596803 171061 596804
rect 168235 588164 168301 588165
rect 168235 588100 168236 588164
rect 168300 588100 168301 588164
rect 168235 588099 168301 588100
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 166211 480860 166277 480861
rect 166211 480796 166212 480860
rect 166276 480796 166277 480860
rect 166211 480795 166277 480796
rect 165475 469844 165541 469845
rect 165475 469780 165476 469844
rect 165540 469780 165541 469844
rect 165475 469779 165541 469780
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163635 341460 163701 341461
rect 163635 341396 163636 341460
rect 163700 341396 163701 341460
rect 163635 341395 163701 341396
rect 162715 323644 162781 323645
rect 162715 323580 162716 323644
rect 162780 323580 162781 323644
rect 162715 323579 162781 323580
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 165478 269789 165538 469779
rect 166214 330581 166274 480795
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 166395 418844 166461 418845
rect 166395 418780 166396 418844
rect 166460 418780 166461 418844
rect 166395 418779 166461 418780
rect 166211 330580 166277 330581
rect 166211 330516 166212 330580
rect 166276 330516 166277 330580
rect 166211 330515 166277 330516
rect 166398 325710 166458 418779
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 166398 325650 166826 325710
rect 166766 313445 166826 325650
rect 166763 313444 166829 313445
rect 166763 313380 166764 313444
rect 166828 313380 166829 313444
rect 166763 313379 166829 313380
rect 166766 285701 166826 313379
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 166947 302428 167013 302429
rect 166947 302364 166948 302428
rect 167012 302364 167013 302428
rect 166947 302363 167013 302364
rect 166950 301613 167010 302363
rect 166947 301612 167013 301613
rect 166947 301548 166948 301612
rect 167012 301548 167013 301612
rect 166947 301547 167013 301548
rect 166763 285700 166829 285701
rect 166763 285636 166764 285700
rect 166828 285636 166829 285700
rect 166763 285635 166829 285636
rect 167514 277174 168134 312618
rect 168238 302429 168298 588099
rect 169339 513364 169405 513365
rect 169339 513300 169340 513364
rect 169404 513300 169405 513364
rect 169339 513299 169405 513300
rect 169342 464405 169402 513299
rect 169523 490516 169589 490517
rect 169523 490452 169524 490516
rect 169588 490452 169589 490516
rect 169523 490451 169589 490452
rect 169339 464404 169405 464405
rect 169339 464340 169340 464404
rect 169404 464340 169405 464404
rect 169339 464339 169405 464340
rect 168971 456244 169037 456245
rect 168971 456180 168972 456244
rect 169036 456180 169037 456244
rect 168971 456179 169037 456180
rect 168235 302428 168301 302429
rect 168235 302364 168236 302428
rect 168300 302364 168301 302428
rect 168235 302363 168301 302364
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 165475 269788 165541 269789
rect 165475 269724 165476 269788
rect 165540 269724 165541 269788
rect 165475 269723 165541 269724
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 160139 234564 160205 234565
rect 160139 234500 160140 234564
rect 160204 234500 160205 234564
rect 160139 234499 160205 234500
rect 161059 234564 161125 234565
rect 161059 234500 161060 234564
rect 161124 234500 161125 234564
rect 161059 234499 161125 234500
rect 160142 233885 160202 234499
rect 160139 233884 160205 233885
rect 160139 233820 160140 233884
rect 160204 233820 160205 233884
rect 160139 233819 160205 233820
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 159219 25532 159285 25533
rect 159219 25468 159220 25532
rect 159284 25468 159285 25532
rect 159219 25467 159285 25468
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 241174 168134 276618
rect 168974 260541 169034 456179
rect 169526 318885 169586 490451
rect 170811 461548 170877 461549
rect 170811 461484 170812 461548
rect 170876 461484 170877 461548
rect 170811 461483 170877 461484
rect 169707 351932 169773 351933
rect 169707 351868 169708 351932
rect 169772 351868 169773 351932
rect 169707 351867 169773 351868
rect 169523 318884 169589 318885
rect 169523 318820 169524 318884
rect 169588 318820 169589 318884
rect 169523 318819 169589 318820
rect 169526 316050 169586 318819
rect 169158 315990 169586 316050
rect 169158 301477 169218 315990
rect 169155 301476 169221 301477
rect 169155 301412 169156 301476
rect 169220 301412 169221 301476
rect 169155 301411 169221 301412
rect 168971 260540 169037 260541
rect 168971 260476 168972 260540
rect 169036 260476 169037 260540
rect 168971 260475 169037 260476
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 169710 237285 169770 351867
rect 170814 319429 170874 461483
rect 170998 386205 171058 596803
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 179275 592788 179341 592789
rect 179275 592724 179276 592788
rect 179340 592724 179341 592788
rect 179275 592723 179341 592724
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 177803 530636 177869 530637
rect 177803 530572 177804 530636
rect 177868 530572 177869 530636
rect 177803 530571 177869 530572
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 172099 489156 172165 489157
rect 172099 489092 172100 489156
rect 172164 489092 172165 489156
rect 172099 489091 172165 489092
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 170995 386204 171061 386205
rect 170995 386140 170996 386204
rect 171060 386140 171061 386204
rect 170995 386139 171061 386140
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 170811 319428 170877 319429
rect 170811 319364 170812 319428
rect 170876 319364 170877 319428
rect 170811 319363 170877 319364
rect 171234 316894 171854 352338
rect 172102 330445 172162 489091
rect 173755 468620 173821 468621
rect 173755 468556 173756 468620
rect 173820 468556 173821 468620
rect 173755 468555 173821 468556
rect 173571 341596 173637 341597
rect 173571 341532 173572 341596
rect 173636 341532 173637 341596
rect 173571 341531 173637 341532
rect 172099 330444 172165 330445
rect 172099 330380 172100 330444
rect 172164 330380 172165 330444
rect 172099 330379 172165 330380
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 173574 253877 173634 341531
rect 173758 337381 173818 468555
rect 174675 467124 174741 467125
rect 174675 467060 174676 467124
rect 174740 467060 174741 467124
rect 174675 467059 174741 467060
rect 173755 337380 173821 337381
rect 173755 337316 173756 337380
rect 173820 337316 173821 337380
rect 173755 337315 173821 337316
rect 174678 258090 174738 467059
rect 173942 258030 174738 258090
rect 174954 464614 175574 500058
rect 176515 476780 176581 476781
rect 176515 476716 176516 476780
rect 176580 476716 176581 476780
rect 176515 476715 176581 476716
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 173942 256053 174002 258030
rect 173939 256052 174005 256053
rect 173939 255988 173940 256052
rect 174004 255988 174005 256052
rect 173939 255987 174005 255988
rect 173571 253876 173637 253877
rect 173571 253812 173572 253876
rect 173636 253812 173637 253876
rect 173571 253811 173637 253812
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 169707 237284 169773 237285
rect 169707 237220 169708 237284
rect 169772 237220 169773 237284
rect 169707 237219 169773 237220
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 173942 46205 174002 255987
rect 174954 248614 175574 284058
rect 176518 270469 176578 476715
rect 177806 398853 177866 530571
rect 179091 454748 179157 454749
rect 179091 454684 179092 454748
rect 179156 454684 179157 454748
rect 179091 454683 179157 454684
rect 177803 398852 177869 398853
rect 177803 398788 177804 398852
rect 177868 398788 177869 398852
rect 177803 398787 177869 398788
rect 179094 351253 179154 454683
rect 179278 413269 179338 592723
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 180195 485892 180261 485893
rect 180195 485828 180196 485892
rect 180260 485828 180261 485892
rect 180195 485827 180261 485828
rect 180011 467804 180077 467805
rect 180011 467740 180012 467804
rect 180076 467740 180077 467804
rect 180011 467739 180077 467740
rect 179275 413268 179341 413269
rect 179275 413204 179276 413268
rect 179340 413204 179341 413268
rect 179275 413203 179341 413204
rect 180014 382397 180074 467739
rect 180198 430677 180258 485827
rect 181483 474060 181549 474061
rect 181483 473996 181484 474060
rect 181548 473996 181549 474060
rect 181483 473995 181549 473996
rect 180195 430676 180261 430677
rect 180195 430612 180196 430676
rect 180260 430612 180261 430676
rect 180195 430611 180261 430612
rect 180563 417484 180629 417485
rect 180563 417420 180564 417484
rect 180628 417420 180629 417484
rect 180563 417419 180629 417420
rect 180011 382396 180077 382397
rect 180011 382332 180012 382396
rect 180076 382332 180077 382396
rect 180011 382331 180077 382332
rect 179091 351252 179157 351253
rect 179091 351188 179092 351252
rect 179156 351188 179157 351252
rect 179091 351187 179157 351188
rect 178539 302564 178605 302565
rect 178539 302500 178540 302564
rect 178604 302500 178605 302564
rect 178539 302499 178605 302500
rect 176515 270468 176581 270469
rect 176515 270404 176516 270468
rect 176580 270404 176581 270468
rect 176515 270403 176581 270404
rect 178542 254013 178602 302499
rect 175779 254012 175845 254013
rect 175779 253948 175780 254012
rect 175844 253948 175845 254012
rect 175779 253947 175845 253948
rect 178539 254012 178605 254013
rect 178539 253948 178540 254012
rect 178604 253948 178605 254012
rect 178539 253947 178605 253948
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 173939 46204 174005 46205
rect 173939 46140 173940 46204
rect 174004 46140 174005 46204
rect 173939 46139 174005 46140
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 68058
rect 175782 40629 175842 253947
rect 180566 242181 180626 417419
rect 181486 370565 181546 473995
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 188291 604620 188357 604621
rect 188291 604556 188292 604620
rect 188356 604556 188357 604620
rect 188291 604555 188357 604556
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 184795 458284 184861 458285
rect 184795 458220 184796 458284
rect 184860 458220 184861 458284
rect 184795 458219 184861 458220
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181483 370564 181549 370565
rect 181483 370500 181484 370564
rect 181548 370500 181549 370564
rect 181483 370499 181549 370500
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 182771 304196 182837 304197
rect 182771 304132 182772 304196
rect 182836 304132 182837 304196
rect 182771 304131 182837 304132
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 180563 242180 180629 242181
rect 180563 242116 180564 242180
rect 180628 242116 180629 242180
rect 180563 242115 180629 242116
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 182774 82109 182834 304131
rect 184798 245717 184858 458219
rect 185514 439174 186134 474618
rect 186819 467260 186885 467261
rect 186819 467196 186820 467260
rect 186884 467196 186885 467260
rect 186819 467195 186885 467196
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185347 305012 185413 305013
rect 185347 304948 185348 305012
rect 185412 304948 185413 305012
rect 185347 304947 185413 304948
rect 185350 291957 185410 304947
rect 185514 295174 186134 330618
rect 186822 305013 186882 467195
rect 188294 446453 188354 604555
rect 189234 586894 189854 622338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 601166 193574 626058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 601166 200414 632898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601166 204134 636618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 601166 207854 604338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 601166 211574 608058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 601166 218414 614898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 601166 222134 618618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 601166 225854 622338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 601166 229574 626058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 601166 236414 632898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601166 240134 636618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 601166 243854 604338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 601166 247574 608058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 601166 254414 614898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 211659 600812 211725 600813
rect 211659 600748 211660 600812
rect 211724 600748 211725 600812
rect 211659 600747 211725 600748
rect 246251 600812 246317 600813
rect 246251 600748 246252 600812
rect 246316 600748 246317 600812
rect 246251 600747 246317 600748
rect 192339 600404 192405 600405
rect 192339 600340 192340 600404
rect 192404 600340 192405 600404
rect 192339 600339 192405 600340
rect 191603 590748 191669 590749
rect 191603 590684 191604 590748
rect 191668 590684 191669 590748
rect 191603 590683 191669 590684
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 191606 575517 191666 590683
rect 191603 575516 191669 575517
rect 191603 575452 191604 575516
rect 191668 575452 191669 575516
rect 191603 575451 191669 575452
rect 192342 570757 192402 600339
rect 197123 599044 197189 599045
rect 197123 598980 197124 599044
rect 197188 598980 197189 599044
rect 197123 598979 197189 598980
rect 203195 599044 203261 599045
rect 203195 598980 203196 599044
rect 203260 598980 203261 599044
rect 203195 598979 203261 598980
rect 207059 599044 207125 599045
rect 207059 598980 207060 599044
rect 207124 598980 207125 599044
rect 207059 598979 207125 598980
rect 210371 599044 210437 599045
rect 210371 598980 210372 599044
rect 210436 598980 210437 599044
rect 210371 598979 210437 598980
rect 193259 598500 193325 598501
rect 193259 598436 193260 598500
rect 193324 598436 193325 598500
rect 193259 598435 193325 598436
rect 193262 589933 193322 598435
rect 193259 589932 193325 589933
rect 193259 589868 193260 589932
rect 193324 589868 193325 589932
rect 193259 589867 193325 589868
rect 193443 575516 193509 575517
rect 193443 575452 193444 575516
rect 193508 575452 193509 575516
rect 193443 575451 193509 575452
rect 192339 570756 192405 570757
rect 192339 570692 192340 570756
rect 192404 570692 192405 570756
rect 192339 570691 192405 570692
rect 193446 567210 193506 575451
rect 193446 567150 193874 567210
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 188843 447404 188909 447405
rect 188843 447340 188844 447404
rect 188908 447340 188909 447404
rect 188843 447339 188909 447340
rect 188291 446452 188357 446453
rect 188291 446388 188292 446452
rect 188356 446388 188357 446452
rect 188291 446387 188357 446388
rect 187555 384436 187621 384437
rect 187555 384372 187556 384436
rect 187620 384372 187621 384436
rect 187555 384371 187621 384372
rect 187558 382261 187618 384371
rect 187555 382260 187621 382261
rect 187555 382196 187556 382260
rect 187620 382196 187621 382260
rect 187555 382195 187621 382196
rect 186819 305012 186885 305013
rect 186819 304948 186820 305012
rect 186884 304948 186885 305012
rect 186819 304947 186885 304948
rect 186267 302564 186333 302565
rect 186267 302500 186268 302564
rect 186332 302500 186333 302564
rect 186267 302499 186333 302500
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185347 291956 185413 291957
rect 185347 291892 185348 291956
rect 185412 291892 185413 291956
rect 185347 291891 185413 291892
rect 185347 274684 185413 274685
rect 185347 274620 185348 274684
rect 185412 274620 185413 274684
rect 185347 274619 185413 274620
rect 184795 245716 184861 245717
rect 184795 245652 184796 245716
rect 184860 245652 184861 245716
rect 184795 245651 184861 245652
rect 185350 205053 185410 274619
rect 185514 259174 186134 294618
rect 186270 285021 186330 302499
rect 186819 296988 186885 296989
rect 186819 296924 186820 296988
rect 186884 296924 186885 296988
rect 186819 296923 186885 296924
rect 186267 285020 186333 285021
rect 186267 284956 186268 285020
rect 186332 284956 186333 285020
rect 186267 284955 186333 284956
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 186822 250477 186882 296923
rect 188846 254149 188906 447339
rect 189234 442894 189854 478338
rect 192954 518614 193574 537166
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 452356 193574 482058
rect 192707 448628 192773 448629
rect 192707 448564 192708 448628
rect 192772 448564 192773 448628
rect 192707 448563 192773 448564
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 192710 378725 192770 448563
rect 192707 378724 192773 378725
rect 192707 378660 192708 378724
rect 192772 378660 192773 378724
rect 192707 378659 192773 378660
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 192954 374614 193574 388356
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 303592 193574 338058
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 193814 275365 193874 567150
rect 197126 493373 197186 598979
rect 197776 579454 198096 579486
rect 197776 579218 197818 579454
rect 198054 579218 198096 579454
rect 197776 579134 198096 579218
rect 197776 578898 197818 579134
rect 198054 578898 198096 579134
rect 197776 578866 198096 578898
rect 197776 543454 198096 543486
rect 197776 543218 197818 543454
rect 198054 543218 198096 543454
rect 197776 543134 198096 543218
rect 197776 542898 197818 543134
rect 198054 542898 198096 543134
rect 197776 542866 198096 542898
rect 199794 525454 200414 537166
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 197123 493372 197189 493373
rect 197123 493308 197124 493372
rect 197188 493308 197189 493372
rect 197123 493307 197189 493308
rect 199794 489454 200414 524898
rect 203198 508469 203258 598979
rect 203514 529174 204134 537166
rect 206139 535532 206205 535533
rect 206139 535468 206140 535532
rect 206204 535468 206205 535532
rect 206139 535467 206205 535468
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203195 508468 203261 508469
rect 203195 508404 203196 508468
rect 203260 508404 203261 508468
rect 203195 508403 203261 508404
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 452356 200414 452898
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 206142 482221 206202 535467
rect 206139 482220 206205 482221
rect 206139 482156 206140 482220
rect 206204 482156 206205 482220
rect 206139 482155 206205 482156
rect 207062 475421 207122 598979
rect 207234 532894 207854 537166
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207059 475420 207125 475421
rect 207059 475356 207060 475420
rect 207124 475356 207125 475420
rect 207059 475355 207125 475356
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 452356 204134 456618
rect 207234 460894 207854 496338
rect 210374 492829 210434 598979
rect 210954 536614 211574 537166
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210371 492828 210437 492829
rect 210371 492764 210372 492828
rect 210436 492764 210437 492828
rect 210371 492763 210437 492764
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 452356 207854 460338
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 452356 211574 464058
rect 211662 462909 211722 600747
rect 219939 600540 220005 600541
rect 219939 600476 219940 600540
rect 220004 600476 220005 600540
rect 219939 600475 220005 600476
rect 229691 600540 229757 600541
rect 229691 600476 229692 600540
rect 229756 600476 229757 600540
rect 229691 600475 229757 600476
rect 237971 600540 238037 600541
rect 237971 600476 237972 600540
rect 238036 600476 238037 600540
rect 237971 600475 238037 600476
rect 215339 600404 215405 600405
rect 215339 600340 215340 600404
rect 215404 600340 215405 600404
rect 215339 600339 215405 600340
rect 213136 561454 213456 561486
rect 213136 561218 213178 561454
rect 213414 561218 213456 561454
rect 213136 561134 213456 561218
rect 213136 560898 213178 561134
rect 213414 560898 213456 561134
rect 213136 560866 213456 560898
rect 215342 483717 215402 600339
rect 216443 599044 216509 599045
rect 216443 598980 216444 599044
rect 216508 598980 216509 599044
rect 216443 598979 216509 598980
rect 216627 599044 216693 599045
rect 216627 598980 216628 599044
rect 216692 598980 216693 599044
rect 216627 598979 216693 598980
rect 218651 599044 218717 599045
rect 218651 598980 218652 599044
rect 218716 598980 218717 599044
rect 218651 598979 218717 598980
rect 216446 493509 216506 598979
rect 216630 509829 216690 598979
rect 216627 509828 216693 509829
rect 216627 509764 216628 509828
rect 216692 509764 216693 509828
rect 216627 509763 216693 509764
rect 217794 507454 218414 537166
rect 218654 512685 218714 598979
rect 219942 522341 220002 600475
rect 226931 600404 226997 600405
rect 226931 600340 226932 600404
rect 226996 600340 226997 600404
rect 226931 600339 226997 600340
rect 222699 599180 222765 599181
rect 222699 599116 222700 599180
rect 222764 599116 222765 599180
rect 222699 599115 222765 599116
rect 223803 599180 223869 599181
rect 223803 599116 223804 599180
rect 223868 599116 223869 599180
rect 223803 599115 223869 599116
rect 220859 599044 220925 599045
rect 220859 598980 220860 599044
rect 220924 598980 220925 599044
rect 220859 598979 220925 598980
rect 219939 522340 220005 522341
rect 219939 522276 219940 522340
rect 220004 522276 220005 522340
rect 219939 522275 220005 522276
rect 218651 512684 218717 512685
rect 218651 512620 218652 512684
rect 218716 512620 218717 512684
rect 218651 512619 218717 512620
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 216443 493508 216509 493509
rect 216443 493444 216444 493508
rect 216508 493444 216509 493508
rect 216443 493443 216509 493444
rect 215339 483716 215405 483717
rect 215339 483652 215340 483716
rect 215404 483652 215405 483716
rect 215339 483651 215405 483652
rect 217794 471454 218414 506898
rect 220862 474061 220922 598979
rect 221514 511174 222134 537166
rect 222702 518125 222762 599115
rect 222699 518124 222765 518125
rect 222699 518060 222700 518124
rect 222764 518060 222765 518124
rect 222699 518059 222765 518060
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 223806 490653 223866 599115
rect 223987 599044 224053 599045
rect 223987 598980 223988 599044
rect 224052 598980 224053 599044
rect 223987 598979 224053 598980
rect 226195 599044 226261 599045
rect 226195 598980 226196 599044
rect 226260 598980 226261 599044
rect 226195 598979 226261 598980
rect 226379 599044 226445 599045
rect 226379 598980 226380 599044
rect 226444 598980 226445 599044
rect 226379 598979 226445 598980
rect 223803 490652 223869 490653
rect 223803 490588 223804 490652
rect 223868 490588 223869 490652
rect 223803 490587 223869 490588
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 220859 474060 220925 474061
rect 220859 473996 220860 474060
rect 220924 473996 220925 474060
rect 220859 473995 220925 473996
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 211659 462908 211725 462909
rect 211659 462844 211660 462908
rect 211724 462844 211725 462908
rect 211659 462843 211725 462844
rect 217794 452356 218414 470898
rect 221514 452356 222134 474618
rect 223990 460325 224050 598979
rect 225234 514894 225854 537166
rect 226198 523701 226258 598979
rect 226195 523700 226261 523701
rect 226195 523636 226196 523700
rect 226260 523636 226261 523700
rect 226195 523635 226261 523636
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 226382 489293 226442 598979
rect 226934 491877 226994 600339
rect 228219 599044 228285 599045
rect 228219 598980 228220 599044
rect 228284 598980 228285 599044
rect 228219 598979 228285 598980
rect 226931 491876 226997 491877
rect 226931 491812 226932 491876
rect 226996 491812 226997 491876
rect 226931 491811 226997 491812
rect 226379 489292 226445 489293
rect 226379 489228 226380 489292
rect 226444 489228 226445 489292
rect 226379 489227 226445 489228
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 223987 460324 224053 460325
rect 223987 460260 223988 460324
rect 224052 460260 224053 460324
rect 223987 460259 224053 460260
rect 225234 452356 225854 478338
rect 228222 458829 228282 598979
rect 228496 579454 228816 579486
rect 228496 579218 228538 579454
rect 228774 579218 228816 579454
rect 228496 579134 228816 579218
rect 228496 578898 228538 579134
rect 228774 578898 228816 579134
rect 228496 578866 228816 578898
rect 228496 543454 228816 543486
rect 228496 543218 228538 543454
rect 228774 543218 228816 543454
rect 228496 543134 228816 543218
rect 228496 542898 228538 543134
rect 228774 542898 228816 543134
rect 228496 542866 228816 542898
rect 228954 518614 229574 537166
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 229694 498813 229754 600475
rect 233003 599044 233069 599045
rect 233003 598980 233004 599044
rect 233068 598980 233069 599044
rect 233003 598979 233069 598980
rect 233187 599044 233253 599045
rect 233187 598980 233188 599044
rect 233252 598980 233253 599044
rect 233187 598979 233253 598980
rect 234659 599044 234725 599045
rect 234659 598980 234660 599044
rect 234724 598980 234725 599044
rect 234659 598979 234725 598980
rect 236499 599044 236565 599045
rect 236499 598980 236500 599044
rect 236564 598980 236565 599044
rect 236499 598979 236565 598980
rect 233006 529141 233066 598979
rect 233003 529140 233069 529141
rect 233003 529076 233004 529140
rect 233068 529076 233069 529140
rect 233003 529075 233069 529076
rect 229691 498812 229757 498813
rect 229691 498748 229692 498812
rect 229756 498748 229757 498812
rect 229691 498747 229757 498748
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228219 458828 228285 458829
rect 228219 458764 228220 458828
rect 228284 458764 228285 458828
rect 228219 458763 228285 458764
rect 228954 452356 229574 482058
rect 233190 458965 233250 598979
rect 234662 478141 234722 598979
rect 235794 525454 236414 537166
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 234659 478140 234725 478141
rect 234659 478076 234660 478140
rect 234724 478076 234725 478140
rect 234659 478075 234725 478076
rect 233187 458964 233253 458965
rect 233187 458900 233188 458964
rect 233252 458900 233253 458964
rect 233187 458899 233253 458900
rect 235794 453454 236414 488898
rect 236502 482221 236562 598979
rect 237974 491197 238034 600475
rect 239259 600404 239325 600405
rect 239259 600340 239260 600404
rect 239324 600340 239325 600404
rect 239259 600339 239325 600340
rect 237971 491196 238037 491197
rect 237971 491132 237972 491196
rect 238036 491132 238037 491196
rect 237971 491131 238037 491132
rect 239262 485077 239322 600339
rect 240731 599044 240797 599045
rect 240731 598980 240732 599044
rect 240796 598980 240797 599044
rect 240731 598979 240797 598980
rect 239514 529174 240134 537166
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239259 485076 239325 485077
rect 239259 485012 239260 485076
rect 239324 485012 239325 485076
rect 239259 485011 239325 485012
rect 236499 482220 236565 482221
rect 236499 482156 236500 482220
rect 236564 482156 236565 482220
rect 236499 482155 236565 482156
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 452356 236414 452898
rect 239514 457174 240134 492618
rect 240734 481541 240794 598979
rect 243856 561454 244176 561486
rect 243856 561218 243898 561454
rect 244134 561218 244176 561454
rect 243856 561134 244176 561218
rect 243856 560898 243898 561134
rect 244134 560898 244176 561134
rect 243856 560866 244176 560898
rect 242939 535532 243005 535533
rect 242939 535468 242940 535532
rect 243004 535468 243005 535532
rect 242939 535467 243005 535468
rect 240731 481540 240797 481541
rect 240731 481476 240732 481540
rect 240796 481476 240797 481540
rect 240731 481475 240797 481476
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 452356 240134 456618
rect 241651 453932 241717 453933
rect 241651 453868 241652 453932
rect 241716 453868 241717 453932
rect 241651 453867 241717 453868
rect 197776 435454 198096 435486
rect 197776 435218 197818 435454
rect 198054 435218 198096 435454
rect 197776 435134 198096 435218
rect 197776 434898 197818 435134
rect 198054 434898 198096 435134
rect 197776 434866 198096 434898
rect 228496 435454 228816 435486
rect 228496 435218 228538 435454
rect 228774 435218 228816 435454
rect 228496 435134 228816 435218
rect 228496 434898 228538 435134
rect 228774 434898 228816 435134
rect 228496 434866 228816 434898
rect 213136 417454 213456 417486
rect 213136 417218 213178 417454
rect 213414 417218 213456 417454
rect 213136 417134 213456 417218
rect 213136 416898 213178 417134
rect 213414 416898 213456 417134
rect 213136 416866 213456 416898
rect 197776 399454 198096 399486
rect 197776 399218 197818 399454
rect 198054 399218 198096 399454
rect 197776 399134 198096 399218
rect 197776 398898 197818 399134
rect 198054 398898 198096 399134
rect 197776 398866 198096 398898
rect 228496 399454 228816 399486
rect 228496 399218 228538 399454
rect 228774 399218 228816 399454
rect 228496 399134 228816 399218
rect 228496 398898 228538 399134
rect 228774 398898 228816 399134
rect 228496 398866 228816 398898
rect 199794 381454 200414 388356
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 194731 308140 194797 308141
rect 194731 308076 194732 308140
rect 194796 308076 194797 308140
rect 194731 308075 194797 308076
rect 194734 300117 194794 308075
rect 199794 303592 200414 308898
rect 203514 385174 204134 388356
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 303592 204134 312618
rect 207234 352894 207854 388356
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 303592 207854 316338
rect 210954 356614 211574 388356
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 303592 211574 320058
rect 217794 363454 218414 388356
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 303592 218414 326898
rect 221514 367174 222134 388356
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 303592 222134 330618
rect 225234 370894 225854 388356
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 303592 225854 334338
rect 228954 374614 229574 388356
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 303592 229574 338058
rect 235794 381454 236414 388356
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 303592 236414 308898
rect 239514 385174 240134 388356
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 241654 377365 241714 453867
rect 241651 377364 241717 377365
rect 241651 377300 241652 377364
rect 241716 377300 241717 377364
rect 241651 377299 241717 377300
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 242942 334661 243002 535467
rect 243234 532894 243854 537166
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 244411 531996 244477 531997
rect 244411 531932 244412 531996
rect 244476 531932 244477 531996
rect 244411 531931 244477 531932
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 452356 243854 460338
rect 243856 417454 244176 417486
rect 243856 417218 243898 417454
rect 244134 417218 244176 417454
rect 243856 417134 244176 417218
rect 243856 416898 243898 417134
rect 244134 416898 244176 417134
rect 243856 416866 244176 416898
rect 244414 389330 244474 531931
rect 245699 523700 245765 523701
rect 245699 523636 245700 523700
rect 245764 523636 245765 523700
rect 245699 523635 245765 523636
rect 244779 500172 244845 500173
rect 244779 500108 244780 500172
rect 244844 500108 244845 500172
rect 244779 500107 244845 500108
rect 244230 389270 244474 389330
rect 244230 389061 244290 389270
rect 244227 389060 244293 389061
rect 244227 388996 244228 389060
rect 244292 388996 244293 389060
rect 244227 388995 244293 388996
rect 243234 352894 243854 388356
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 242939 334660 243005 334661
rect 242939 334596 242940 334660
rect 243004 334596 243005 334660
rect 242939 334595 243005 334596
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 303592 240134 312618
rect 243234 316894 243854 352338
rect 244230 351117 244290 388995
rect 244227 351116 244293 351117
rect 244227 351052 244228 351116
rect 244292 351052 244293 351116
rect 244227 351051 244293 351052
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 303592 243854 316338
rect 244782 301069 244842 500107
rect 245702 460950 245762 523635
rect 246254 466037 246314 600747
rect 247723 599044 247789 599045
rect 247723 598980 247724 599044
rect 247788 598980 247789 599044
rect 247723 598979 247789 598980
rect 251035 599044 251101 599045
rect 251035 598980 251036 599044
rect 251100 598980 251101 599044
rect 251035 598979 251101 598980
rect 252507 599044 252573 599045
rect 252507 598980 252508 599044
rect 252572 598980 252573 599044
rect 252507 598979 252573 598980
rect 246954 536614 247574 537166
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246251 466036 246317 466037
rect 246251 465972 246252 466036
rect 246316 465972 246317 466036
rect 246251 465971 246317 465972
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 245702 460890 245946 460950
rect 245886 450261 245946 460890
rect 246954 452356 247574 464058
rect 247726 456109 247786 598979
rect 249011 531316 249077 531317
rect 249011 531252 249012 531316
rect 249076 531252 249077 531316
rect 249011 531251 249077 531252
rect 249014 516765 249074 531251
rect 249747 529140 249813 529141
rect 249747 529076 249748 529140
rect 249812 529076 249813 529140
rect 249747 529075 249813 529076
rect 249011 516764 249077 516765
rect 249011 516700 249012 516764
rect 249076 516700 249077 516764
rect 249011 516699 249077 516700
rect 249011 481540 249077 481541
rect 249011 481476 249012 481540
rect 249076 481476 249077 481540
rect 249011 481475 249077 481476
rect 247723 456108 247789 456109
rect 247723 456044 247724 456108
rect 247788 456044 247789 456108
rect 247723 456043 247789 456044
rect 245883 450260 245949 450261
rect 245883 450196 245884 450260
rect 245948 450196 245949 450260
rect 245883 450195 245949 450196
rect 245699 449716 245765 449717
rect 245699 449652 245700 449716
rect 245764 449652 245765 449716
rect 245699 449651 245765 449652
rect 245702 337381 245762 449651
rect 245886 359141 245946 450195
rect 247723 449716 247789 449717
rect 247723 449652 247724 449716
rect 247788 449652 247789 449716
rect 247723 449651 247789 449652
rect 245883 359140 245949 359141
rect 245883 359076 245884 359140
rect 245948 359076 245949 359140
rect 245883 359075 245949 359076
rect 246954 356614 247574 388356
rect 247726 364989 247786 449651
rect 249014 390965 249074 481475
rect 249011 390964 249077 390965
rect 249011 390900 249012 390964
rect 249076 390900 249077 390964
rect 249011 390899 249077 390900
rect 248459 381716 248525 381717
rect 248459 381652 248460 381716
rect 248524 381652 248525 381716
rect 248459 381651 248525 381652
rect 247723 364988 247789 364989
rect 247723 364924 247724 364988
rect 247788 364924 247789 364988
rect 247723 364923 247789 364924
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 245699 337380 245765 337381
rect 245699 337316 245700 337380
rect 245764 337316 245765 337380
rect 245699 337315 245765 337316
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 303592 247574 320058
rect 244779 301068 244845 301069
rect 244779 301004 244780 301068
rect 244844 301004 244845 301068
rect 244779 301003 244845 301004
rect 248462 300797 248522 381651
rect 249750 303789 249810 529075
rect 251038 492693 251098 598979
rect 252510 496093 252570 598979
rect 254531 595236 254597 595237
rect 254531 595172 254532 595236
rect 254596 595172 254597 595236
rect 254531 595171 254597 595172
rect 253794 507454 254414 537166
rect 254534 507925 254594 595171
rect 256739 586532 256805 586533
rect 256739 586468 256740 586532
rect 256804 586468 256805 586532
rect 256739 586467 256805 586468
rect 254715 508468 254781 508469
rect 254715 508404 254716 508468
rect 254780 508404 254781 508468
rect 254715 508403 254781 508404
rect 254531 507924 254597 507925
rect 254531 507860 254532 507924
rect 254596 507860 254597 507924
rect 254531 507859 254597 507860
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 252507 496092 252573 496093
rect 252507 496028 252508 496092
rect 252572 496028 252573 496092
rect 252507 496027 252573 496028
rect 252507 493372 252573 493373
rect 252507 493308 252508 493372
rect 252572 493308 252573 493372
rect 252507 493307 252573 493308
rect 251035 492692 251101 492693
rect 251035 492628 251036 492692
rect 251100 492628 251101 492692
rect 251035 492627 251101 492628
rect 252510 422310 252570 493307
rect 253794 471454 254414 506898
rect 254718 489930 254778 508403
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 452356 254414 470898
rect 254534 489870 254778 489930
rect 253979 452164 254045 452165
rect 253979 452100 253980 452164
rect 254044 452100 254045 452164
rect 253979 452099 254045 452100
rect 253982 446181 254042 452099
rect 253979 446180 254045 446181
rect 253979 446116 253980 446180
rect 254044 446116 254045 446180
rect 253979 446115 254045 446116
rect 254534 440469 254594 489870
rect 256555 466716 256621 466717
rect 256555 466652 256556 466716
rect 256620 466652 256621 466716
rect 256555 466651 256621 466652
rect 254531 440468 254597 440469
rect 254531 440404 254532 440468
rect 254596 440404 254597 440468
rect 254531 440403 254597 440404
rect 256558 437613 256618 466651
rect 256555 437612 256621 437613
rect 256555 437548 256556 437612
rect 256620 437548 256621 437612
rect 256555 437547 256621 437548
rect 252510 422250 253122 422310
rect 252875 404836 252941 404837
rect 252875 404772 252876 404836
rect 252940 404772 252941 404836
rect 252875 404771 252941 404772
rect 252878 393330 252938 404771
rect 253062 397357 253122 422250
rect 253059 397356 253125 397357
rect 253059 397292 253060 397356
rect 253124 397292 253125 397356
rect 253059 397291 253125 397292
rect 253979 396948 254045 396949
rect 253979 396884 253980 396948
rect 254044 396884 254045 396948
rect 253979 396883 254045 396884
rect 252694 393270 252938 393330
rect 251035 388516 251101 388517
rect 251035 388452 251036 388516
rect 251100 388452 251101 388516
rect 251035 388451 251101 388452
rect 249747 303788 249813 303789
rect 249747 303724 249748 303788
rect 249812 303724 249813 303788
rect 249747 303723 249813 303724
rect 248459 300796 248525 300797
rect 248459 300732 248460 300796
rect 248524 300732 248525 300796
rect 248459 300731 248525 300732
rect 194731 300116 194797 300117
rect 194731 300052 194732 300116
rect 194796 300052 194797 300116
rect 194731 300051 194797 300052
rect 197776 291454 198096 291486
rect 197776 291218 197818 291454
rect 198054 291218 198096 291454
rect 197776 291134 198096 291218
rect 197776 290898 197818 291134
rect 198054 290898 198096 291134
rect 197776 290866 198096 290898
rect 228496 291454 228816 291486
rect 228496 291218 228538 291454
rect 228774 291218 228816 291454
rect 228496 291134 228816 291218
rect 228496 290898 228538 291134
rect 228774 290898 228816 291134
rect 228496 290866 228816 290898
rect 193811 275364 193877 275365
rect 193811 275300 193812 275364
rect 193876 275300 193877 275364
rect 193811 275299 193877 275300
rect 213136 273454 213456 273486
rect 213136 273218 213178 273454
rect 213414 273218 213456 273454
rect 213136 273134 213456 273218
rect 213136 272898 213178 273134
rect 213414 272898 213456 273134
rect 213136 272866 213456 272898
rect 243856 273454 244176 273486
rect 243856 273218 243898 273454
rect 244134 273218 244176 273454
rect 243856 273134 244176 273218
rect 243856 272898 243898 273134
rect 244134 272898 244176 273134
rect 243856 272866 244176 272898
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 188843 254148 188909 254149
rect 188843 254084 188844 254148
rect 188908 254084 188909 254148
rect 188843 254083 188909 254084
rect 186819 250476 186885 250477
rect 186819 250412 186820 250476
rect 186884 250412 186885 250476
rect 186819 250411 186885 250412
rect 188291 248572 188357 248573
rect 188291 248508 188292 248572
rect 188356 248508 188357 248572
rect 188291 248507 188357 248508
rect 187555 241500 187621 241501
rect 187555 241436 187556 241500
rect 187620 241436 187621 241500
rect 187555 241435 187621 241436
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185347 205052 185413 205053
rect 185347 204988 185348 205052
rect 185412 204988 185413 205052
rect 185347 204987 185413 204988
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 184059 120732 184125 120733
rect 184059 120668 184060 120732
rect 184124 120668 184125 120732
rect 184059 120667 184125 120668
rect 182771 82108 182837 82109
rect 182771 82044 182772 82108
rect 182836 82044 182837 82108
rect 182771 82043 182837 82044
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 175779 40628 175845 40629
rect 175779 40564 175780 40628
rect 175844 40564 175845 40628
rect 175779 40563 175845 40564
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 74898
rect 184062 74493 184122 120667
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 187558 81429 187618 241435
rect 188294 202197 188354 248507
rect 189234 226894 189854 262338
rect 197776 255454 198096 255486
rect 197776 255218 197818 255454
rect 198054 255218 198096 255454
rect 197776 255134 198096 255218
rect 197776 254898 197818 255134
rect 198054 254898 198096 255134
rect 197776 254866 198096 254898
rect 228496 255454 228816 255486
rect 228496 255218 228538 255454
rect 228774 255218 228816 255454
rect 228496 255134 228816 255218
rect 228496 254898 228538 255134
rect 228774 254898 228816 255134
rect 228496 254866 228816 254898
rect 191787 249116 191853 249117
rect 191787 249052 191788 249116
rect 191852 249052 191853 249116
rect 191787 249051 191853 249052
rect 191790 242861 191850 249051
rect 192339 247484 192405 247485
rect 192339 247420 192340 247484
rect 192404 247420 192405 247484
rect 192339 247419 192405 247420
rect 191787 242860 191853 242861
rect 191787 242796 191788 242860
rect 191852 242796 191853 242860
rect 191787 242795 191853 242796
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188291 202196 188357 202197
rect 188291 202132 188292 202196
rect 188356 202132 188357 202196
rect 188291 202131 188357 202132
rect 189234 190894 189854 226338
rect 192342 222053 192402 247419
rect 193443 245852 193509 245853
rect 193443 245788 193444 245852
rect 193508 245850 193509 245852
rect 193508 245790 193874 245850
rect 193508 245788 193509 245790
rect 193443 245787 193509 245788
rect 193259 243540 193325 243541
rect 193259 243476 193260 243540
rect 193324 243476 193325 243540
rect 193259 243475 193325 243476
rect 193262 242045 193322 243475
rect 193259 242044 193325 242045
rect 193259 241980 193260 242044
rect 193324 241980 193325 242044
rect 193259 241979 193325 241980
rect 192954 230614 193574 239592
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 193814 230485 193874 245790
rect 251038 242045 251098 388451
rect 252694 367029 252754 393270
rect 253982 392053 254042 396883
rect 254531 394636 254597 394637
rect 254531 394572 254532 394636
rect 254596 394572 254597 394636
rect 254531 394571 254597 394572
rect 253979 392052 254045 392053
rect 253979 391988 253980 392052
rect 254044 391988 254045 392052
rect 253979 391987 254045 391988
rect 252691 367028 252757 367029
rect 252691 366964 252692 367028
rect 252756 366964 252757 367028
rect 252691 366963 252757 366964
rect 253794 363454 254414 388356
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 252507 330580 252573 330581
rect 252507 330516 252508 330580
rect 252572 330516 252573 330580
rect 252507 330515 252573 330516
rect 252510 268970 252570 330515
rect 253794 327454 254414 362898
rect 254534 345677 254594 394571
rect 254715 392596 254781 392597
rect 254715 392532 254716 392596
rect 254780 392532 254781 392596
rect 254715 392531 254781 392532
rect 254718 388109 254778 392531
rect 254715 388108 254781 388109
rect 254715 388044 254716 388108
rect 254780 388044 254781 388108
rect 254715 388043 254781 388044
rect 256742 362269 256802 586467
rect 257514 583174 258134 618618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 259499 606116 259565 606117
rect 259499 606052 259500 606116
rect 259564 606052 259565 606116
rect 259499 606051 259565 606052
rect 258395 600676 258461 600677
rect 258395 600612 258396 600676
rect 258460 600612 258461 600676
rect 258395 600611 258461 600612
rect 258398 586530 258458 600611
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 256739 362268 256805 362269
rect 256739 362204 256740 362268
rect 256804 362204 256805 362268
rect 256739 362203 256805 362204
rect 254531 345676 254597 345677
rect 254531 345612 254532 345676
rect 254596 345612 254597 345676
rect 254531 345611 254597 345612
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 303592 254414 326898
rect 257514 331174 258134 366618
rect 258214 586470 258458 586530
rect 258214 334250 258274 586470
rect 258395 366348 258461 366349
rect 258395 366284 258396 366348
rect 258460 366284 258461 366348
rect 258395 366283 258461 366284
rect 258398 340890 258458 366283
rect 259502 356693 259562 606051
rect 261234 586894 261854 622338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 266307 594964 266373 594965
rect 266307 594900 266308 594964
rect 266372 594900 266373 594964
rect 266307 594899 266373 594900
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 262259 589388 262325 589389
rect 262259 589324 262260 589388
rect 262324 589324 262325 589388
rect 262259 589323 262325 589324
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 259499 356692 259565 356693
rect 259499 356628 259500 356692
rect 259564 356628 259565 356692
rect 259499 356627 259565 356628
rect 258398 340830 258826 340890
rect 258214 334190 258642 334250
rect 258582 333301 258642 334190
rect 258579 333300 258645 333301
rect 258579 333236 258580 333300
rect 258644 333236 258645 333300
rect 258579 333235 258645 333236
rect 258766 331230 258826 340830
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 256739 317388 256805 317389
rect 256739 317324 256740 317388
rect 256804 317324 256805 317388
rect 256739 317323 256805 317324
rect 252691 301612 252757 301613
rect 252691 301548 252692 301612
rect 252756 301548 252757 301612
rect 252691 301547 252757 301548
rect 252694 273270 252754 301547
rect 256742 298757 256802 317323
rect 256739 298756 256805 298757
rect 256739 298692 256740 298756
rect 256804 298692 256805 298756
rect 256739 298691 256805 298692
rect 257514 295174 258134 330618
rect 258398 331170 258826 331230
rect 261234 334894 261854 370338
rect 262262 363629 262322 589323
rect 263547 580276 263613 580277
rect 263547 580212 263548 580276
rect 263612 580212 263613 580276
rect 263547 580211 263613 580212
rect 262443 536076 262509 536077
rect 262443 536012 262444 536076
rect 262508 536012 262509 536076
rect 262443 536011 262509 536012
rect 262259 363628 262325 363629
rect 262259 363564 262260 363628
rect 262324 363564 262325 363628
rect 262259 363563 262325 363564
rect 262446 349757 262506 536011
rect 262443 349756 262509 349757
rect 262443 349692 262444 349756
rect 262508 349692 262509 349756
rect 262443 349691 262509 349692
rect 263550 340890 263610 580211
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 263731 351796 263797 351797
rect 263731 351732 263732 351796
rect 263796 351732 263797 351796
rect 263731 351731 263797 351732
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 258398 325710 258458 331170
rect 260971 329220 261037 329221
rect 260971 329156 260972 329220
rect 261036 329156 261037 329220
rect 260971 329155 261037 329156
rect 259499 327316 259565 327317
rect 259499 327252 259500 327316
rect 259564 327252 259565 327316
rect 259499 327251 259565 327252
rect 258398 325650 258826 325710
rect 258579 325004 258645 325005
rect 258579 324940 258580 325004
rect 258644 324940 258645 325004
rect 258579 324939 258645 324940
rect 258582 324050 258642 324939
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 252694 273210 253122 273270
rect 252510 268910 252938 268970
rect 252878 265981 252938 268910
rect 252875 265980 252941 265981
rect 252875 265916 252876 265980
rect 252940 265916 252941 265980
rect 252875 265915 252941 265916
rect 253062 263610 253122 273210
rect 252694 263550 253122 263610
rect 251035 242044 251101 242045
rect 251035 241980 251036 242044
rect 251100 241980 251101 242044
rect 251035 241979 251101 241980
rect 251771 242044 251837 242045
rect 251771 241980 251772 242044
rect 251836 241980 251837 242044
rect 251771 241979 251837 241980
rect 199794 237454 200414 239592
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 193811 230484 193877 230485
rect 193811 230420 193812 230484
rect 193876 230420 193877 230484
rect 193811 230419 193877 230420
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192339 222052 192405 222053
rect 192339 221988 192340 222052
rect 192404 221988 192405 222052
rect 192339 221987 192405 221988
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 188291 169012 188357 169013
rect 188291 168948 188292 169012
rect 188356 168948 188357 169012
rect 188291 168947 188357 168948
rect 188294 144805 188354 168947
rect 189234 154894 189854 190338
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 189947 174588 190013 174589
rect 189947 174524 189948 174588
rect 190012 174524 190013 174588
rect 189947 174523 190013 174524
rect 189950 164389 190010 174523
rect 189947 164388 190013 164389
rect 189947 164324 189948 164388
rect 190012 164324 190013 164388
rect 189947 164323 190013 164324
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 188291 144804 188357 144805
rect 188291 144740 188292 144804
rect 188356 144740 188357 144804
rect 188291 144739 188357 144740
rect 189234 118894 189854 154338
rect 189950 132565 190010 164323
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192339 149156 192405 149157
rect 192339 149092 192340 149156
rect 192404 149092 192405 149156
rect 192339 149091 192405 149092
rect 192342 146301 192402 149091
rect 192339 146300 192405 146301
rect 192339 146236 192340 146300
rect 192404 146236 192405 146300
rect 192339 146235 192405 146236
rect 192342 142170 192402 146235
rect 192954 143035 193574 158058
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 193995 153916 194061 153917
rect 193995 153852 193996 153916
rect 194060 153852 194061 153916
rect 193995 153851 194061 153852
rect 193259 142900 193325 142901
rect 193259 142836 193260 142900
rect 193324 142836 193325 142900
rect 193259 142835 193325 142836
rect 192342 142110 192770 142170
rect 189947 132564 190013 132565
rect 189947 132500 189948 132564
rect 190012 132500 190013 132564
rect 189947 132499 190013 132500
rect 192710 123861 192770 142110
rect 193262 138685 193322 142835
rect 193259 138684 193325 138685
rect 193259 138620 193260 138684
rect 193324 138620 193325 138684
rect 193259 138619 193325 138620
rect 193998 132510 194058 153851
rect 194547 148340 194613 148341
rect 194547 148276 194548 148340
rect 194612 148276 194613 148340
rect 194547 148275 194613 148276
rect 194550 139090 194610 148275
rect 199794 143035 200414 164898
rect 203514 205174 204134 239592
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 200619 157996 200685 157997
rect 200619 157932 200620 157996
rect 200684 157932 200685 157996
rect 200619 157931 200685 157932
rect 197859 142220 197925 142221
rect 197859 142156 197860 142220
rect 197924 142156 197925 142220
rect 197859 142155 197925 142156
rect 196571 140452 196637 140453
rect 196571 140388 196572 140452
rect 196636 140388 196637 140452
rect 196571 140387 196637 140388
rect 194182 139030 194610 139090
rect 194182 138821 194242 139030
rect 194179 138820 194245 138821
rect 194179 138756 194180 138820
rect 194244 138756 194245 138820
rect 194179 138755 194245 138756
rect 193446 132450 194058 132510
rect 193446 124133 193506 132450
rect 193811 131476 193877 131477
rect 193811 131412 193812 131476
rect 193876 131412 193877 131476
rect 193811 131411 193877 131412
rect 193443 124132 193509 124133
rect 193443 124068 193444 124132
rect 193508 124068 193509 124132
rect 193443 124067 193509 124068
rect 192707 123860 192773 123861
rect 192707 123796 192708 123860
rect 192772 123796 192773 123860
rect 192707 123795 192773 123796
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 188291 96660 188357 96661
rect 188291 96596 188292 96660
rect 188356 96596 188357 96660
rect 188291 96595 188357 96596
rect 188294 89453 188354 96595
rect 188475 96116 188541 96117
rect 188475 96052 188476 96116
rect 188540 96052 188541 96116
rect 188475 96051 188541 96052
rect 188478 91221 188538 96051
rect 188475 91220 188541 91221
rect 188475 91156 188476 91220
rect 188540 91156 188541 91220
rect 188475 91155 188541 91156
rect 188291 89452 188357 89453
rect 188291 89388 188292 89452
rect 188356 89388 188357 89452
rect 188291 89387 188357 89388
rect 189234 82894 189854 118338
rect 192710 87549 192770 123795
rect 192707 87548 192773 87549
rect 192707 87484 192708 87548
rect 192772 87484 192773 87548
rect 192707 87483 192773 87484
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 187555 81428 187621 81429
rect 187555 81364 187556 81428
rect 187620 81364 187621 81428
rect 187555 81363 187621 81364
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 184059 74492 184125 74493
rect 184059 74428 184060 74492
rect 184124 74428 184125 74492
rect 184059 74427 184125 74428
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 86614 193574 90782
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 193814 80749 193874 131411
rect 193811 80748 193877 80749
rect 193811 80684 193812 80748
rect 193876 80684 193877 80748
rect 193811 80683 193877 80684
rect 196574 79525 196634 140387
rect 196571 79524 196637 79525
rect 196571 79460 196572 79524
rect 196636 79460 196637 79524
rect 196571 79459 196637 79460
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 197862 26893 197922 142155
rect 199388 111454 199708 111486
rect 199388 111218 199430 111454
rect 199666 111218 199708 111454
rect 199388 111134 199708 111218
rect 199388 110898 199430 111134
rect 199666 110898 199708 111134
rect 199388 110866 199708 110898
rect 200622 93397 200682 157931
rect 203514 143035 204134 168618
rect 207234 208894 207854 239592
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 205587 158132 205653 158133
rect 205587 158068 205588 158132
rect 205652 158068 205653 158132
rect 205587 158067 205653 158068
rect 203195 140452 203261 140453
rect 203195 140388 203196 140452
rect 203260 140388 203261 140452
rect 203195 140387 203261 140388
rect 200619 93396 200685 93397
rect 200619 93332 200620 93396
rect 200684 93332 200685 93396
rect 200619 93331 200685 93332
rect 199794 57454 200414 90782
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 197859 26892 197925 26893
rect 197859 26828 197860 26892
rect 197924 26828 197925 26892
rect 197859 26827 197925 26828
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 203198 21317 203258 140387
rect 204264 129454 204584 129486
rect 204264 129218 204306 129454
rect 204542 129218 204584 129454
rect 204264 129134 204584 129218
rect 204264 128898 204306 129134
rect 204542 128898 204584 129134
rect 204264 128866 204584 128898
rect 205590 93397 205650 158067
rect 207234 143035 207854 172338
rect 210954 212614 211574 239592
rect 213131 229940 213197 229941
rect 213131 229876 213132 229940
rect 213196 229876 213197 229940
rect 213131 229875 213197 229876
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 209819 155956 209885 155957
rect 209819 155892 209820 155956
rect 209884 155892 209885 155956
rect 209819 155891 209885 155892
rect 208163 140452 208229 140453
rect 208163 140388 208164 140452
rect 208228 140388 208229 140452
rect 208163 140387 208229 140388
rect 205587 93396 205653 93397
rect 205587 93332 205588 93396
rect 205652 93332 205653 93396
rect 205587 93331 205653 93332
rect 203514 61174 204134 90782
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203195 21316 203261 21317
rect 203195 21252 203196 21316
rect 203260 21252 203261 21316
rect 203195 21251 203261 21252
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 90782
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 208166 39269 208226 140387
rect 209140 111454 209460 111486
rect 209140 111218 209182 111454
rect 209418 111218 209460 111454
rect 209140 111134 209460 111218
rect 209140 110898 209182 111134
rect 209418 110898 209460 111134
rect 209140 110866 209460 110898
rect 209822 92309 209882 155891
rect 210954 143035 211574 176058
rect 211659 163436 211725 163437
rect 211659 163372 211660 163436
rect 211724 163372 211725 163436
rect 211659 163371 211725 163372
rect 210003 140588 210069 140589
rect 210003 140524 210004 140588
rect 210068 140524 210069 140588
rect 210003 140523 210069 140524
rect 210006 93397 210066 140523
rect 211662 93397 211722 163371
rect 210003 93396 210069 93397
rect 210003 93332 210004 93396
rect 210068 93332 210069 93396
rect 210003 93331 210069 93332
rect 211659 93396 211725 93397
rect 211659 93332 211660 93396
rect 211724 93332 211725 93396
rect 211659 93331 211725 93332
rect 213134 92989 213194 229875
rect 215339 224228 215405 224229
rect 215339 224164 215340 224228
rect 215404 224164 215405 224228
rect 215339 224163 215405 224164
rect 214016 129454 214336 129486
rect 214016 129218 214058 129454
rect 214294 129218 214336 129454
rect 214016 129134 214336 129218
rect 214016 128898 214058 129134
rect 214294 128898 214336 129134
rect 214016 128866 214336 128898
rect 213131 92988 213197 92989
rect 213131 92924 213132 92988
rect 213196 92924 213197 92988
rect 213131 92923 213197 92924
rect 209819 92308 209885 92309
rect 209819 92244 209820 92308
rect 209884 92244 209885 92308
rect 209819 92243 209885 92244
rect 210954 68614 211574 90782
rect 215342 90269 215402 224163
rect 217794 219454 218414 239592
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 143035 218414 146898
rect 221514 223174 222134 239592
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 225234 226894 225854 239592
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 223619 192540 223685 192541
rect 223619 192476 223620 192540
rect 223684 192476 223685 192540
rect 223619 192475 223685 192476
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 143035 222134 150618
rect 223622 143581 223682 192475
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 228954 230614 229574 239592
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 226379 182884 226445 182885
rect 226379 182820 226380 182884
rect 226444 182820 226445 182884
rect 226379 182819 226445 182820
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 224355 143716 224421 143717
rect 224355 143652 224356 143716
rect 224420 143652 224421 143716
rect 224355 143651 224421 143652
rect 223619 143580 223685 143581
rect 223619 143516 223620 143580
rect 223684 143516 223685 143580
rect 223619 143515 223685 143516
rect 223622 132510 223682 143515
rect 224358 133381 224418 143651
rect 225234 143035 225854 154338
rect 224907 141132 224973 141133
rect 224907 141068 224908 141132
rect 224972 141068 224973 141132
rect 224907 141067 224973 141068
rect 224355 133380 224421 133381
rect 224355 133316 224356 133380
rect 224420 133316 224421 133380
rect 224355 133315 224421 133316
rect 223622 132450 224418 132510
rect 224358 129709 224418 132450
rect 224355 129708 224421 129709
rect 224355 129644 224356 129708
rect 224420 129644 224421 129708
rect 224355 129643 224421 129644
rect 224910 120053 224970 141067
rect 226382 134741 226442 182819
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 227667 151060 227733 151061
rect 227667 150996 227668 151060
rect 227732 150996 227733 151060
rect 227667 150995 227733 150996
rect 226379 134740 226445 134741
rect 226379 134676 226380 134740
rect 226444 134676 226445 134740
rect 226379 134675 226445 134676
rect 227670 121141 227730 150995
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 227667 121140 227733 121141
rect 227667 121076 227668 121140
rect 227732 121076 227733 121140
rect 227667 121075 227733 121076
rect 224907 120052 224973 120053
rect 224907 119988 224908 120052
rect 224972 119988 224973 120052
rect 224907 119987 224973 119988
rect 218892 111454 219212 111486
rect 218892 111218 218934 111454
rect 219170 111218 219212 111454
rect 218892 111134 219212 111218
rect 218892 110898 218934 111134
rect 219170 110898 219212 111134
rect 218892 110866 219212 110898
rect 226379 107812 226445 107813
rect 226379 107748 226380 107812
rect 226444 107748 226445 107812
rect 226379 107747 226445 107748
rect 224723 97476 224789 97477
rect 224723 97412 224724 97476
rect 224788 97412 224789 97476
rect 224723 97411 224789 97412
rect 224355 95844 224421 95845
rect 224355 95780 224356 95844
rect 224420 95780 224421 95844
rect 224355 95779 224421 95780
rect 224358 92853 224418 95779
rect 224726 93397 224786 97411
rect 224723 93396 224789 93397
rect 224723 93332 224724 93396
rect 224788 93332 224789 93396
rect 224723 93331 224789 93332
rect 224355 92852 224421 92853
rect 224355 92788 224356 92852
rect 224420 92788 224421 92852
rect 224355 92787 224421 92788
rect 215339 90268 215405 90269
rect 215339 90204 215340 90268
rect 215404 90204 215405 90268
rect 215339 90203 215405 90204
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 208163 39268 208229 39269
rect 208163 39204 208164 39268
rect 208228 39204 208229 39268
rect 208163 39203 208229 39204
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 90782
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 90782
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 90782
rect 226382 84149 226442 107747
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 226379 84148 226445 84149
rect 226379 84084 226380 84148
rect 226444 84084 226445 84148
rect 226379 84083 226445 84084
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 237454 236414 239592
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 205174 240134 239592
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 208894 243854 239592
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 212614 247574 239592
rect 251774 230077 251834 241979
rect 251771 230076 251837 230077
rect 251771 230012 251772 230076
rect 251836 230012 251837 230076
rect 251771 230011 251837 230012
rect 252694 229941 252754 263550
rect 257514 259174 258134 294618
rect 258214 323990 258642 324050
rect 258214 290050 258274 323990
rect 258766 320650 258826 325650
rect 258398 320590 258826 320650
rect 258398 299490 258458 320590
rect 258398 299430 258826 299490
rect 258579 290052 258645 290053
rect 258579 290050 258580 290052
rect 258214 289990 258580 290050
rect 258579 289988 258580 289990
rect 258644 289988 258645 290052
rect 258579 289987 258645 289988
rect 258766 289830 258826 299430
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 258398 289770 258826 289830
rect 258398 258909 258458 289770
rect 259502 288829 259562 327251
rect 259683 307188 259749 307189
rect 259683 307124 259684 307188
rect 259748 307124 259749 307188
rect 259683 307123 259749 307124
rect 259686 296717 259746 307123
rect 259683 296716 259749 296717
rect 259683 296652 259684 296716
rect 259748 296652 259749 296716
rect 259683 296651 259749 296652
rect 260974 291685 261034 329155
rect 261234 298894 261854 334338
rect 263366 340830 263610 340890
rect 263366 331230 263426 340830
rect 263366 331170 263610 331230
rect 263550 330445 263610 331170
rect 263547 330444 263613 330445
rect 263547 330380 263548 330444
rect 263612 330380 263613 330444
rect 263547 330379 263613 330380
rect 262443 304196 262509 304197
rect 262443 304132 262444 304196
rect 262508 304132 262509 304196
rect 262443 304131 262509 304132
rect 262259 303652 262325 303653
rect 262259 303588 262260 303652
rect 262324 303588 262325 303652
rect 262259 303587 262325 303588
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 260971 291684 261037 291685
rect 260971 291620 260972 291684
rect 261036 291620 261037 291684
rect 260971 291619 261037 291620
rect 260974 291277 261034 291619
rect 260971 291276 261037 291277
rect 260971 291212 260972 291276
rect 261036 291212 261037 291276
rect 260971 291211 261037 291212
rect 259499 288828 259565 288829
rect 259499 288764 259500 288828
rect 259564 288764 259565 288828
rect 259499 288763 259565 288764
rect 260971 267068 261037 267069
rect 260971 267004 260972 267068
rect 261036 267004 261037 267068
rect 260971 267003 261037 267004
rect 260974 260541 261034 267003
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 260971 260540 261037 260541
rect 260971 260476 260972 260540
rect 261036 260476 261037 260540
rect 260971 260475 261037 260476
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 258395 258908 258461 258909
rect 258395 258844 258396 258908
rect 258460 258844 258461 258908
rect 258395 258843 258461 258844
rect 256739 253740 256805 253741
rect 256739 253676 256740 253740
rect 256804 253676 256805 253740
rect 256739 253675 256805 253676
rect 256742 245717 256802 253675
rect 254531 245716 254597 245717
rect 254531 245652 254532 245716
rect 254596 245652 254597 245716
rect 254531 245651 254597 245652
rect 256739 245716 256805 245717
rect 256739 245652 256740 245716
rect 256804 245652 256805 245716
rect 256739 245651 256805 245652
rect 253611 243268 253677 243269
rect 253611 243204 253612 243268
rect 253676 243204 253677 243268
rect 253611 243203 253677 243204
rect 253614 240957 253674 243203
rect 253611 240956 253677 240957
rect 253611 240892 253612 240956
rect 253676 240892 253677 240956
rect 253611 240891 253677 240892
rect 254534 239733 254594 245651
rect 256739 243404 256805 243405
rect 256739 243340 256740 243404
rect 256804 243340 256805 243404
rect 256739 243339 256805 243340
rect 254531 239732 254597 239733
rect 254531 239668 254532 239732
rect 254596 239668 254597 239732
rect 254531 239667 254597 239668
rect 252691 229940 252757 229941
rect 252691 229876 252692 229940
rect 252756 229876 252757 229940
rect 252691 229875 252757 229876
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 219454 254414 239592
rect 256742 237285 256802 243339
rect 256739 237284 256805 237285
rect 256739 237220 256740 237284
rect 256804 237220 256805 237284
rect 256739 237219 256805 237220
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 223174 258134 258618
rect 258398 258090 258458 258843
rect 258214 258030 258458 258090
rect 258214 248430 258274 258030
rect 258214 248370 258458 248430
rect 258398 241501 258458 248370
rect 259499 246396 259565 246397
rect 259499 246332 259500 246396
rect 259564 246332 259565 246396
rect 259499 246331 259565 246332
rect 258395 241500 258461 241501
rect 258395 241436 258396 241500
rect 258460 241436 258461 241500
rect 258395 241435 258461 241436
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 259502 217293 259562 246331
rect 260974 231165 261034 260475
rect 260971 231164 261037 231165
rect 260971 231100 260972 231164
rect 261036 231100 261037 231164
rect 260971 231099 261037 231100
rect 261234 226894 261854 262338
rect 262262 235245 262322 303587
rect 262446 265573 262506 304131
rect 263734 270469 263794 351731
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 263915 330716 263981 330717
rect 263915 330652 263916 330716
rect 263980 330652 263981 330716
rect 263915 330651 263981 330652
rect 263731 270468 263797 270469
rect 263731 270404 263732 270468
rect 263796 270404 263797 270468
rect 263731 270403 263797 270404
rect 262443 265572 262509 265573
rect 262443 265508 262444 265572
rect 262508 265508 262509 265572
rect 262443 265507 262509 265508
rect 262446 265165 262506 265507
rect 262443 265164 262509 265165
rect 262443 265100 262444 265164
rect 262508 265100 262509 265164
rect 262443 265099 262509 265100
rect 263918 262717 263978 330651
rect 264954 302614 265574 338058
rect 265755 325820 265821 325821
rect 265755 325756 265756 325820
rect 265820 325756 265821 325820
rect 265755 325755 265821 325756
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 265758 267750 265818 325755
rect 266310 312085 266370 594899
rect 267779 578372 267845 578373
rect 267779 578308 267780 578372
rect 267844 578308 267845 578372
rect 267779 578307 267845 578308
rect 267782 334117 267842 578307
rect 267963 563412 268029 563413
rect 267963 563348 267964 563412
rect 268028 563348 268029 563412
rect 267963 563347 268029 563348
rect 267966 345813 268026 563347
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 269067 559060 269133 559061
rect 269067 558996 269068 559060
rect 269132 558996 269133 559060
rect 269067 558995 269133 558996
rect 267963 345812 268029 345813
rect 267963 345748 267964 345812
rect 268028 345748 268029 345812
rect 267963 345747 268029 345748
rect 269070 344317 269130 558995
rect 270539 542740 270605 542741
rect 270539 542676 270540 542740
rect 270604 542676 270605 542740
rect 270539 542675 270605 542676
rect 269067 344316 269133 344317
rect 269067 344252 269068 344316
rect 269132 344252 269133 344316
rect 269067 344251 269133 344252
rect 268331 341460 268397 341461
rect 268331 341396 268332 341460
rect 268396 341396 268397 341460
rect 268331 341395 268397 341396
rect 267963 334660 268029 334661
rect 267963 334596 267964 334660
rect 268028 334596 268029 334660
rect 267963 334595 268029 334596
rect 267779 334116 267845 334117
rect 267779 334052 267780 334116
rect 267844 334052 267845 334116
rect 267779 334051 267845 334052
rect 267966 316050 268026 334595
rect 267782 315990 268026 316050
rect 266307 312084 266373 312085
rect 266307 312020 266308 312084
rect 266372 312020 266373 312084
rect 266307 312019 266373 312020
rect 265758 267690 266002 267750
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 263915 262716 263981 262717
rect 263915 262652 263916 262716
rect 263980 262652 263981 262716
rect 263915 262651 263981 262652
rect 263547 261492 263613 261493
rect 263547 261428 263548 261492
rect 263612 261428 263613 261492
rect 263547 261427 263613 261428
rect 263550 261085 263610 261427
rect 263547 261084 263613 261085
rect 263547 261020 263548 261084
rect 263612 261020 263613 261084
rect 263547 261019 263613 261020
rect 262443 257276 262509 257277
rect 262443 257212 262444 257276
rect 262508 257212 262509 257276
rect 262443 257211 262509 257212
rect 262259 235244 262325 235245
rect 262259 235180 262260 235244
rect 262324 235180 262325 235244
rect 262259 235179 262325 235180
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 259499 217292 259565 217293
rect 259499 217228 259500 217292
rect 259564 217228 259565 217292
rect 259499 217227 259565 217228
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 190894 261854 226338
rect 262446 222189 262506 257211
rect 262443 222188 262509 222189
rect 262443 222124 262444 222188
rect 262508 222124 262509 222188
rect 262443 222123 262509 222124
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 263550 189685 263610 261019
rect 263731 259996 263797 259997
rect 263731 259932 263732 259996
rect 263796 259932 263797 259996
rect 263731 259931 263797 259932
rect 263734 229805 263794 259931
rect 264954 230614 265574 266058
rect 265942 252517 266002 267690
rect 265939 252516 266005 252517
rect 265939 252452 265940 252516
rect 266004 252452 266005 252516
rect 265939 252451 266005 252452
rect 265755 252108 265821 252109
rect 265755 252044 265756 252108
rect 265820 252044 265821 252108
rect 265755 252043 265821 252044
rect 265758 234565 265818 252043
rect 266310 236741 266370 312019
rect 266491 311404 266557 311405
rect 266491 311340 266492 311404
rect 266556 311340 266557 311404
rect 266491 311339 266557 311340
rect 266494 247757 266554 311339
rect 266491 247756 266557 247757
rect 266491 247692 266492 247756
rect 266556 247692 266557 247756
rect 266491 247691 266557 247692
rect 266307 236740 266373 236741
rect 266307 236676 266308 236740
rect 266372 236676 266373 236740
rect 266307 236675 266373 236676
rect 265755 234564 265821 234565
rect 265755 234500 265756 234564
rect 265820 234500 265821 234564
rect 265755 234499 265821 234500
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 263731 229804 263797 229805
rect 263731 229740 263732 229804
rect 263796 229740 263797 229804
rect 263731 229739 263797 229740
rect 264954 194614 265574 230058
rect 266494 219333 266554 247691
rect 267782 244221 267842 315990
rect 268334 286109 268394 341395
rect 269067 319428 269133 319429
rect 269067 319364 269068 319428
rect 269132 319364 269133 319428
rect 269067 319363 269133 319364
rect 268331 286108 268397 286109
rect 268331 286044 268332 286108
rect 268396 286044 268397 286108
rect 268331 286043 268397 286044
rect 268334 285837 268394 286043
rect 268331 285836 268397 285837
rect 268331 285772 268332 285836
rect 268396 285772 268397 285836
rect 268331 285771 268397 285772
rect 267963 250068 268029 250069
rect 267963 250004 267964 250068
rect 268028 250004 268029 250068
rect 267963 250003 268029 250004
rect 267779 244220 267845 244221
rect 267779 244156 267780 244220
rect 267844 244156 267845 244220
rect 267779 244155 267845 244156
rect 267966 231845 268026 250003
rect 269070 242317 269130 319363
rect 270542 313989 270602 542675
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 280291 584084 280357 584085
rect 280291 584020 280292 584084
rect 280356 584020 280357 584084
rect 280291 584019 280357 584020
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 276243 539748 276309 539749
rect 276243 539684 276244 539748
rect 276308 539684 276309 539748
rect 276243 539683 276309 539684
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 273483 465084 273549 465085
rect 273483 465020 273484 465084
rect 273548 465020 273549 465084
rect 273483 465019 273549 465020
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271091 447812 271157 447813
rect 271091 447748 271092 447812
rect 271156 447748 271157 447812
rect 271091 447747 271157 447748
rect 271094 385661 271154 447747
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271091 385660 271157 385661
rect 271091 385596 271092 385660
rect 271156 385596 271157 385660
rect 271091 385595 271157 385596
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 270723 364988 270789 364989
rect 270723 364924 270724 364988
rect 270788 364924 270789 364988
rect 270723 364923 270789 364924
rect 270539 313988 270605 313989
rect 270539 313924 270540 313988
rect 270604 313924 270605 313988
rect 270539 313923 270605 313924
rect 270726 262445 270786 364923
rect 271794 345454 272414 380898
rect 273299 378996 273365 378997
rect 273299 378932 273300 378996
rect 273364 378932 273365 378996
rect 273299 378931 273365 378932
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 273115 298212 273181 298213
rect 273115 298148 273116 298212
rect 273180 298148 273181 298212
rect 273115 298147 273181 298148
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 270723 262444 270789 262445
rect 270723 262380 270724 262444
rect 270788 262380 270789 262444
rect 270723 262379 270789 262380
rect 271091 259452 271157 259453
rect 271091 259388 271092 259452
rect 271156 259388 271157 259452
rect 271091 259387 271157 259388
rect 271094 258365 271154 259387
rect 271091 258364 271157 258365
rect 271091 258300 271092 258364
rect 271156 258300 271157 258364
rect 271091 258299 271157 258300
rect 269619 244220 269685 244221
rect 269619 244156 269620 244220
rect 269684 244156 269685 244220
rect 269619 244155 269685 244156
rect 269067 242316 269133 242317
rect 269067 242252 269068 242316
rect 269132 242252 269133 242316
rect 269067 242251 269133 242252
rect 267963 231844 268029 231845
rect 267963 231780 267964 231844
rect 268028 231780 268029 231844
rect 267963 231779 268029 231780
rect 266491 219332 266557 219333
rect 266491 219268 266492 219332
rect 266556 219268 266557 219332
rect 266491 219267 266557 219268
rect 269622 210901 269682 244155
rect 271094 222189 271154 258299
rect 271794 237454 272414 272898
rect 273118 251157 273178 298147
rect 273302 260269 273362 378931
rect 273486 356829 273546 465019
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 273483 356828 273549 356829
rect 273483 356764 273484 356828
rect 273548 356764 273549 356828
rect 273483 356763 273549 356764
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 276246 316709 276306 539683
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 277163 452708 277229 452709
rect 277163 452644 277164 452708
rect 277228 452644 277229 452708
rect 277163 452643 277229 452644
rect 276427 376684 276493 376685
rect 276427 376620 276428 376684
rect 276492 376620 276493 376684
rect 276427 376619 276493 376620
rect 276243 316708 276309 316709
rect 276243 316644 276244 316708
rect 276308 316644 276309 316708
rect 276243 316643 276309 316644
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 276243 285836 276309 285837
rect 276243 285772 276244 285836
rect 276308 285772 276309 285836
rect 276243 285771 276309 285772
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 273667 262172 273733 262173
rect 273667 262108 273668 262172
rect 273732 262108 273733 262172
rect 273667 262107 273733 262108
rect 273670 261221 273730 262107
rect 273667 261220 273733 261221
rect 273667 261156 273668 261220
rect 273732 261156 273733 261220
rect 273667 261155 273733 261156
rect 273299 260268 273365 260269
rect 273299 260204 273300 260268
rect 273364 260204 273365 260268
rect 273299 260203 273365 260204
rect 273115 251156 273181 251157
rect 273115 251092 273116 251156
rect 273180 251092 273181 251156
rect 273115 251091 273181 251092
rect 273118 250610 273178 251091
rect 273118 250550 273546 250610
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271091 222188 271157 222189
rect 271091 222124 271092 222188
rect 271156 222124 271157 222188
rect 271091 222123 271157 222124
rect 269619 210900 269685 210901
rect 269619 210836 269620 210900
rect 269684 210836 269685 210900
rect 269619 210835 269685 210836
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263547 189684 263613 189685
rect 263547 189620 263548 189684
rect 263612 189620 263613 189684
rect 263547 189619 263613 189620
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 201454 272414 236898
rect 273486 235245 273546 250550
rect 273483 235244 273549 235245
rect 273483 235180 273484 235244
rect 273548 235180 273549 235244
rect 273483 235179 273549 235180
rect 273670 203557 273730 261155
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 273667 203556 273733 203557
rect 273667 203492 273668 203556
rect 273732 203492 273733 203556
rect 273667 203491 273733 203492
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 276246 156637 276306 285771
rect 276430 259453 276490 376619
rect 276427 259452 276493 259453
rect 276427 259388 276428 259452
rect 276492 259388 276493 259452
rect 276427 259387 276493 259388
rect 277166 244221 277226 452643
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 280294 383670 280354 584019
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 287099 472156 287165 472157
rect 287099 472092 287100 472156
rect 287164 472092 287165 472156
rect 287099 472091 287165 472092
rect 285627 466580 285693 466581
rect 285627 466516 285628 466580
rect 285692 466516 285693 466580
rect 285627 466515 285693 466516
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 284339 457468 284405 457469
rect 284339 457404 284340 457468
rect 284404 457404 284405 457468
rect 284339 457403 284405 457404
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 281579 416668 281645 416669
rect 281579 416604 281580 416668
rect 281644 416604 281645 416668
rect 281579 416603 281645 416604
rect 280110 383610 280354 383670
rect 280110 355333 280170 383610
rect 280291 380764 280357 380765
rect 280291 380700 280292 380764
rect 280356 380700 280357 380764
rect 280291 380699 280357 380700
rect 280107 355332 280173 355333
rect 280107 355268 280108 355332
rect 280172 355268 280173 355332
rect 280107 355267 280173 355268
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 280294 246397 280354 380699
rect 281582 262853 281642 416603
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 281763 283660 281829 283661
rect 281763 283596 281764 283660
rect 281828 283596 281829 283660
rect 281763 283595 281829 283596
rect 281579 262852 281645 262853
rect 281579 262788 281580 262852
rect 281644 262788 281645 262852
rect 281579 262787 281645 262788
rect 280291 246396 280357 246397
rect 280291 246332 280292 246396
rect 280356 246332 280357 246396
rect 280291 246331 280357 246332
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 277163 244220 277229 244221
rect 277163 244156 277164 244220
rect 277228 244156 277229 244220
rect 277163 244155 277229 244156
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 276243 156636 276309 156637
rect 276243 156572 276244 156636
rect 276308 156572 276309 156636
rect 276243 156571 276309 156572
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 136894 279854 172338
rect 281766 159357 281826 283595
rect 282954 248614 283574 284058
rect 284342 261493 284402 457403
rect 284339 261492 284405 261493
rect 284339 261428 284340 261492
rect 284404 261428 284405 261492
rect 284339 261427 284405 261428
rect 285630 258229 285690 466515
rect 285627 258228 285693 258229
rect 285627 258164 285628 258228
rect 285692 258164 285693 258228
rect 285627 258163 285693 258164
rect 287102 253877 287162 472091
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 288387 378044 288453 378045
rect 288387 377980 288388 378044
rect 288452 377980 288453 378044
rect 288387 377979 288453 377980
rect 288390 267069 288450 377979
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 288387 267068 288453 267069
rect 288387 267004 288388 267068
rect 288452 267004 288453 267068
rect 288387 267003 288453 267004
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 287099 253876 287165 253877
rect 287099 253812 287100 253876
rect 287164 253812 287165 253876
rect 287099 253811 287165 253812
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281763 159356 281829 159357
rect 281763 159292 281764 159356
rect 281828 159292 281829 159356
rect 281763 159291 281829 159292
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 73721 543218 73957 543454
rect 73721 542898 73957 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77686 561218 77922 561454
rect 77686 560898 77922 561134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 74387 255218 74623 255454
rect 74387 254898 74623 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73721 111218 73957 111454
rect 73721 110898 73957 111134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 81651 543218 81887 543454
rect 81651 542898 81887 543134
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 85617 561218 85853 561454
rect 85617 560898 85853 561134
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 79019 273218 79255 273454
rect 79019 272898 79255 273134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 83651 255218 83887 255454
rect 83651 254898 83887 255134
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 89582 543218 89818 543454
rect 89582 542898 89818 543134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 88283 273218 88519 273454
rect 88283 272898 88519 273134
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 92915 255218 93151 255454
rect 92915 254898 93151 255134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 77686 129218 77922 129454
rect 77686 128898 77922 129134
rect 85617 129218 85853 129454
rect 85617 128898 85853 129134
rect 81651 111218 81887 111454
rect 81651 110898 81887 111134
rect 89582 111218 89818 111454
rect 89582 110898 89818 111134
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 197818 579218 198054 579454
rect 197818 578898 198054 579134
rect 197818 543218 198054 543454
rect 197818 542898 198054 543134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 213178 561218 213414 561454
rect 213178 560898 213414 561134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228538 579218 228774 579454
rect 228538 578898 228774 579134
rect 228538 543218 228774 543454
rect 228538 542898 228774 543134
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 243898 561218 244134 561454
rect 243898 560898 244134 561134
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 197818 435218 198054 435454
rect 197818 434898 198054 435134
rect 228538 435218 228774 435454
rect 228538 434898 228774 435134
rect 213178 417218 213414 417454
rect 213178 416898 213414 417134
rect 197818 399218 198054 399454
rect 197818 398898 198054 399134
rect 228538 399218 228774 399454
rect 228538 398898 228774 399134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243898 417218 244134 417454
rect 243898 416898 244134 417134
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 197818 291218 198054 291454
rect 197818 290898 198054 291134
rect 228538 291218 228774 291454
rect 228538 290898 228774 291134
rect 213178 273218 213414 273454
rect 213178 272898 213414 273134
rect 243898 273218 244134 273454
rect 243898 272898 244134 273134
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 197818 255218 198054 255454
rect 197818 254898 198054 255134
rect 228538 255218 228774 255454
rect 228538 254898 228774 255134
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 199430 111218 199666 111454
rect 199430 110898 199666 111134
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 204306 129218 204542 129454
rect 204306 128898 204542 129134
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 209182 111218 209418 111454
rect 209182 110898 209418 111134
rect 214058 129218 214294 129454
rect 214058 128898 214294 129134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 218934 111218 219170 111454
rect 218934 110898 219170 111134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 197818 579454
rect 198054 579218 228538 579454
rect 228774 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 197818 579134
rect 198054 578898 228538 579134
rect 228774 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 77686 561454
rect 77922 561218 85617 561454
rect 85853 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 213178 561454
rect 213414 561218 243898 561454
rect 244134 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 77686 561134
rect 77922 560898 85617 561134
rect 85853 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 213178 561134
rect 213414 560898 243898 561134
rect 244134 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73721 543454
rect 73957 543218 81651 543454
rect 81887 543218 89582 543454
rect 89818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 197818 543454
rect 198054 543218 228538 543454
rect 228774 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73721 543134
rect 73957 542898 81651 543134
rect 81887 542898 89582 543134
rect 89818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 197818 543134
rect 198054 542898 228538 543134
rect 228774 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 197818 435454
rect 198054 435218 228538 435454
rect 228774 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 197818 435134
rect 198054 434898 228538 435134
rect 228774 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 213178 417454
rect 213414 417218 243898 417454
rect 244134 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 213178 417134
rect 213414 416898 243898 417134
rect 244134 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 197818 399454
rect 198054 399218 228538 399454
rect 228774 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 197818 399134
rect 198054 398898 228538 399134
rect 228774 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 197818 291454
rect 198054 291218 228538 291454
rect 228774 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 197818 291134
rect 198054 290898 228538 291134
rect 228774 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 79019 273454
rect 79255 273218 88283 273454
rect 88519 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 213178 273454
rect 213414 273218 243898 273454
rect 244134 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 79019 273134
rect 79255 272898 88283 273134
rect 88519 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 213178 273134
rect 213414 272898 243898 273134
rect 244134 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74387 255454
rect 74623 255218 83651 255454
rect 83887 255218 92915 255454
rect 93151 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 197818 255454
rect 198054 255218 228538 255454
rect 228774 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74387 255134
rect 74623 254898 83651 255134
rect 83887 254898 92915 255134
rect 93151 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 197818 255134
rect 198054 254898 228538 255134
rect 228774 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 77686 129454
rect 77922 129218 85617 129454
rect 85853 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 204306 129454
rect 204542 129218 214058 129454
rect 214294 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 77686 129134
rect 77922 128898 85617 129134
rect 85853 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 204306 129134
rect 204542 128898 214058 129134
rect 214294 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73721 111454
rect 73957 111218 81651 111454
rect 81887 111218 89582 111454
rect 89818 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 199430 111454
rect 199666 111218 209182 111454
rect 209418 111218 218934 111454
rect 219170 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73721 111134
rect 73957 110898 81651 111134
rect 81887 110898 89582 111134
rect 89818 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 199430 111134
rect 199666 110898 209182 111134
rect 209418 110898 218934 111134
rect 219170 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use zube_wrapped_project  zube_wrapped_project_5
timestamp 1636029542
transform 1 0 193568 0 1 241592
box 0 0 60000 60000
use wrapped_ws2812  wrapped_ws2812_4
timestamp 1636029542
transform 1 0 193568 0 1 92782
box 0 0 31475 48253
use wrapped_vga_clock  wrapped_vga_clock_2
timestamp 1636029542
transform 1 0 68770 0 1 390356
box 0 0 44000 44000
use wrapped_tpm2137  wrapped_tpm2137_3
timestamp 1636029542
transform 1 0 68770 0 1 539166
box 0 0 26000 42000
use wrapped_rgb_mixer  wrapped_rgb_mixer_0
timestamp 1636029542
transform 1 0 68770 0 1 92782
box 0 0 26000 42000
use wrapped_nco  wrapped_nco_7
timestamp 1636029542
transform 1 0 193568 0 1 539166
box 0 0 60000 60000
use wrapped_hack_soc  wrapped_hack_soc_6
timestamp 1636029542
transform 1 0 193568 0 1 390356
box 0 0 60000 60000
use wrapped_frequency_counter  wrapped_frequency_counter_1
timestamp 1636029542
transform 1 0 68770 0 1 241592
box 0 0 30000 42000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 136782 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 143035 218414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 303592 218414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 303592 254414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 436356 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 452356 218414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 452356 254414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 583166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 436356 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 601166 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 601166 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 136782 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 143035 222134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 303592 222134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 436356 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 452356 222134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 583166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 436356 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 601166 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 136782 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 143035 225854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 303592 225854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 436356 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 452356 225854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 583166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 601166 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 136782 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 143035 193574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 303592 193574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 303592 229574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 436356 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 452356 193574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 452356 229574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 583166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 601166 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 601166 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 90782 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 143035 207854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 303592 207854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 303592 243854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 452356 207854 537166 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 452356 243854 537166 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 436356 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 601166 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 601166 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 136782 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 143035 211574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 303592 211574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 303592 247574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 436356 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 452356 211574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 452356 247574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 583166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 436356 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 601166 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 601166 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 136782 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 143035 200414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 303592 200414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 303592 236414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 436356 92414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 452356 200414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 452356 236414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 583166 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 601166 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 601166 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 136782 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 143035 204134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 303592 204134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 303592 240134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 436356 96134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 452356 204134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 452356 240134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 583166 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 601166 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 601166 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
