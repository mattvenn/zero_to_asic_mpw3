magic
tech sky130A
magscale 1 2
timestamp 1636115455
<< metal1 >>
rect 242802 703128 242808 703180
rect 242860 703168 242866 703180
rect 348786 703168 348792 703180
rect 242860 703140 348792 703168
rect 242860 703128 242866 703140
rect 348786 703128 348792 703140
rect 348844 703128 348850 703180
rect 268378 703060 268384 703112
rect 268436 703100 268442 703112
rect 413646 703100 413652 703112
rect 268436 703072 413652 703100
rect 268436 703060 268442 703072
rect 413646 703060 413652 703072
rect 413704 703060 413710 703112
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 218974 702992 218980 703044
rect 219032 703032 219038 703044
rect 269114 703032 269120 703044
rect 219032 703004 269120 703032
rect 219032 702992 219038 703004
rect 269114 702992 269120 703004
rect 269172 702992 269178 703044
rect 280798 702992 280804 703044
rect 280856 703032 280862 703044
rect 429838 703032 429844 703044
rect 280856 703004 429844 703032
rect 280856 702992 280862 703004
rect 429838 702992 429844 703004
rect 429896 702992 429902 703044
rect 179322 702924 179328 702976
rect 179380 702964 179386 702976
rect 332502 702964 332508 702976
rect 179380 702936 332508 702964
rect 179380 702924 179386 702936
rect 332502 702924 332508 702936
rect 332560 702924 332566 702976
rect 188338 702856 188344 702908
rect 188396 702896 188402 702908
rect 235166 702896 235172 702908
rect 188396 702868 235172 702896
rect 188396 702856 188402 702868
rect 235166 702856 235172 702868
rect 235224 702856 235230 702908
rect 249702 702856 249708 702908
rect 249760 702896 249766 702908
rect 494790 702896 494796 702908
rect 249760 702868 494796 702896
rect 249760 702856 249766 702868
rect 494790 702856 494796 702868
rect 494848 702856 494854 702908
rect 154114 702788 154120 702840
rect 154172 702828 154178 702840
rect 233234 702828 233240 702840
rect 154172 702800 233240 702828
rect 154172 702788 154178 702800
rect 233234 702788 233240 702800
rect 233292 702788 233298 702840
rect 285582 702788 285588 702840
rect 285640 702828 285646 702840
rect 462314 702828 462320 702840
rect 285640 702800 462320 702828
rect 285640 702788 285646 702800
rect 462314 702788 462320 702800
rect 462372 702788 462378 702840
rect 187602 702720 187608 702772
rect 187660 702760 187666 702772
rect 364978 702760 364984 702772
rect 187660 702732 364984 702760
rect 187660 702720 187666 702732
rect 364978 702720 364984 702732
rect 365036 702720 365042 702772
rect 205634 702652 205640 702704
rect 205692 702692 205698 702704
rect 397362 702692 397368 702704
rect 205692 702664 397368 702692
rect 205692 702652 205698 702664
rect 397362 702652 397368 702664
rect 397420 702652 397426 702704
rect 24302 702584 24308 702636
rect 24360 702624 24366 702636
rect 85574 702624 85580 702636
rect 24360 702596 85580 702624
rect 24360 702584 24366 702596
rect 85574 702584 85580 702596
rect 85632 702584 85638 702636
rect 137830 702584 137836 702636
rect 137888 702624 137894 702636
rect 215294 702624 215300 702636
rect 137888 702596 215300 702624
rect 137888 702584 137894 702596
rect 215294 702584 215300 702596
rect 215352 702584 215358 702636
rect 222838 702584 222844 702636
rect 222896 702624 222902 702636
rect 478506 702624 478512 702636
rect 222896 702596 478512 702624
rect 222896 702584 222902 702596
rect 478506 702584 478512 702596
rect 478564 702584 478570 702636
rect 67634 702516 67640 702568
rect 67692 702556 67698 702568
rect 170306 702556 170312 702568
rect 67692 702528 170312 702556
rect 67692 702516 67698 702528
rect 170306 702516 170312 702528
rect 170364 702556 170370 702568
rect 224218 702556 224224 702568
rect 170364 702528 224224 702556
rect 170364 702516 170370 702528
rect 224218 702516 224224 702528
rect 224276 702516 224282 702568
rect 255958 702516 255964 702568
rect 256016 702556 256022 702568
rect 543458 702556 543464 702568
rect 256016 702528 543464 702556
rect 256016 702516 256022 702528
rect 543458 702516 543464 702528
rect 543516 702516 543522 702568
rect 8110 702448 8116 702500
rect 8168 702488 8174 702500
rect 96614 702488 96620 702500
rect 8168 702460 96620 702488
rect 8168 702448 8174 702460
rect 96614 702448 96620 702460
rect 96672 702448 96678 702500
rect 166350 702448 166356 702500
rect 166408 702488 166414 702500
rect 527174 702488 527180 702500
rect 166408 702460 527180 702488
rect 166408 702448 166414 702460
rect 527174 702448 527180 702460
rect 527232 702448 527238 702500
rect 71038 700272 71044 700324
rect 71096 700312 71102 700324
rect 105446 700312 105452 700324
rect 71096 700284 105452 700312
rect 71096 700272 71102 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 251818 700272 251824 700324
rect 251876 700312 251882 700324
rect 283834 700312 283840 700324
rect 251876 700284 283840 700312
rect 251876 700272 251882 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 559650 700272 559656 700324
rect 559708 700312 559714 700324
rect 582834 700312 582840 700324
rect 559708 700284 582840 700312
rect 559708 700272 559714 700284
rect 582834 700272 582840 700284
rect 582892 700272 582898 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 33778 683176 33784 683188
rect 3476 683148 33784 683176
rect 3476 683136 3482 683148
rect 33778 683136 33784 683148
rect 33836 683136 33842 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 15838 670732 15844 670744
rect 3568 670704 15844 670732
rect 3568 670692 3574 670704
rect 15838 670692 15844 670704
rect 15896 670692 15902 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 74534 656928 74540 656940
rect 3476 656900 74540 656928
rect 3476 656888 3482 656900
rect 74534 656888 74540 656900
rect 74592 656888 74598 656940
rect 81434 620984 81440 621036
rect 81492 621024 81498 621036
rect 201494 621024 201500 621036
rect 81492 620996 201500 621024
rect 81492 620984 81498 620996
rect 201494 620984 201500 620996
rect 201552 621024 201558 621036
rect 202138 621024 202144 621036
rect 201552 620996 202144 621024
rect 201552 620984 201558 620996
rect 202138 620984 202144 620996
rect 202196 620984 202202 621036
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 57238 618304 57244 618316
rect 3568 618276 57244 618304
rect 3568 618264 3574 618276
rect 57238 618264 57244 618276
rect 57296 618264 57302 618316
rect 164142 618264 164148 618316
rect 164200 618304 164206 618316
rect 226334 618304 226340 618316
rect 164200 618276 226340 618304
rect 164200 618264 164206 618276
rect 226334 618264 226340 618276
rect 226392 618264 226398 618316
rect 161382 616836 161388 616888
rect 161440 616876 161446 616888
rect 242894 616876 242900 616888
rect 161440 616848 242900 616876
rect 161440 616836 161446 616848
rect 242894 616836 242900 616848
rect 242952 616836 242958 616888
rect 233234 615952 233240 616004
rect 233292 615992 233298 616004
rect 233878 615992 233884 616004
rect 233292 615964 233884 615992
rect 233292 615952 233298 615964
rect 233878 615952 233884 615964
rect 233936 615952 233942 616004
rect 167638 615544 167644 615596
rect 167696 615584 167702 615596
rect 233234 615584 233240 615596
rect 167696 615556 233240 615584
rect 167696 615544 167702 615556
rect 233234 615544 233240 615556
rect 233292 615544 233298 615596
rect 155586 615476 155592 615528
rect 155644 615516 155650 615528
rect 231854 615516 231860 615528
rect 155644 615488 231860 615516
rect 155644 615476 155650 615488
rect 231854 615476 231860 615488
rect 231912 615476 231918 615528
rect 147582 614184 147588 614236
rect 147640 614224 147646 614236
rect 215938 614224 215944 614236
rect 147640 614196 215944 614224
rect 147640 614184 147646 614196
rect 215938 614184 215944 614196
rect 215996 614184 216002 614236
rect 173802 614116 173808 614168
rect 173860 614156 173866 614168
rect 251910 614156 251916 614168
rect 173860 614128 251916 614156
rect 173860 614116 173866 614128
rect 251910 614116 251916 614128
rect 251968 614116 251974 614168
rect 166258 612824 166264 612876
rect 166316 612864 166322 612876
rect 237466 612864 237472 612876
rect 166316 612836 237472 612864
rect 166316 612824 166322 612836
rect 237466 612824 237472 612836
rect 237524 612824 237530 612876
rect 184290 612756 184296 612808
rect 184348 612796 184354 612808
rect 259454 612796 259460 612808
rect 184348 612768 259460 612796
rect 184348 612756 184354 612768
rect 259454 612756 259460 612768
rect 259512 612756 259518 612808
rect 152550 611396 152556 611448
rect 152608 611436 152614 611448
rect 213178 611436 213184 611448
rect 152608 611408 213184 611436
rect 152608 611396 152614 611408
rect 213178 611396 213184 611408
rect 213236 611396 213242 611448
rect 66162 611328 66168 611380
rect 66220 611368 66226 611380
rect 254118 611368 254124 611380
rect 66220 611340 254124 611368
rect 66220 611328 66226 611340
rect 254118 611328 254124 611340
rect 254176 611328 254182 611380
rect 137922 610036 137928 610088
rect 137980 610076 137986 610088
rect 213086 610076 213092 610088
rect 137980 610048 213092 610076
rect 137980 610036 137986 610048
rect 213086 610036 213092 610048
rect 213144 610036 213150 610088
rect 160738 609968 160744 610020
rect 160796 610008 160802 610020
rect 255314 610008 255320 610020
rect 160796 609980 255320 610008
rect 160796 609968 160802 609980
rect 255314 609968 255320 609980
rect 255372 609968 255378 610020
rect 202138 609288 202144 609340
rect 202196 609328 202202 609340
rect 223022 609328 223028 609340
rect 202196 609300 223028 609328
rect 202196 609288 202202 609300
rect 223022 609288 223028 609300
rect 223080 609288 223086 609340
rect 219342 609220 219348 609272
rect 219400 609260 219406 609272
rect 582834 609260 582840 609272
rect 219400 609232 582840 609260
rect 219400 609220 219406 609232
rect 582834 609220 582840 609232
rect 582892 609220 582898 609272
rect 140682 608608 140688 608660
rect 140740 608648 140746 608660
rect 205726 608648 205732 608660
rect 140740 608620 205732 608648
rect 140740 608608 140746 608620
rect 205726 608608 205732 608620
rect 205784 608608 205790 608660
rect 182818 607248 182824 607300
rect 182876 607288 182882 607300
rect 217686 607288 217692 607300
rect 182876 607260 217692 607288
rect 182876 607248 182882 607260
rect 217686 607248 217692 607260
rect 217744 607248 217750 607300
rect 177298 607180 177304 607232
rect 177356 607220 177362 607232
rect 216950 607220 216956 607232
rect 177356 607192 216956 607220
rect 177356 607180 177362 607192
rect 216950 607180 216956 607192
rect 217008 607180 217014 607232
rect 218790 607180 218796 607232
rect 218848 607220 218854 607232
rect 278038 607220 278044 607232
rect 218848 607192 278044 607220
rect 218848 607180 218854 607192
rect 278038 607180 278044 607192
rect 278096 607180 278102 607232
rect 215938 607112 215944 607164
rect 215996 607152 216002 607164
rect 582374 607152 582380 607164
rect 215996 607124 582380 607152
rect 215996 607112 216002 607124
rect 582374 607112 582380 607124
rect 582432 607112 582438 607164
rect 176562 605888 176568 605940
rect 176620 605928 176626 605940
rect 212534 605928 212540 605940
rect 176620 605900 212540 605928
rect 176620 605888 176626 605900
rect 212534 605888 212540 605900
rect 212592 605888 212598 605940
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 94682 605860 94688 605872
rect 3568 605832 94688 605860
rect 3568 605820 3574 605832
rect 94682 605820 94688 605832
rect 94740 605820 94746 605872
rect 98638 605820 98644 605872
rect 98696 605860 98702 605872
rect 142798 605860 142804 605872
rect 98696 605832 142804 605860
rect 98696 605820 98702 605832
rect 142798 605820 142804 605832
rect 142856 605860 142862 605872
rect 245470 605860 245476 605872
rect 142856 605832 245476 605860
rect 142856 605820 142862 605832
rect 245470 605820 245476 605832
rect 245528 605820 245534 605872
rect 172422 604528 172428 604580
rect 172480 604568 172486 604580
rect 205542 604568 205548 604580
rect 172480 604540 205548 604568
rect 172480 604528 172486 604540
rect 205542 604528 205548 604540
rect 205600 604528 205606 604580
rect 115198 604460 115204 604512
rect 115256 604500 115262 604512
rect 238478 604500 238484 604512
rect 115256 604472 238484 604500
rect 115256 604460 115262 604472
rect 238478 604460 238484 604472
rect 238536 604460 238542 604512
rect 241790 604460 241796 604512
rect 241848 604500 241854 604512
rect 242802 604500 242808 604512
rect 241848 604472 242808 604500
rect 241848 604460 241854 604472
rect 242802 604460 242808 604472
rect 242860 604500 242866 604512
rect 271874 604500 271880 604512
rect 242860 604472 271880 604500
rect 242860 604460 242866 604472
rect 271874 604460 271880 604472
rect 271932 604460 271938 604512
rect 289722 604460 289728 604512
rect 289780 604500 289786 604512
rect 582834 604500 582840 604512
rect 289780 604472 582840 604500
rect 289780 604460 289786 604472
rect 582834 604460 582840 604472
rect 582892 604460 582898 604512
rect 169018 603168 169024 603220
rect 169076 603208 169082 603220
rect 199102 603208 199108 603220
rect 169076 603180 199108 603208
rect 169076 603168 169082 603180
rect 199102 603168 199108 603180
rect 199160 603168 199166 603220
rect 244918 603168 244924 603220
rect 244976 603208 244982 603220
rect 254670 603208 254676 603220
rect 244976 603180 254676 603208
rect 244976 603168 244982 603180
rect 254670 603168 254676 603180
rect 254728 603168 254734 603220
rect 181806 603100 181812 603152
rect 181864 603140 181870 603152
rect 214374 603140 214380 603152
rect 181864 603112 214380 603140
rect 181864 603100 181870 603112
rect 214374 603100 214380 603112
rect 214432 603100 214438 603152
rect 249702 603100 249708 603152
rect 249760 603140 249766 603152
rect 263594 603140 263600 603152
rect 249760 603112 263600 603140
rect 249760 603100 249766 603112
rect 263594 603100 263600 603112
rect 263652 603100 263658 603152
rect 180058 601740 180064 601792
rect 180116 601780 180122 601792
rect 229094 601780 229100 601792
rect 180116 601752 229100 601780
rect 180116 601740 180122 601752
rect 229094 601740 229100 601752
rect 229152 601740 229158 601792
rect 241054 601740 241060 601792
rect 241112 601780 241118 601792
rect 285674 601780 285680 601792
rect 241112 601752 285680 601780
rect 241112 601740 241118 601752
rect 285674 601740 285680 601752
rect 285732 601740 285738 601792
rect 104158 601672 104164 601724
rect 104216 601712 104222 601724
rect 211246 601712 211252 601724
rect 104216 601684 211252 601712
rect 104216 601672 104222 601684
rect 211246 601672 211252 601684
rect 211304 601672 211310 601724
rect 582742 601712 582748 601724
rect 213196 601684 582748 601712
rect 213196 601656 213224 601684
rect 582742 601672 582748 601684
rect 582800 601672 582806 601724
rect 211798 601604 211804 601656
rect 211856 601644 211862 601656
rect 213178 601644 213184 601656
rect 211856 601616 213184 601644
rect 211856 601604 211862 601616
rect 213178 601604 213184 601616
rect 213236 601604 213242 601656
rect 224218 601604 224224 601656
rect 224276 601644 224282 601656
rect 225230 601644 225236 601656
rect 224276 601616 225236 601644
rect 224276 601604 224282 601616
rect 225230 601604 225236 601616
rect 225288 601604 225294 601656
rect 221366 600788 221372 600840
rect 221424 600828 221430 600840
rect 226334 600828 226340 600840
rect 221424 600800 226340 600828
rect 221424 600788 221430 600800
rect 226334 600788 226340 600800
rect 226392 600788 226398 600840
rect 233878 600652 233884 600704
rect 233936 600692 233942 600704
rect 235350 600692 235356 600704
rect 233936 600664 235356 600692
rect 233936 600652 233942 600664
rect 235350 600652 235356 600664
rect 235408 600652 235414 600704
rect 141418 600380 141424 600432
rect 141476 600420 141482 600432
rect 200390 600420 200396 600432
rect 141476 600392 200396 600420
rect 141476 600380 141482 600392
rect 200390 600380 200396 600392
rect 200448 600380 200454 600432
rect 192478 600312 192484 600364
rect 192536 600352 192542 600364
rect 195422 600352 195428 600364
rect 192536 600324 195428 600352
rect 192536 600312 192542 600324
rect 195422 600312 195428 600324
rect 195480 600312 195486 600364
rect 212442 600312 212448 600364
rect 212500 600352 212506 600364
rect 219526 600352 219532 600364
rect 212500 600324 219532 600352
rect 212500 600312 212506 600324
rect 219526 600312 219532 600324
rect 219584 600312 219590 600364
rect 226334 600312 226340 600364
rect 226392 600352 226398 600364
rect 231762 600352 231768 600364
rect 226392 600324 231768 600352
rect 226392 600312 226398 600324
rect 231762 600312 231768 600324
rect 231820 600312 231826 600364
rect 232222 600312 232228 600364
rect 232280 600352 232286 600364
rect 248322 600352 248328 600364
rect 232280 600324 248328 600352
rect 232280 600312 232286 600324
rect 248322 600312 248328 600324
rect 248380 600312 248386 600364
rect 86954 599564 86960 599616
rect 87012 599604 87018 599616
rect 147674 599604 147680 599616
rect 87012 599576 147680 599604
rect 87012 599564 87018 599576
rect 147674 599564 147680 599576
rect 147732 599564 147738 599616
rect 222654 599428 222660 599480
rect 222712 599468 222718 599480
rect 223022 599468 223028 599480
rect 222712 599440 223028 599468
rect 222712 599428 222718 599440
rect 223022 599428 223028 599440
rect 223080 599428 223086 599480
rect 238726 599168 258074 599196
rect 193398 599088 193404 599140
rect 193456 599128 193462 599140
rect 193456 599100 200114 599128
rect 193456 599088 193462 599100
rect 184198 599020 184204 599072
rect 184256 599060 184262 599072
rect 197630 599060 197636 599072
rect 184256 599032 197636 599060
rect 184256 599020 184262 599032
rect 197630 599020 197636 599032
rect 197688 599020 197694 599072
rect 191190 598952 191196 599004
rect 191248 598992 191254 599004
rect 195606 598992 195612 599004
rect 191248 598964 195612 598992
rect 191248 598952 191254 598964
rect 195606 598952 195612 598964
rect 195664 598952 195670 599004
rect 200086 598992 200114 599100
rect 228634 599020 228640 599072
rect 228692 599060 228698 599072
rect 238726 599060 238754 599168
rect 228692 599032 238754 599060
rect 228692 599020 228698 599032
rect 251450 599020 251456 599072
rect 251508 599060 251514 599072
rect 253290 599060 253296 599072
rect 251508 599032 253296 599060
rect 251508 599020 251514 599032
rect 253290 599020 253296 599032
rect 253348 599020 253354 599072
rect 258046 599060 258074 599168
rect 271966 599060 271972 599072
rect 258046 599032 271972 599060
rect 271966 599020 271972 599032
rect 272024 599020 272030 599072
rect 214742 598992 214748 599004
rect 200086 598964 214748 598992
rect 214742 598952 214748 598964
rect 214800 598952 214806 599004
rect 222838 598952 222844 599004
rect 222896 598992 222902 599004
rect 276106 598992 276112 599004
rect 222896 598964 276112 598992
rect 222896 598952 222902 598964
rect 276106 598952 276112 598964
rect 276164 598952 276170 599004
rect 203334 598924 203340 598936
rect 200086 598896 203340 598924
rect 150158 597592 150164 597644
rect 150216 597632 150222 597644
rect 191006 597632 191012 597644
rect 150216 597604 191012 597632
rect 150216 597592 150222 597604
rect 191006 597592 191012 597604
rect 191064 597592 191070 597644
rect 84102 597524 84108 597576
rect 84160 597564 84166 597576
rect 133690 597564 133696 597576
rect 84160 597536 133696 597564
rect 84160 597524 84166 597536
rect 133690 597524 133696 597536
rect 133748 597524 133754 597576
rect 190362 597524 190368 597576
rect 190420 597564 190426 597576
rect 200086 597564 200114 598896
rect 203334 598884 203340 598896
rect 203392 598884 203398 598936
rect 247678 598884 247684 598936
rect 247736 598884 247742 598936
rect 249058 598884 249064 598936
rect 249116 598924 249122 598936
rect 253474 598924 253480 598936
rect 249116 598896 253480 598924
rect 249116 598884 249122 598896
rect 253474 598884 253480 598896
rect 253532 598884 253538 598936
rect 253906 598896 258074 598924
rect 247696 598856 247724 598884
rect 253906 598856 253934 598896
rect 247696 598828 253934 598856
rect 258046 598244 258074 598896
rect 295334 598244 295340 598256
rect 258046 598216 295340 598244
rect 295334 598204 295340 598216
rect 295392 598204 295398 598256
rect 190420 597536 200114 597564
rect 190420 597524 190426 597536
rect 253474 597524 253480 597576
rect 253532 597564 253538 597576
rect 273254 597564 273260 597576
rect 253532 597536 273260 597564
rect 253532 597524 253538 597536
rect 273254 597524 273260 597536
rect 273312 597524 273318 597576
rect 253382 596776 253388 596828
rect 253440 596816 253446 596828
rect 293954 596816 293960 596828
rect 253440 596788 293960 596816
rect 253440 596776 253446 596788
rect 293954 596776 293960 596788
rect 294012 596776 294018 596828
rect 146938 596232 146944 596284
rect 146996 596272 147002 596284
rect 191374 596272 191380 596284
rect 146996 596244 191380 596272
rect 146996 596232 147002 596244
rect 191374 596232 191380 596244
rect 191432 596232 191438 596284
rect 97258 596164 97264 596216
rect 97316 596204 97322 596216
rect 188246 596204 188252 596216
rect 97316 596176 188252 596204
rect 97316 596164 97322 596176
rect 188246 596164 188252 596176
rect 188304 596164 188310 596216
rect 166350 595416 166356 595468
rect 166408 595456 166414 595468
rect 192662 595456 192668 595468
rect 166408 595428 192668 595456
rect 166408 595416 166414 595428
rect 192662 595416 192668 595428
rect 192720 595416 192726 595468
rect 256602 595416 256608 595468
rect 256660 595456 256666 595468
rect 287054 595456 287060 595468
rect 256660 595428 287060 595456
rect 256660 595416 256666 595428
rect 287054 595416 287060 595428
rect 287112 595416 287118 595468
rect 92474 594804 92480 594856
rect 92532 594844 92538 594856
rect 166350 594844 166356 594856
rect 92532 594816 166356 594844
rect 92532 594804 92538 594816
rect 166350 594804 166356 594816
rect 166408 594844 166414 594856
rect 166626 594844 166632 594856
rect 166408 594816 166632 594844
rect 166408 594804 166414 594816
rect 166626 594804 166632 594816
rect 166684 594804 166690 594856
rect 69842 593376 69848 593428
rect 69900 593416 69906 593428
rect 142614 593416 142620 593428
rect 69900 593388 142620 593416
rect 69900 593376 69906 593388
rect 142614 593376 142620 593388
rect 142672 593376 142678 593428
rect 164878 593376 164884 593428
rect 164936 593416 164942 593428
rect 191282 593416 191288 593428
rect 164936 593388 191288 593416
rect 164936 593376 164942 593388
rect 191282 593376 191288 593388
rect 191340 593376 191346 593428
rect 255406 593376 255412 593428
rect 255464 593416 255470 593428
rect 261018 593416 261024 593428
rect 255464 593388 261024 593416
rect 255464 593376 255470 593388
rect 261018 593376 261024 593388
rect 261076 593416 261082 593428
rect 582650 593416 582656 593428
rect 261076 593388 582656 593416
rect 261076 593376 261082 593388
rect 582650 593376 582656 593388
rect 582708 593376 582714 593428
rect 89714 592628 89720 592680
rect 89772 592668 89778 592680
rect 192570 592668 192576 592680
rect 89772 592640 192576 592668
rect 89772 592628 89778 592640
rect 192570 592628 192576 592640
rect 192628 592628 192634 592680
rect 255406 592628 255412 592680
rect 255464 592668 255470 592680
rect 291194 592668 291200 592680
rect 255464 592640 291200 592668
rect 255464 592628 255470 592640
rect 291194 592628 291200 592640
rect 291252 592668 291258 592680
rect 299474 592668 299480 592680
rect 291252 592640 299480 592668
rect 291252 592628 291258 592640
rect 299474 592628 299480 592640
rect 299532 592628 299538 592680
rect 162118 592016 162124 592068
rect 162176 592056 162182 592068
rect 191374 592056 191380 592068
rect 162176 592028 191380 592056
rect 162176 592016 162182 592028
rect 191374 592016 191380 592028
rect 191432 592016 191438 592068
rect 71774 591268 71780 591320
rect 71832 591308 71838 591320
rect 184290 591308 184296 591320
rect 71832 591280 184296 591308
rect 71832 591268 71838 591280
rect 184290 591268 184296 591280
rect 184348 591268 184354 591320
rect 253382 591268 253388 591320
rect 253440 591308 253446 591320
rect 296714 591308 296720 591320
rect 253440 591280 296720 591308
rect 253440 591268 253446 591280
rect 296714 591268 296720 591280
rect 296772 591268 296778 591320
rect 157978 590656 157984 590708
rect 158036 590696 158042 590708
rect 191282 590696 191288 590708
rect 158036 590668 191288 590696
rect 158036 590656 158042 590668
rect 191282 590656 191288 590668
rect 191340 590656 191346 590708
rect 125502 589908 125508 589960
rect 125560 589948 125566 589960
rect 188430 589948 188436 589960
rect 125560 589920 188436 589948
rect 125560 589908 125566 589920
rect 188430 589908 188436 589920
rect 188488 589908 188494 589960
rect 91370 589296 91376 589348
rect 91428 589336 91434 589348
rect 124214 589336 124220 589348
rect 91428 589308 124220 589336
rect 91428 589296 91434 589308
rect 124214 589296 124220 589308
rect 124272 589336 124278 589348
rect 125502 589336 125508 589348
rect 124272 589308 125508 589336
rect 124272 589296 124278 589308
rect 125502 589296 125508 589308
rect 125560 589296 125566 589348
rect 179230 589296 179236 589348
rect 179288 589336 179294 589348
rect 191374 589336 191380 589348
rect 179288 589308 191380 589336
rect 179288 589296 179294 589308
rect 191374 589296 191380 589308
rect 191432 589296 191438 589348
rect 255406 589296 255412 589348
rect 255464 589336 255470 589348
rect 262398 589336 262404 589348
rect 255464 589308 262404 589336
rect 255464 589296 255470 589308
rect 262398 589296 262404 589308
rect 262456 589296 262462 589348
rect 78122 588616 78128 588668
rect 78180 588656 78186 588668
rect 88242 588656 88248 588668
rect 78180 588628 88248 588656
rect 78180 588616 78186 588628
rect 88242 588616 88248 588628
rect 88300 588656 88306 588668
rect 125594 588656 125600 588668
rect 88300 588628 125600 588656
rect 88300 588616 88306 588628
rect 125594 588616 125600 588628
rect 125652 588616 125658 588668
rect 40034 588548 40040 588600
rect 40092 588588 40098 588600
rect 95326 588588 95332 588600
rect 40092 588560 95332 588588
rect 40092 588548 40098 588560
rect 95326 588548 95332 588560
rect 95384 588548 95390 588600
rect 170398 588548 170404 588600
rect 170456 588588 170462 588600
rect 191650 588588 191656 588600
rect 170456 588560 191656 588588
rect 170456 588548 170462 588560
rect 191650 588548 191656 588560
rect 191708 588548 191714 588600
rect 254670 588548 254676 588600
rect 254728 588588 254734 588600
rect 274726 588588 274732 588600
rect 254728 588560 274732 588588
rect 254728 588548 254734 588560
rect 274726 588548 274732 588560
rect 274784 588548 274790 588600
rect 177942 587120 177948 587172
rect 178000 587160 178006 587172
rect 192478 587160 192484 587172
rect 178000 587132 192484 587160
rect 178000 587120 178006 587132
rect 192478 587120 192484 587132
rect 192536 587120 192542 587172
rect 176010 586508 176016 586560
rect 176068 586548 176074 586560
rect 190454 586548 190460 586560
rect 176068 586520 190460 586548
rect 176068 586508 176074 586520
rect 190454 586508 190460 586520
rect 190512 586508 190518 586560
rect 169662 585828 169668 585880
rect 169720 585868 169726 585880
rect 190546 585868 190552 585880
rect 169720 585840 190552 585868
rect 169720 585828 169726 585840
rect 190546 585828 190552 585840
rect 190604 585828 190610 585880
rect 147490 585760 147496 585812
rect 147548 585800 147554 585812
rect 191742 585800 191748 585812
rect 147548 585772 191748 585800
rect 147548 585760 147554 585772
rect 191742 585760 191748 585772
rect 191800 585760 191806 585812
rect 65978 585148 65984 585200
rect 66036 585188 66042 585200
rect 122190 585188 122196 585200
rect 66036 585160 122196 585188
rect 66036 585148 66042 585160
rect 122190 585148 122196 585160
rect 122248 585148 122254 585200
rect 260742 585148 260748 585200
rect 260800 585188 260806 585200
rect 266354 585188 266360 585200
rect 260800 585160 266360 585188
rect 260800 585148 260806 585160
rect 266354 585148 266360 585160
rect 266412 585148 266418 585200
rect 181438 584400 181444 584452
rect 181496 584440 181502 584452
rect 193398 584440 193404 584452
rect 181496 584412 193404 584440
rect 181496 584400 181502 584412
rect 193398 584400 193404 584412
rect 193456 584400 193462 584452
rect 255406 584400 255412 584452
rect 255464 584440 255470 584452
rect 259454 584440 259460 584452
rect 255464 584412 259460 584440
rect 255464 584400 255470 584412
rect 259454 584400 259460 584412
rect 259512 584440 259518 584452
rect 274818 584440 274824 584452
rect 259512 584412 274824 584440
rect 259512 584400 259518 584412
rect 274818 584400 274824 584412
rect 274876 584440 274882 584452
rect 582374 584440 582380 584452
rect 274876 584412 582380 584440
rect 274876 584400 274882 584412
rect 582374 584400 582380 584412
rect 582432 584400 582438 584452
rect 79962 583788 79968 583840
rect 80020 583828 80026 583840
rect 98546 583828 98552 583840
rect 80020 583800 98552 583828
rect 80020 583788 80026 583800
rect 98546 583788 98552 583800
rect 98604 583788 98610 583840
rect 74258 583720 74264 583772
rect 74316 583760 74322 583772
rect 122098 583760 122104 583772
rect 74316 583732 122104 583760
rect 74316 583720 74322 583732
rect 122098 583720 122104 583732
rect 122156 583720 122162 583772
rect 171778 583720 171784 583772
rect 171836 583760 171842 583772
rect 191742 583760 191748 583772
rect 171836 583732 191748 583760
rect 171836 583720 171842 583732
rect 191742 583720 191748 583732
rect 191800 583720 191806 583772
rect 255498 583720 255504 583772
rect 255556 583760 255562 583772
rect 266354 583760 266360 583772
rect 255556 583732 266360 583760
rect 255556 583720 255562 583732
rect 266354 583720 266360 583732
rect 266412 583720 266418 583772
rect 88242 583176 88248 583228
rect 88300 583216 88306 583228
rect 88978 583216 88984 583228
rect 88300 583188 88984 583216
rect 88300 583176 88306 583188
rect 88978 583176 88984 583188
rect 89036 583176 89042 583228
rect 259362 583040 259368 583092
rect 259420 583080 259426 583092
rect 268378 583080 268384 583092
rect 259420 583052 268384 583080
rect 259420 583040 259426 583052
rect 268378 583040 268384 583052
rect 268436 583040 268442 583092
rect 151722 582972 151728 583024
rect 151780 583012 151786 583024
rect 189718 583012 189724 583024
rect 151780 582984 189724 583012
rect 151780 582972 151786 582984
rect 189718 582972 189724 582984
rect 189776 582972 189782 583024
rect 254578 582972 254584 583024
rect 254636 583012 254642 583024
rect 283098 583012 283104 583024
rect 254636 582984 283104 583012
rect 254636 582972 254642 582984
rect 283098 582972 283104 582984
rect 283156 582972 283162 583024
rect 84102 582632 84108 582684
rect 84160 582672 84166 582684
rect 85022 582672 85028 582684
rect 84160 582644 85028 582672
rect 84160 582632 84166 582644
rect 85022 582632 85028 582644
rect 85080 582632 85086 582684
rect 55122 582428 55128 582480
rect 55180 582468 55186 582480
rect 82998 582468 83004 582480
rect 55180 582440 83004 582468
rect 55180 582428 55186 582440
rect 82998 582428 83004 582440
rect 83056 582428 83062 582480
rect 91002 582428 91008 582480
rect 91060 582468 91066 582480
rect 123478 582468 123484 582480
rect 91060 582440 123484 582468
rect 91060 582428 91066 582440
rect 123478 582428 123484 582440
rect 123536 582428 123542 582480
rect 67358 582360 67364 582412
rect 67416 582400 67422 582412
rect 71038 582400 71044 582412
rect 67416 582372 71044 582400
rect 67416 582360 67422 582372
rect 71038 582360 71044 582372
rect 71096 582360 71102 582412
rect 80698 582360 80704 582412
rect 80756 582400 80762 582412
rect 130470 582400 130476 582412
rect 80756 582372 130476 582400
rect 80756 582360 80762 582372
rect 130470 582360 130476 582372
rect 130528 582360 130534 582412
rect 255406 582360 255412 582412
rect 255464 582400 255470 582412
rect 258166 582400 258172 582412
rect 255464 582372 258172 582400
rect 255464 582360 255470 582372
rect 258166 582360 258172 582372
rect 258224 582400 258230 582412
rect 259362 582400 259368 582412
rect 258224 582372 259368 582400
rect 258224 582360 258230 582372
rect 259362 582360 259368 582372
rect 259420 582360 259426 582412
rect 76282 581068 76288 581120
rect 76340 581108 76346 581120
rect 108298 581108 108304 581120
rect 76340 581080 108304 581108
rect 76340 581068 76346 581080
rect 108298 581068 108304 581080
rect 108356 581068 108362 581120
rect 184842 581068 184848 581120
rect 184900 581108 184906 581120
rect 191190 581108 191196 581120
rect 184900 581080 191196 581108
rect 184900 581068 184906 581080
rect 191190 581068 191196 581080
rect 191248 581068 191254 581120
rect 80238 581040 80244 581052
rect 4172 581012 80244 581040
rect 3326 580932 3332 580984
rect 3384 580972 3390 580984
rect 4172 580972 4200 581012
rect 80238 581000 80244 581012
rect 80296 581000 80302 581052
rect 86586 581000 86592 581052
rect 86644 581040 86650 581052
rect 105538 581040 105544 581052
rect 86644 581012 105544 581040
rect 86644 581000 86650 581012
rect 105538 581000 105544 581012
rect 105596 581000 105602 581052
rect 173158 581000 173164 581052
rect 173216 581040 173222 581052
rect 191742 581040 191748 581052
rect 173216 581012 191748 581040
rect 173216 581000 173222 581012
rect 191742 581000 191748 581012
rect 191800 581000 191806 581052
rect 3384 580944 4200 580972
rect 3384 580932 3390 580944
rect 69014 580660 69020 580712
rect 69072 580660 69078 580712
rect 79042 580660 79048 580712
rect 79100 580700 79106 580712
rect 79100 580672 84194 580700
rect 79100 580660 79106 580672
rect 61930 579708 61936 579760
rect 61988 579748 61994 579760
rect 66898 579748 66904 579760
rect 61988 579720 66904 579748
rect 61988 579708 61994 579720
rect 66898 579708 66904 579720
rect 66956 579708 66962 579760
rect 53742 579640 53748 579692
rect 53800 579680 53806 579692
rect 69032 579680 69060 580660
rect 53800 579652 69060 579680
rect 84166 579680 84194 580672
rect 179046 580388 179052 580440
rect 179104 580428 179110 580440
rect 191006 580428 191012 580440
rect 179104 580400 191012 580428
rect 179104 580388 179110 580400
rect 191006 580388 191012 580400
rect 191064 580388 191070 580440
rect 159358 580252 159364 580304
rect 159416 580292 159422 580304
rect 179322 580292 179328 580304
rect 159416 580264 179328 580292
rect 159416 580252 159422 580264
rect 179322 580252 179328 580264
rect 179380 580292 179386 580304
rect 188430 580292 188436 580304
rect 179380 580264 188436 580292
rect 179380 580252 179386 580264
rect 188430 580252 188436 580264
rect 188488 580252 188494 580304
rect 255498 579708 255504 579760
rect 255556 579748 255562 579760
rect 262214 579748 262220 579760
rect 255556 579720 262220 579748
rect 255556 579708 255562 579720
rect 262214 579708 262220 579720
rect 262272 579708 262278 579760
rect 159358 579680 159364 579692
rect 84166 579652 159364 579680
rect 53800 579640 53806 579652
rect 159358 579640 159364 579652
rect 159416 579640 159422 579692
rect 255406 579640 255412 579692
rect 255464 579680 255470 579692
rect 288710 579680 288716 579692
rect 255464 579652 288716 579680
rect 255464 579640 255470 579652
rect 288710 579640 288716 579652
rect 288768 579640 288774 579692
rect 94958 579572 94964 579624
rect 95016 579612 95022 579624
rect 96706 579612 96712 579624
rect 95016 579584 96712 579612
rect 95016 579572 95022 579584
rect 96706 579572 96712 579584
rect 96764 579572 96770 579624
rect 188982 578280 188988 578332
rect 189040 578320 189046 578332
rect 190914 578320 190920 578332
rect 189040 578292 190920 578320
rect 189040 578280 189046 578292
rect 190914 578280 190920 578292
rect 190972 578280 190978 578332
rect 96890 578212 96896 578264
rect 96948 578252 96954 578264
rect 134518 578252 134524 578264
rect 96948 578224 134524 578252
rect 96948 578212 96954 578224
rect 134518 578212 134524 578224
rect 134576 578212 134582 578264
rect 148962 578212 148968 578264
rect 149020 578252 149026 578264
rect 191650 578252 191656 578264
rect 149020 578224 191656 578252
rect 149020 578212 149026 578224
rect 191650 578212 191656 578224
rect 191708 578212 191714 578264
rect 255314 578212 255320 578264
rect 255372 578252 255378 578264
rect 302234 578252 302240 578264
rect 255372 578224 302240 578252
rect 255372 578212 255378 578224
rect 302234 578212 302240 578224
rect 302292 578212 302298 578264
rect 98546 578144 98552 578196
rect 98604 578184 98610 578196
rect 191742 578184 191748 578196
rect 98604 578156 191748 578184
rect 98604 578144 98610 578156
rect 191742 578144 191748 578156
rect 191800 578144 191806 578196
rect 255406 577056 255412 577108
rect 255464 577096 255470 577108
rect 259546 577096 259552 577108
rect 255464 577068 259552 577096
rect 255464 577056 255470 577068
rect 259546 577056 259552 577068
rect 259604 577056 259610 577108
rect 255406 576852 255412 576904
rect 255464 576892 255470 576904
rect 267734 576892 267740 576904
rect 255464 576864 267740 576892
rect 255464 576852 255470 576864
rect 267734 576852 267740 576864
rect 267792 576852 267798 576904
rect 3418 576784 3424 576836
rect 3476 576824 3482 576836
rect 66162 576824 66168 576836
rect 3476 576796 66168 576824
rect 3476 576784 3482 576796
rect 66162 576784 66168 576796
rect 66220 576784 66226 576836
rect 97902 576784 97908 576836
rect 97960 576824 97966 576836
rect 160738 576824 160744 576836
rect 97960 576796 160744 576824
rect 97960 576784 97966 576796
rect 160738 576784 160744 576796
rect 160796 576784 160802 576836
rect 95878 576104 95884 576156
rect 95936 576144 95942 576156
rect 111058 576144 111064 576156
rect 95936 576116 111064 576144
rect 95936 576104 95942 576116
rect 111058 576104 111064 576116
rect 111116 576104 111122 576156
rect 186130 575560 186136 575612
rect 186188 575600 186194 575612
rect 191650 575600 191656 575612
rect 186188 575572 191656 575600
rect 186188 575560 186194 575572
rect 191650 575560 191656 575572
rect 191708 575560 191714 575612
rect 116578 575492 116584 575544
rect 116636 575532 116642 575544
rect 191742 575532 191748 575544
rect 116636 575504 191748 575532
rect 116636 575492 116642 575504
rect 191742 575492 191748 575504
rect 191800 575492 191806 575544
rect 255406 575492 255412 575544
rect 255464 575532 255470 575544
rect 278774 575532 278780 575544
rect 255464 575504 278780 575532
rect 255464 575492 255470 575504
rect 278774 575492 278780 575504
rect 278832 575492 278838 575544
rect 97902 574744 97908 574796
rect 97960 574784 97966 574796
rect 166442 574784 166448 574796
rect 97960 574756 166448 574784
rect 97960 574744 97966 574756
rect 166442 574744 166448 574756
rect 166500 574744 166506 574796
rect 168282 574744 168288 574796
rect 168340 574784 168346 574796
rect 191282 574784 191288 574796
rect 168340 574756 191288 574784
rect 168340 574744 168346 574756
rect 191282 574744 191288 574756
rect 191340 574744 191346 574796
rect 66070 574064 66076 574116
rect 66128 574104 66134 574116
rect 67358 574104 67364 574116
rect 66128 574076 67364 574104
rect 66128 574064 66134 574076
rect 67358 574064 67364 574076
rect 67416 574064 67422 574116
rect 157242 574064 157248 574116
rect 157300 574104 157306 574116
rect 190822 574104 190828 574116
rect 157300 574076 190828 574104
rect 157300 574064 157306 574076
rect 190822 574064 190828 574076
rect 190880 574064 190886 574116
rect 255406 574064 255412 574116
rect 255464 574104 255470 574116
rect 270494 574104 270500 574116
rect 255464 574076 270500 574104
rect 255464 574064 255470 574076
rect 270494 574064 270500 574076
rect 270552 574064 270558 574116
rect 97994 573316 98000 573368
rect 98052 573356 98058 573368
rect 137094 573356 137100 573368
rect 98052 573328 137100 573356
rect 98052 573316 98058 573328
rect 137094 573316 137100 573328
rect 137152 573316 137158 573368
rect 255958 573316 255964 573368
rect 256016 573356 256022 573368
rect 284294 573356 284300 573368
rect 256016 573328 284300 573356
rect 256016 573316 256022 573328
rect 284294 573316 284300 573328
rect 284352 573316 284358 573368
rect 97534 572976 97540 573028
rect 97592 573016 97598 573028
rect 100754 573016 100760 573028
rect 97592 572988 100760 573016
rect 97592 572976 97598 572988
rect 100754 572976 100760 572988
rect 100812 572976 100818 573028
rect 64782 572704 64788 572756
rect 64840 572744 64846 572756
rect 66806 572744 66812 572756
rect 64840 572716 66812 572744
rect 64840 572704 64846 572716
rect 66806 572704 66812 572716
rect 66864 572704 66870 572756
rect 136634 572704 136640 572756
rect 136692 572744 136698 572756
rect 137094 572744 137100 572756
rect 136692 572716 137100 572744
rect 136692 572704 136698 572716
rect 137094 572704 137100 572716
rect 137152 572744 137158 572756
rect 191742 572744 191748 572756
rect 137152 572716 191748 572744
rect 137152 572704 137158 572716
rect 191742 572704 191748 572716
rect 191800 572704 191806 572756
rect 188430 572636 188436 572688
rect 188488 572676 188494 572688
rect 190822 572676 190828 572688
rect 188488 572648 190828 572676
rect 188488 572636 188494 572648
rect 190822 572636 190828 572648
rect 190880 572636 190886 572688
rect 100754 571956 100760 572008
rect 100812 571996 100818 572008
rect 179414 571996 179420 572008
rect 100812 571968 179420 571996
rect 100812 571956 100818 571968
rect 179414 571956 179420 571968
rect 179472 571956 179478 572008
rect 255406 571412 255412 571464
rect 255464 571452 255470 571464
rect 277486 571452 277492 571464
rect 255464 571424 277492 571452
rect 255464 571412 255470 571424
rect 277486 571412 277492 571424
rect 277544 571412 277550 571464
rect 97718 571344 97724 571396
rect 97776 571384 97782 571396
rect 101398 571384 101404 571396
rect 97776 571356 101404 571384
rect 97776 571344 97782 571356
rect 101398 571344 101404 571356
rect 101456 571344 101462 571396
rect 255498 571344 255504 571396
rect 255556 571384 255562 571396
rect 286318 571384 286324 571396
rect 255556 571356 286324 571384
rect 255556 571344 255562 571356
rect 286318 571344 286324 571356
rect 286376 571344 286382 571396
rect 255406 571276 255412 571328
rect 255464 571316 255470 571328
rect 582558 571316 582564 571328
rect 255464 571288 582564 571316
rect 255464 571276 255470 571288
rect 582558 571276 582564 571288
rect 582616 571276 582622 571328
rect 105538 570596 105544 570648
rect 105596 570636 105602 570648
rect 160094 570636 160100 570648
rect 105596 570608 160100 570636
rect 105596 570596 105602 570608
rect 160094 570596 160100 570608
rect 160152 570596 160158 570648
rect 179414 570596 179420 570648
rect 179472 570636 179478 570648
rect 180518 570636 180524 570648
rect 179472 570608 180524 570636
rect 179472 570596 179478 570608
rect 180518 570596 180524 570608
rect 180576 570636 180582 570648
rect 191742 570636 191748 570648
rect 180576 570608 191748 570636
rect 180576 570596 180582 570608
rect 191742 570596 191748 570608
rect 191800 570596 191806 570648
rect 97902 569916 97908 569968
rect 97960 569956 97966 569968
rect 112530 569956 112536 569968
rect 97960 569928 112536 569956
rect 97960 569916 97966 569928
rect 112530 569916 112536 569928
rect 112588 569916 112594 569968
rect 160094 569916 160100 569968
rect 160152 569956 160158 569968
rect 191742 569956 191748 569968
rect 160152 569928 191748 569956
rect 160152 569916 160158 569928
rect 191742 569916 191748 569928
rect 191800 569916 191806 569968
rect 97902 569168 97908 569220
rect 97960 569208 97966 569220
rect 178678 569208 178684 569220
rect 97960 569180 178684 569208
rect 97960 569168 97966 569180
rect 178678 569168 178684 569180
rect 178736 569168 178742 569220
rect 255498 568624 255504 568676
rect 255556 568664 255562 568676
rect 267918 568664 267924 568676
rect 255556 568636 267924 568664
rect 255556 568624 255562 568636
rect 267918 568624 267924 568636
rect 267976 568624 267982 568676
rect 255406 568556 255412 568608
rect 255464 568596 255470 568608
rect 284386 568596 284392 568608
rect 255464 568568 284392 568596
rect 255464 568556 255470 568568
rect 284386 568556 284392 568568
rect 284444 568556 284450 568608
rect 130378 567808 130384 567860
rect 130436 567848 130442 567860
rect 178770 567848 178776 567860
rect 130436 567820 178776 567848
rect 130436 567808 130442 567820
rect 178770 567808 178776 567820
rect 178828 567808 178834 567860
rect 255682 567808 255688 567860
rect 255740 567848 255746 567860
rect 289814 567848 289820 567860
rect 255740 567820 289820 567848
rect 255740 567808 255746 567820
rect 289814 567808 289820 567820
rect 289872 567808 289878 567860
rect 59262 567196 59268 567248
rect 59320 567236 59326 567248
rect 66898 567236 66904 567248
rect 59320 567208 66904 567236
rect 59320 567196 59326 567208
rect 66898 567196 66904 567208
rect 66956 567196 66962 567248
rect 97902 567196 97908 567248
rect 97960 567236 97966 567248
rect 130378 567236 130384 567248
rect 97960 567208 130384 567236
rect 97960 567196 97966 567208
rect 130378 567196 130384 567208
rect 130436 567196 130442 567248
rect 187050 567196 187056 567248
rect 187108 567236 187114 567248
rect 191374 567236 191380 567248
rect 187108 567208 191380 567236
rect 187108 567196 187114 567208
rect 191374 567196 191380 567208
rect 191432 567196 191438 567248
rect 281994 566448 282000 566500
rect 282052 566488 282058 566500
rect 582466 566488 582472 566500
rect 282052 566460 582472 566488
rect 282052 566448 282058 566460
rect 582466 566448 582472 566460
rect 582524 566448 582530 566500
rect 255498 565904 255504 565956
rect 255556 565944 255562 565956
rect 281534 565944 281540 565956
rect 255556 565916 281540 565944
rect 255556 565904 255562 565916
rect 281534 565904 281540 565916
rect 281592 565944 281598 565956
rect 281994 565944 282000 565956
rect 281592 565916 282000 565944
rect 281592 565904 281598 565916
rect 281994 565904 282000 565916
rect 282052 565904 282058 565956
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 39298 565876 39304 565888
rect 3476 565848 39304 565876
rect 3476 565836 3482 565848
rect 39298 565836 39304 565848
rect 39356 565836 39362 565888
rect 52362 565836 52368 565888
rect 52420 565876 52426 565888
rect 67634 565876 67640 565888
rect 52420 565848 67640 565876
rect 52420 565836 52426 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 255590 565836 255596 565888
rect 255648 565876 255654 565888
rect 282914 565876 282920 565888
rect 255648 565848 282920 565876
rect 255648 565836 255654 565848
rect 282914 565836 282920 565848
rect 282972 565836 282978 565888
rect 169570 565156 169576 565208
rect 169628 565196 169634 565208
rect 187602 565196 187608 565208
rect 169628 565168 187608 565196
rect 169628 565156 169634 565168
rect 187602 565156 187608 565168
rect 187660 565196 187666 565208
rect 191742 565196 191748 565208
rect 187660 565168 191748 565196
rect 187660 565156 187666 565168
rect 191742 565156 191748 565168
rect 191800 565156 191806 565208
rect 150250 565088 150256 565140
rect 150308 565128 150314 565140
rect 186958 565128 186964 565140
rect 150308 565100 186964 565128
rect 150308 565088 150314 565100
rect 186958 565088 186964 565100
rect 187016 565088 187022 565140
rect 63402 564408 63408 564460
rect 63460 564448 63466 564460
rect 66438 564448 66444 564460
rect 63460 564420 66444 564448
rect 63460 564408 63466 564420
rect 66438 564408 66444 564420
rect 66496 564408 66502 564460
rect 187694 564408 187700 564460
rect 187752 564448 187758 564460
rect 191282 564448 191288 564460
rect 187752 564420 191288 564448
rect 187752 564408 187758 564420
rect 191282 564408 191288 564420
rect 191340 564408 191346 564460
rect 255498 564408 255504 564460
rect 255556 564448 255562 564460
rect 259454 564448 259460 564460
rect 255556 564420 259460 564448
rect 255556 564408 255562 564420
rect 259454 564408 259460 564420
rect 259512 564408 259518 564460
rect 122190 563660 122196 563712
rect 122248 563700 122254 563712
rect 122742 563700 122748 563712
rect 122248 563672 122748 563700
rect 122248 563660 122254 563672
rect 122742 563660 122748 563672
rect 122800 563700 122806 563712
rect 191742 563700 191748 563712
rect 122800 563672 191748 563700
rect 122800 563660 122806 563672
rect 191742 563660 191748 563672
rect 191800 563660 191806 563712
rect 97902 562300 97908 562352
rect 97960 562340 97966 562352
rect 106182 562340 106188 562352
rect 97960 562312 106188 562340
rect 97960 562300 97966 562312
rect 106182 562300 106188 562312
rect 106240 562340 106246 562352
rect 169018 562340 169024 562352
rect 106240 562312 169024 562340
rect 106240 562300 106246 562312
rect 169018 562300 169024 562312
rect 169076 562300 169082 562352
rect 177850 561688 177856 561740
rect 177908 561728 177914 561740
rect 190914 561728 190920 561740
rect 177908 561700 190920 561728
rect 177908 561688 177914 561700
rect 190914 561688 190920 561700
rect 190972 561688 190978 561740
rect 97902 560940 97908 560992
rect 97960 560980 97966 560992
rect 180058 560980 180064 560992
rect 97960 560952 180064 560980
rect 97960 560940 97966 560952
rect 180058 560940 180064 560952
rect 180116 560940 180122 560992
rect 64690 560328 64696 560380
rect 64748 560368 64754 560380
rect 66806 560368 66812 560380
rect 64748 560340 66812 560368
rect 64748 560328 64754 560340
rect 66806 560328 66812 560340
rect 66864 560328 66870 560380
rect 169478 560260 169484 560312
rect 169536 560300 169542 560312
rect 190822 560300 190828 560312
rect 169536 560272 190828 560300
rect 169536 560260 169542 560272
rect 190822 560260 190828 560272
rect 190880 560260 190886 560312
rect 255498 560260 255504 560312
rect 255556 560300 255562 560312
rect 266446 560300 266452 560312
rect 255556 560272 266452 560300
rect 255556 560260 255562 560272
rect 266446 560260 266452 560272
rect 266504 560260 266510 560312
rect 164050 559512 164056 559564
rect 164108 559552 164114 559564
rect 187694 559552 187700 559564
rect 164108 559524 187700 559552
rect 164108 559512 164114 559524
rect 187694 559512 187700 559524
rect 187752 559512 187758 559564
rect 255498 558968 255504 559020
rect 255556 559008 255562 559020
rect 269206 559008 269212 559020
rect 255556 558980 269212 559008
rect 255556 558968 255562 558980
rect 269206 558968 269212 558980
rect 269264 558968 269270 559020
rect 60642 558900 60648 558952
rect 60700 558940 60706 558952
rect 66806 558940 66812 558952
rect 60700 558912 66812 558940
rect 60700 558900 60706 558912
rect 66806 558900 66812 558912
rect 66864 558900 66870 558952
rect 96890 558900 96896 558952
rect 96948 558940 96954 558952
rect 113818 558940 113824 558952
rect 96948 558912 113824 558940
rect 96948 558900 96954 558912
rect 113818 558900 113824 558912
rect 113876 558900 113882 558952
rect 174538 558900 174544 558952
rect 174596 558940 174602 558952
rect 191742 558940 191748 558952
rect 174596 558912 191748 558940
rect 174596 558900 174602 558912
rect 191742 558900 191748 558912
rect 191800 558900 191806 558952
rect 255590 558900 255596 558952
rect 255648 558940 255654 558952
rect 273346 558940 273352 558952
rect 255648 558912 273352 558940
rect 255648 558900 255654 558912
rect 273346 558900 273352 558912
rect 273404 558900 273410 558952
rect 95142 558832 95148 558884
rect 95200 558872 95206 558884
rect 95326 558872 95332 558884
rect 95200 558844 95332 558872
rect 95200 558832 95206 558844
rect 95326 558832 95332 558844
rect 95384 558872 95390 558884
rect 184198 558872 184204 558884
rect 95384 558844 184204 558872
rect 95384 558832 95390 558844
rect 184198 558832 184204 558844
rect 184256 558832 184262 558884
rect 62022 557540 62028 557592
rect 62080 557580 62086 557592
rect 66806 557580 66812 557592
rect 62080 557552 66812 557580
rect 62080 557540 62086 557552
rect 66806 557540 66812 557552
rect 66864 557540 66870 557592
rect 159910 557540 159916 557592
rect 159968 557580 159974 557592
rect 191742 557580 191748 557592
rect 159968 557552 191748 557580
rect 159968 557540 159974 557552
rect 191742 557540 191748 557552
rect 191800 557540 191806 557592
rect 255590 557540 255596 557592
rect 255648 557580 255654 557592
rect 274634 557580 274640 557592
rect 255648 557552 274640 557580
rect 255648 557540 255654 557552
rect 274634 557540 274640 557552
rect 274692 557540 274698 557592
rect 97902 556792 97908 556844
rect 97960 556832 97966 556844
rect 115198 556832 115204 556844
rect 97960 556804 115204 556832
rect 97960 556792 97966 556804
rect 115198 556792 115204 556804
rect 115256 556792 115262 556844
rect 160830 556792 160836 556844
rect 160888 556832 160894 556844
rect 166350 556832 166356 556844
rect 160888 556804 166356 556832
rect 160888 556792 160894 556804
rect 166350 556792 166356 556804
rect 166408 556792 166414 556844
rect 166350 556180 166356 556232
rect 166408 556220 166414 556232
rect 191742 556220 191748 556232
rect 166408 556192 191748 556220
rect 166408 556180 166414 556192
rect 191742 556180 191748 556192
rect 191800 556180 191806 556232
rect 255590 556180 255596 556232
rect 255648 556220 255654 556232
rect 263686 556220 263692 556232
rect 255648 556192 263692 556220
rect 255648 556180 255654 556192
rect 263686 556180 263692 556192
rect 263744 556180 263750 556232
rect 173710 554820 173716 554872
rect 173768 554860 173774 554872
rect 191466 554860 191472 554872
rect 173768 554832 191472 554860
rect 173768 554820 173774 554832
rect 191466 554820 191472 554832
rect 191524 554820 191530 554872
rect 63310 554752 63316 554804
rect 63368 554792 63374 554804
rect 66530 554792 66536 554804
rect 63368 554764 66536 554792
rect 63368 554752 63374 554764
rect 66530 554752 66536 554764
rect 66588 554752 66594 554804
rect 162210 554752 162216 554804
rect 162268 554792 162274 554804
rect 180058 554792 180064 554804
rect 162268 554764 180064 554792
rect 162268 554752 162274 554764
rect 180058 554752 180064 554764
rect 180116 554752 180122 554804
rect 173250 554004 173256 554056
rect 173308 554044 173314 554056
rect 189718 554044 189724 554056
rect 173308 554016 189724 554044
rect 173308 554004 173314 554016
rect 189718 554004 189724 554016
rect 189776 554004 189782 554056
rect 3418 553664 3424 553716
rect 3476 553704 3482 553716
rect 7558 553704 7564 553716
rect 3476 553676 7564 553704
rect 3476 553664 3482 553676
rect 7558 553664 7564 553676
rect 7616 553664 7622 553716
rect 255590 553460 255596 553512
rect 255648 553500 255654 553512
rect 269482 553500 269488 553512
rect 255648 553472 269488 553500
rect 255648 553460 255654 553472
rect 269482 553460 269488 553472
rect 269540 553460 269546 553512
rect 56410 553392 56416 553444
rect 56468 553432 56474 553444
rect 66898 553432 66904 553444
rect 56468 553404 66904 553432
rect 56468 553392 56474 553404
rect 66898 553392 66904 553404
rect 66956 553392 66962 553444
rect 255682 553392 255688 553444
rect 255740 553432 255746 553444
rect 277578 553432 277584 553444
rect 255740 553404 277584 553432
rect 255740 553392 255746 553404
rect 277578 553392 277584 553404
rect 277636 553392 277642 553444
rect 255590 552644 255596 552696
rect 255648 552684 255654 552696
rect 260742 552684 260748 552696
rect 255648 552656 260748 552684
rect 255648 552644 255654 552656
rect 260742 552644 260748 552656
rect 260800 552684 260806 552696
rect 265066 552684 265072 552696
rect 260800 552656 265072 552684
rect 260800 552644 260806 552656
rect 265066 552644 265072 552656
rect 265124 552644 265130 552696
rect 180610 552100 180616 552152
rect 180668 552140 180674 552152
rect 191098 552140 191104 552152
rect 180668 552112 191104 552140
rect 180668 552100 180674 552112
rect 191098 552100 191104 552112
rect 191156 552100 191162 552152
rect 97902 552032 97908 552084
rect 97960 552072 97966 552084
rect 102042 552072 102048 552084
rect 97960 552044 102048 552072
rect 97960 552032 97966 552044
rect 102042 552032 102048 552044
rect 102100 552072 102106 552084
rect 184198 552072 184204 552084
rect 102100 552044 184204 552072
rect 102100 552032 102106 552044
rect 184198 552032 184204 552044
rect 184256 552032 184262 552084
rect 106182 551284 106188 551336
rect 106240 551324 106246 551336
rect 114738 551324 114744 551336
rect 106240 551296 114744 551324
rect 106240 551284 106246 551296
rect 114738 551284 114744 551296
rect 114796 551284 114802 551336
rect 122098 551284 122104 551336
rect 122156 551324 122162 551336
rect 160186 551324 160192 551336
rect 122156 551296 160192 551324
rect 122156 551284 122162 551296
rect 160186 551284 160192 551296
rect 160244 551284 160250 551336
rect 255590 550672 255596 550724
rect 255648 550712 255654 550724
rect 259638 550712 259644 550724
rect 255648 550684 259644 550712
rect 255648 550672 255654 550684
rect 259638 550672 259644 550684
rect 259696 550672 259702 550724
rect 160186 550604 160192 550656
rect 160244 550644 160250 550656
rect 160738 550644 160744 550656
rect 160244 550616 160744 550644
rect 160244 550604 160250 550616
rect 160738 550604 160744 550616
rect 160796 550644 160802 550656
rect 191742 550644 191748 550656
rect 160796 550616 191748 550644
rect 160796 550604 160802 550616
rect 191742 550604 191748 550616
rect 191800 550604 191806 550656
rect 97810 549856 97816 549908
rect 97868 549896 97874 549908
rect 162302 549896 162308 549908
rect 97868 549868 162308 549896
rect 97868 549856 97874 549868
rect 162302 549856 162308 549868
rect 162360 549856 162366 549908
rect 255590 549856 255596 549908
rect 255648 549896 255654 549908
rect 258074 549896 258080 549908
rect 255648 549868 258080 549896
rect 255648 549856 255654 549868
rect 258074 549856 258080 549868
rect 258132 549896 258138 549908
rect 269114 549896 269120 549908
rect 258132 549868 269120 549896
rect 258132 549856 258138 549868
rect 269114 549856 269120 549868
rect 269172 549856 269178 549908
rect 186038 549312 186044 549364
rect 186096 549352 186102 549364
rect 191742 549352 191748 549364
rect 186096 549324 191748 549352
rect 186096 549312 186102 549324
rect 191742 549312 191748 549324
rect 191800 549312 191806 549364
rect 162302 549244 162308 549296
rect 162360 549284 162366 549296
rect 188522 549284 188528 549296
rect 162360 549256 188528 549284
rect 162360 549244 162366 549256
rect 188522 549244 188528 549256
rect 188580 549244 188586 549296
rect 102042 548496 102048 548548
rect 102100 548536 102106 548548
rect 112438 548536 112444 548548
rect 102100 548508 112444 548536
rect 102100 548496 102106 548508
rect 112438 548496 112444 548508
rect 112496 548496 112502 548548
rect 112530 548496 112536 548548
rect 112588 548536 112594 548548
rect 188430 548536 188436 548548
rect 112588 548508 188436 548536
rect 112588 548496 112594 548508
rect 188430 548496 188436 548508
rect 188488 548496 188494 548548
rect 187510 547884 187516 547936
rect 187568 547924 187574 547936
rect 190638 547924 190644 547936
rect 187568 547896 190644 547924
rect 187568 547884 187574 547896
rect 190638 547884 190644 547896
rect 190696 547884 190702 547936
rect 255590 547884 255596 547936
rect 255648 547924 255654 547936
rect 262306 547924 262312 547936
rect 255648 547896 262312 547924
rect 255648 547884 255654 547896
rect 262306 547884 262312 547896
rect 262364 547884 262370 547936
rect 156598 546524 156604 546576
rect 156656 546564 156662 546576
rect 191650 546564 191656 546576
rect 156656 546536 191656 546564
rect 156656 546524 156662 546536
rect 191650 546524 191656 546536
rect 191708 546524 191714 546576
rect 99374 546456 99380 546508
rect 99432 546496 99438 546508
rect 191558 546496 191564 546508
rect 99432 546468 191564 546496
rect 99432 546456 99438 546468
rect 191558 546456 191564 546468
rect 191616 546456 191622 546508
rect 255498 546456 255504 546508
rect 255556 546496 255562 546508
rect 276198 546496 276204 546508
rect 255556 546468 276204 546496
rect 255556 546456 255562 546468
rect 276198 546456 276204 546468
rect 276256 546456 276262 546508
rect 106918 545708 106924 545760
rect 106976 545748 106982 545760
rect 186958 545748 186964 545760
rect 106976 545720 186964 545748
rect 106976 545708 106982 545720
rect 186958 545708 186964 545720
rect 187016 545708 187022 545760
rect 97074 545232 97080 545284
rect 97132 545272 97138 545284
rect 100018 545272 100024 545284
rect 97132 545244 100024 545272
rect 97132 545232 97138 545244
rect 100018 545232 100024 545244
rect 100076 545232 100082 545284
rect 255498 545232 255504 545284
rect 255556 545272 255562 545284
rect 258350 545272 258356 545284
rect 255556 545244 258356 545272
rect 255556 545232 255562 545244
rect 258350 545232 258356 545244
rect 258408 545232 258414 545284
rect 168190 545096 168196 545148
rect 168248 545136 168254 545148
rect 191650 545136 191656 545148
rect 168248 545108 191656 545136
rect 168248 545096 168254 545108
rect 191650 545096 191656 545108
rect 191708 545096 191714 545148
rect 180058 545028 180064 545080
rect 180116 545068 180122 545080
rect 191558 545068 191564 545080
rect 180116 545040 191564 545068
rect 180116 545028 180122 545040
rect 191558 545028 191564 545040
rect 191616 545028 191622 545080
rect 50982 543736 50988 543788
rect 51040 543776 51046 543788
rect 66806 543776 66812 543788
rect 51040 543748 66812 543776
rect 51040 543736 51046 543748
rect 66806 543736 66812 543748
rect 66864 543736 66870 543788
rect 97534 543736 97540 543788
rect 97592 543776 97598 543788
rect 104250 543776 104256 543788
rect 97592 543748 104256 543776
rect 97592 543736 97598 543748
rect 104250 543736 104256 543748
rect 104308 543736 104314 543788
rect 184750 543736 184756 543788
rect 184808 543776 184814 543788
rect 191006 543776 191012 543788
rect 184808 543748 191012 543776
rect 184808 543736 184814 543748
rect 191006 543736 191012 543748
rect 191064 543736 191070 543788
rect 33778 543668 33784 543720
rect 33836 543708 33842 543720
rect 66254 543708 66260 543720
rect 33836 543680 66260 543708
rect 33836 543668 33842 543680
rect 66254 543668 66260 543680
rect 66312 543668 66318 543720
rect 166442 542988 166448 543040
rect 166500 543028 166506 543040
rect 181530 543028 181536 543040
rect 166500 543000 181536 543028
rect 166500 542988 166506 543000
rect 181530 542988 181536 543000
rect 181588 542988 181594 543040
rect 255590 542444 255596 542496
rect 255648 542484 255654 542496
rect 264974 542484 264980 542496
rect 255648 542456 264980 542484
rect 255648 542444 255654 542456
rect 264974 542444 264980 542456
rect 265032 542444 265038 542496
rect 97534 542376 97540 542428
rect 97592 542416 97598 542428
rect 158806 542416 158812 542428
rect 97592 542388 158812 542416
rect 97592 542376 97598 542388
rect 158806 542376 158812 542388
rect 158864 542416 158870 542428
rect 186314 542416 186320 542428
rect 158864 542388 186320 542416
rect 158864 542376 158870 542388
rect 186314 542376 186320 542388
rect 186372 542376 186378 542428
rect 255498 542376 255504 542428
rect 255556 542416 255562 542428
rect 267826 542416 267832 542428
rect 255556 542388 267832 542416
rect 255556 542376 255562 542388
rect 267826 542376 267832 542388
rect 267884 542376 267890 542428
rect 184658 542308 184664 542360
rect 184716 542348 184722 542360
rect 187050 542348 187056 542360
rect 184716 542320 187056 542348
rect 184716 542308 184722 542320
rect 187050 542308 187056 542320
rect 187108 542308 187114 542360
rect 123478 541696 123484 541748
rect 123536 541736 123542 541748
rect 155770 541736 155776 541748
rect 123536 541708 155776 541736
rect 123536 541696 123542 541708
rect 155770 541696 155776 541708
rect 155828 541696 155834 541748
rect 15838 541628 15844 541680
rect 15896 541668 15902 541680
rect 39942 541668 39948 541680
rect 15896 541640 39948 541668
rect 15896 541628 15902 541640
rect 39942 541628 39948 541640
rect 40000 541628 40006 541680
rect 97902 541628 97908 541680
rect 97960 541668 97966 541680
rect 146938 541668 146944 541680
rect 97960 541640 146944 541668
rect 97960 541628 97966 541640
rect 146938 541628 146944 541640
rect 146996 541628 147002 541680
rect 178402 541628 178408 541680
rect 178460 541668 178466 541680
rect 179138 541668 179144 541680
rect 178460 541640 179144 541668
rect 178460 541628 178466 541640
rect 179138 541628 179144 541640
rect 179196 541668 179202 541680
rect 188338 541668 188344 541680
rect 179196 541640 188344 541668
rect 179196 541628 179202 541640
rect 188338 541628 188344 541640
rect 188396 541628 188402 541680
rect 278038 541628 278044 541680
rect 278096 541668 278102 541680
rect 287146 541668 287152 541680
rect 278096 541640 287152 541668
rect 278096 541628 278102 541640
rect 287146 541628 287152 541640
rect 287204 541628 287210 541680
rect 39942 540948 39948 541000
rect 40000 540988 40006 541000
rect 66254 540988 66260 541000
rect 40000 540960 66260 540988
rect 40000 540948 40006 540960
rect 66254 540948 66260 540960
rect 66312 540948 66318 541000
rect 155770 540948 155776 541000
rect 155828 540988 155834 541000
rect 178402 540988 178408 541000
rect 155828 540960 178408 540988
rect 155828 540948 155834 540960
rect 178402 540948 178408 540960
rect 178460 540948 178466 541000
rect 188522 540540 188528 540592
rect 188580 540580 188586 540592
rect 191650 540580 191656 540592
rect 188580 540552 191656 540580
rect 188580 540540 188586 540552
rect 191650 540540 191656 540552
rect 191708 540540 191714 540592
rect 177390 540200 177396 540252
rect 177448 540240 177454 540252
rect 184750 540240 184756 540252
rect 177448 540212 184756 540240
rect 177448 540200 177454 540212
rect 184750 540200 184756 540212
rect 184808 540200 184814 540252
rect 67818 539792 67824 539844
rect 67876 539832 67882 539844
rect 71774 539832 71780 539844
rect 67876 539804 71780 539832
rect 67876 539792 67882 539804
rect 71774 539792 71780 539804
rect 71832 539792 71838 539844
rect 94130 539656 94136 539708
rect 94188 539696 94194 539708
rect 94774 539696 94780 539708
rect 94188 539668 94780 539696
rect 94188 539656 94194 539668
rect 94774 539656 94780 539668
rect 94832 539656 94838 539708
rect 259546 539696 259552 539708
rect 251468 539668 259552 539696
rect 57790 539588 57796 539640
rect 57848 539628 57854 539640
rect 66254 539628 66260 539640
rect 57848 539600 66260 539628
rect 57848 539588 57854 539600
rect 66254 539588 66260 539600
rect 66312 539588 66318 539640
rect 88150 539588 88156 539640
rect 88208 539628 88214 539640
rect 134610 539628 134616 539640
rect 88208 539600 134616 539628
rect 88208 539588 88214 539600
rect 134610 539588 134616 539600
rect 134668 539628 134674 539640
rect 164326 539628 164332 539640
rect 134668 539600 164332 539628
rect 134668 539588 134674 539600
rect 164326 539588 164332 539600
rect 164384 539588 164390 539640
rect 251468 539368 251496 539668
rect 259546 539656 259552 539668
rect 259604 539656 259610 539708
rect 255498 539588 255504 539640
rect 255556 539628 255562 539640
rect 278866 539628 278872 539640
rect 255556 539600 278872 539628
rect 255556 539588 255562 539600
rect 278866 539588 278872 539600
rect 278924 539588 278930 539640
rect 251450 539316 251456 539368
rect 251508 539316 251514 539368
rect 250438 539248 250444 539300
rect 250496 539288 250502 539300
rect 255774 539288 255780 539300
rect 250496 539260 255780 539288
rect 250496 539248 250502 539260
rect 255774 539248 255780 539260
rect 255832 539248 255838 539300
rect 67634 538840 67640 538892
rect 67692 538880 67698 538892
rect 83458 538880 83464 538892
rect 67692 538852 83464 538880
rect 67692 538840 67698 538852
rect 83458 538840 83464 538852
rect 83516 538840 83522 538892
rect 119338 538840 119344 538892
rect 119396 538880 119402 538892
rect 150434 538880 150440 538892
rect 119396 538852 150440 538880
rect 119396 538840 119402 538852
rect 150434 538840 150440 538852
rect 150492 538840 150498 538892
rect 43438 538296 43444 538348
rect 43496 538336 43502 538348
rect 94590 538336 94596 538348
rect 43496 538308 94596 538336
rect 43496 538296 43502 538308
rect 94590 538296 94596 538308
rect 94648 538336 94654 538348
rect 104158 538336 104164 538348
rect 94648 538308 104164 538336
rect 94648 538296 94654 538308
rect 104158 538296 104164 538308
rect 104216 538296 104222 538348
rect 186314 538296 186320 538348
rect 186372 538336 186378 538348
rect 221366 538336 221372 538348
rect 186372 538308 221372 538336
rect 186372 538296 186378 538308
rect 221366 538296 221372 538308
rect 221424 538296 221430 538348
rect 255498 538296 255504 538348
rect 255556 538336 255562 538348
rect 277394 538336 277400 538348
rect 255556 538308 277400 538336
rect 255556 538296 255562 538308
rect 277394 538296 277400 538308
rect 277452 538296 277458 538348
rect 85574 538228 85580 538280
rect 85632 538268 85638 538280
rect 85758 538268 85764 538280
rect 85632 538240 85764 538268
rect 85632 538228 85638 538240
rect 85758 538228 85764 538240
rect 85816 538268 85822 538280
rect 99374 538268 99380 538280
rect 85816 538240 99380 538268
rect 85816 538228 85822 538240
rect 99374 538228 99380 538240
rect 99432 538228 99438 538280
rect 150434 538228 150440 538280
rect 150492 538268 150498 538280
rect 151630 538268 151636 538280
rect 150492 538240 151636 538268
rect 150492 538228 150498 538240
rect 151630 538228 151636 538240
rect 151688 538268 151694 538280
rect 216398 538268 216404 538280
rect 151688 538240 216404 538268
rect 151688 538228 151694 538240
rect 216398 538228 216404 538240
rect 216456 538228 216462 538280
rect 224678 538228 224684 538280
rect 224736 538268 224742 538280
rect 582926 538268 582932 538280
rect 224736 538240 582932 538268
rect 224736 538228 224742 538240
rect 582926 538228 582932 538240
rect 582984 538228 582990 538280
rect 7558 538160 7564 538212
rect 7616 538200 7622 538212
rect 70670 538200 70676 538212
rect 7616 538172 70676 538200
rect 7616 538160 7622 538172
rect 70670 538160 70676 538172
rect 70728 538160 70734 538212
rect 79962 538160 79968 538212
rect 80020 538200 80026 538212
rect 116578 538200 116584 538212
rect 80020 538172 116584 538200
rect 80020 538160 80026 538172
rect 116578 538160 116584 538172
rect 116636 538160 116642 538212
rect 184198 538160 184204 538212
rect 184256 538200 184262 538212
rect 200390 538200 200396 538212
rect 184256 538172 200396 538200
rect 184256 538160 184262 538172
rect 200390 538160 200396 538172
rect 200448 538160 200454 538212
rect 239214 538160 239220 538212
rect 239272 538200 239278 538212
rect 239398 538200 239404 538212
rect 239272 538172 239404 538200
rect 239272 538160 239278 538172
rect 239398 538160 239404 538172
rect 239456 538200 239462 538212
rect 582374 538200 582380 538212
rect 239456 538172 582380 538200
rect 239456 538160 239462 538172
rect 582374 538160 582380 538172
rect 582432 538160 582438 538212
rect 178678 538092 178684 538144
rect 178736 538132 178742 538144
rect 244366 538132 244372 538144
rect 178736 538104 244372 538132
rect 178736 538092 178742 538104
rect 244366 538092 244372 538104
rect 244424 538092 244430 538144
rect 79226 537684 79232 537736
rect 79284 537724 79290 537736
rect 79962 537724 79968 537736
rect 79284 537696 79968 537724
rect 79284 537684 79290 537696
rect 79962 537684 79968 537696
rect 80020 537684 80026 537736
rect 66070 537480 66076 537532
rect 66128 537520 66134 537532
rect 143626 537520 143632 537532
rect 66128 537492 143632 537520
rect 66128 537480 66134 537492
rect 143626 537480 143632 537492
rect 143684 537480 143690 537532
rect 70670 536800 70676 536852
rect 70728 536840 70734 536852
rect 71038 536840 71044 536852
rect 70728 536812 71044 536840
rect 70728 536800 70734 536812
rect 71038 536800 71044 536812
rect 71096 536800 71102 536852
rect 57238 536732 57244 536784
rect 57296 536772 57302 536784
rect 73246 536772 73252 536784
rect 57296 536744 73252 536772
rect 57296 536732 57302 536744
rect 73246 536732 73252 536744
rect 73304 536732 73310 536784
rect 87690 536732 87696 536784
rect 87748 536772 87754 536784
rect 215294 536772 215300 536784
rect 87748 536744 215300 536772
rect 87748 536732 87754 536744
rect 215294 536732 215300 536744
rect 215352 536732 215358 536784
rect 82170 536664 82176 536716
rect 82228 536704 82234 536716
rect 88150 536704 88156 536716
rect 82228 536676 88156 536704
rect 82228 536664 82234 536676
rect 88150 536664 88156 536676
rect 88208 536664 88214 536716
rect 211982 536664 211988 536716
rect 212040 536704 212046 536716
rect 280798 536704 280804 536716
rect 212040 536676 280804 536704
rect 212040 536664 212046 536676
rect 280798 536664 280804 536676
rect 280856 536664 280862 536716
rect 39298 536052 39304 536104
rect 39356 536092 39362 536104
rect 53650 536092 53656 536104
rect 39356 536064 53656 536092
rect 39356 536052 39362 536064
rect 53650 536052 53656 536064
rect 53708 536092 53714 536104
rect 69382 536092 69388 536104
rect 53708 536064 69388 536092
rect 53708 536052 53714 536064
rect 69382 536052 69388 536064
rect 69440 536052 69446 536104
rect 73246 536052 73252 536104
rect 73304 536092 73310 536104
rect 81434 536092 81440 536104
rect 73304 536064 81440 536092
rect 73304 536052 73310 536064
rect 81434 536052 81440 536064
rect 81492 536052 81498 536104
rect 188338 536052 188344 536104
rect 188396 536092 188402 536104
rect 205542 536092 205548 536104
rect 188396 536064 205548 536092
rect 188396 536052 188402 536064
rect 205542 536052 205548 536064
rect 205600 536052 205606 536104
rect 253198 536052 253204 536104
rect 253256 536092 253262 536104
rect 260834 536092 260840 536104
rect 253256 536064 260840 536092
rect 253256 536052 253262 536064
rect 260834 536052 260840 536064
rect 260892 536052 260898 536104
rect 225230 535984 225236 536036
rect 225288 536024 225294 536036
rect 226978 536024 226984 536036
rect 225288 535996 226984 536024
rect 225288 535984 225294 535996
rect 226978 535984 226984 535996
rect 227036 535984 227042 536036
rect 233418 535780 233424 535832
rect 233476 535820 233482 535832
rect 236638 535820 236644 535832
rect 233476 535792 236644 535820
rect 233476 535780 233482 535792
rect 236638 535780 236644 535792
rect 236696 535780 236702 535832
rect 220078 535508 220084 535560
rect 220136 535548 220142 535560
rect 223390 535548 223396 535560
rect 220136 535520 223396 535548
rect 220136 535508 220142 535520
rect 223390 535508 223396 535520
rect 223448 535508 223454 535560
rect 86218 535440 86224 535492
rect 86276 535480 86282 535492
rect 89806 535480 89812 535492
rect 86276 535452 89812 535480
rect 86276 535440 86282 535452
rect 89806 535440 89812 535452
rect 89864 535440 89870 535492
rect 91002 535440 91008 535492
rect 91060 535480 91066 535492
rect 91830 535480 91836 535492
rect 91060 535452 91836 535480
rect 91060 535440 91066 535452
rect 91830 535440 91836 535452
rect 91888 535440 91894 535492
rect 206370 535440 206376 535492
rect 206428 535480 206434 535492
rect 209958 535480 209964 535492
rect 206428 535452 209964 535480
rect 206428 535440 206434 535452
rect 209958 535440 209964 535452
rect 210016 535440 210022 535492
rect 215938 535440 215944 535492
rect 215996 535480 216002 535492
rect 218974 535480 218980 535492
rect 215996 535452 218980 535480
rect 215996 535440 216002 535452
rect 218974 535440 218980 535452
rect 219032 535440 219038 535492
rect 222838 535440 222844 535492
rect 222896 535480 222902 535492
rect 223942 535480 223948 535492
rect 222896 535452 223948 535480
rect 222896 535440 222902 535452
rect 223942 535440 223948 535452
rect 224000 535440 224006 535492
rect 229646 535440 229652 535492
rect 229704 535480 229710 535492
rect 233878 535480 233884 535492
rect 229704 535452 233884 535480
rect 229704 535440 229710 535452
rect 233878 535440 233884 535452
rect 233936 535440 233942 535492
rect 242986 535440 242992 535492
rect 243044 535480 243050 535492
rect 250622 535480 250628 535492
rect 243044 535452 250628 535480
rect 243044 535440 243050 535452
rect 250622 535440 250628 535452
rect 250680 535440 250686 535492
rect 88242 535372 88248 535424
rect 88300 535412 88306 535424
rect 95418 535412 95424 535424
rect 88300 535384 95424 535412
rect 88300 535372 88306 535384
rect 95418 535372 95424 535384
rect 95476 535372 95482 535424
rect 186958 535372 186964 535424
rect 187016 535412 187022 535424
rect 238202 535412 238208 535424
rect 187016 535384 238208 535412
rect 187016 535372 187022 535384
rect 238202 535372 238208 535384
rect 238260 535412 238266 535424
rect 238662 535412 238668 535424
rect 238260 535384 238668 535412
rect 238260 535372 238266 535384
rect 238662 535372 238668 535384
rect 238720 535372 238726 535424
rect 164326 535304 164332 535356
rect 164384 535344 164390 535356
rect 197998 535344 198004 535356
rect 164384 535316 198004 535344
rect 164384 535304 164390 535316
rect 197998 535304 198004 535316
rect 198056 535304 198062 535356
rect 249058 534760 249064 534812
rect 249116 534800 249122 534812
rect 258166 534800 258172 534812
rect 249116 534772 258172 534800
rect 249116 534760 249122 534772
rect 258166 534760 258172 534772
rect 258224 534760 258230 534812
rect 82722 534692 82728 534744
rect 82780 534732 82786 534744
rect 94682 534732 94688 534744
rect 82780 534704 94688 534732
rect 82780 534692 82786 534704
rect 94682 534692 94688 534704
rect 94740 534692 94746 534744
rect 216030 534692 216036 534744
rect 216088 534732 216094 534744
rect 230382 534732 230388 534744
rect 216088 534704 230388 534732
rect 216088 534692 216094 534704
rect 230382 534692 230388 534704
rect 230440 534692 230446 534744
rect 246390 534692 246396 534744
rect 246448 534732 246454 534744
rect 256878 534732 256884 534744
rect 246448 534704 256884 534732
rect 246448 534692 246454 534704
rect 256878 534692 256884 534704
rect 256936 534692 256942 534744
rect 211982 534420 211988 534472
rect 212040 534460 212046 534472
rect 212718 534460 212724 534472
rect 212040 534432 212724 534460
rect 212040 534420 212046 534432
rect 212718 534420 212724 534432
rect 212776 534420 212782 534472
rect 130470 534012 130476 534064
rect 130528 534052 130534 534064
rect 130930 534052 130936 534064
rect 130528 534024 130936 534052
rect 130528 534012 130534 534024
rect 130930 534012 130936 534024
rect 130988 534052 130994 534064
rect 242986 534052 242992 534064
rect 130988 534024 242992 534052
rect 130988 534012 130994 534024
rect 242986 534012 242992 534024
rect 243044 534012 243050 534064
rect 81434 533400 81440 533452
rect 81492 533440 81498 533452
rect 102778 533440 102784 533452
rect 81492 533412 102784 533440
rect 81492 533400 81498 533412
rect 102778 533400 102784 533412
rect 102836 533400 102842 533452
rect 195974 533400 195980 533452
rect 196032 533440 196038 533452
rect 198826 533440 198832 533452
rect 196032 533412 198832 533440
rect 196032 533400 196038 533412
rect 198826 533400 198832 533412
rect 198884 533400 198890 533452
rect 233418 533440 233424 533452
rect 219406 533412 233424 533440
rect 59170 533332 59176 533384
rect 59228 533372 59234 533384
rect 73154 533372 73160 533384
rect 59228 533344 73160 533372
rect 59228 533332 59234 533344
rect 73154 533332 73160 533344
rect 73212 533332 73218 533384
rect 75822 533332 75828 533384
rect 75880 533372 75886 533384
rect 96798 533372 96804 533384
rect 75880 533344 96804 533372
rect 75880 533332 75886 533344
rect 96798 533332 96804 533344
rect 96856 533332 96862 533384
rect 212534 533332 212540 533384
rect 212592 533372 212598 533384
rect 213454 533372 213460 533384
rect 212592 533344 213460 533372
rect 212592 533332 212598 533344
rect 213454 533332 213460 533344
rect 213512 533332 213518 533384
rect 216674 533332 216680 533384
rect 216732 533372 216738 533384
rect 217318 533372 217324 533384
rect 216732 533344 217324 533372
rect 216732 533332 216738 533344
rect 217318 533332 217324 533344
rect 217376 533332 217382 533384
rect 213178 533196 213184 533248
rect 213236 533236 213242 533248
rect 219406 533236 219434 533412
rect 233418 533400 233424 533412
rect 233476 533400 233482 533452
rect 246942 533400 246948 533452
rect 247000 533440 247006 533452
rect 255866 533440 255872 533452
rect 247000 533412 255872 533440
rect 247000 533400 247006 533412
rect 255866 533400 255872 533412
rect 255924 533400 255930 533452
rect 233234 533332 233240 533384
rect 233292 533372 233298 533384
rect 233694 533372 233700 533384
rect 233292 533344 233700 533372
rect 233292 533332 233298 533344
rect 233694 533332 233700 533344
rect 233752 533332 233758 533384
rect 234614 533332 234620 533384
rect 234672 533372 234678 533384
rect 234982 533372 234988 533384
rect 234672 533344 234988 533372
rect 234672 533332 234678 533344
rect 234982 533332 234988 533344
rect 235040 533332 235046 533384
rect 237374 533332 237380 533384
rect 237432 533372 237438 533384
rect 237558 533372 237564 533384
rect 237432 533344 237564 533372
rect 237432 533332 237438 533344
rect 237558 533332 237564 533344
rect 237616 533332 237622 533384
rect 240134 533332 240140 533384
rect 240192 533372 240198 533384
rect 240686 533372 240692 533384
rect 240192 533344 240692 533372
rect 240192 533332 240198 533344
rect 240686 533332 240692 533344
rect 240744 533332 240750 533384
rect 247034 533332 247040 533384
rect 247092 533372 247098 533384
rect 247678 533372 247684 533384
rect 247092 533344 247684 533372
rect 247092 533332 247098 533344
rect 247678 533332 247684 533344
rect 247736 533332 247742 533384
rect 251910 533332 251916 533384
rect 251968 533372 251974 533384
rect 280338 533372 280344 533384
rect 251968 533344 280344 533372
rect 251968 533332 251974 533344
rect 280338 533332 280344 533344
rect 280396 533332 280402 533384
rect 213236 533208 219434 533236
rect 213236 533196 213242 533208
rect 201494 532720 201500 532772
rect 201552 532760 201558 532772
rect 202046 532760 202052 532772
rect 201552 532732 202052 532760
rect 201552 532720 201558 532732
rect 202046 532720 202052 532732
rect 202104 532720 202110 532772
rect 231854 532720 231860 532772
rect 231912 532760 231918 532772
rect 232406 532760 232412 532772
rect 231912 532732 232412 532760
rect 231912 532720 231918 532732
rect 232406 532720 232412 532732
rect 232464 532720 232470 532772
rect 179138 532652 179144 532704
rect 179196 532692 179202 532704
rect 206830 532692 206836 532704
rect 179196 532664 206836 532692
rect 179196 532652 179202 532664
rect 206830 532652 206836 532664
rect 206888 532652 206894 532704
rect 83090 532040 83096 532092
rect 83148 532080 83154 532092
rect 109678 532080 109684 532092
rect 83148 532052 109684 532080
rect 83148 532040 83154 532052
rect 109678 532040 109684 532052
rect 109736 532040 109742 532092
rect 244366 532040 244372 532092
rect 244424 532080 244430 532092
rect 266538 532080 266544 532092
rect 244424 532052 266544 532080
rect 244424 532040 244430 532052
rect 266538 532040 266544 532052
rect 266596 532040 266602 532092
rect 48222 531972 48228 532024
rect 48280 532012 48286 532024
rect 96890 532012 96896 532024
rect 48280 531984 96896 532012
rect 48280 531972 48286 531984
rect 96890 531972 96896 531984
rect 96948 531972 96954 532024
rect 100018 531972 100024 532024
rect 100076 532012 100082 532024
rect 128998 532012 129004 532024
rect 100076 531984 129004 532012
rect 100076 531972 100082 531984
rect 128998 531972 129004 531984
rect 129056 531972 129062 532024
rect 173158 531972 173164 532024
rect 173216 532012 173222 532024
rect 195422 532012 195428 532024
rect 173216 531984 195428 532012
rect 173216 531972 173222 531984
rect 195422 531972 195428 531984
rect 195480 531972 195486 532024
rect 202966 531972 202972 532024
rect 203024 532012 203030 532024
rect 270586 532012 270592 532024
rect 203024 531984 270592 532012
rect 203024 531972 203030 531984
rect 270586 531972 270592 531984
rect 270644 531972 270650 532024
rect 93118 531292 93124 531344
rect 93176 531332 93182 531344
rect 94038 531332 94044 531344
rect 93176 531304 94044 531332
rect 93176 531292 93182 531304
rect 94038 531292 94044 531304
rect 94096 531292 94102 531344
rect 183370 530612 183376 530664
rect 183428 530652 183434 530664
rect 254210 530652 254216 530664
rect 183428 530624 254216 530652
rect 183428 530612 183434 530624
rect 254210 530612 254216 530624
rect 254268 530612 254274 530664
rect 81986 530544 81992 530596
rect 82044 530584 82050 530596
rect 187602 530584 187608 530596
rect 82044 530556 187608 530584
rect 82044 530544 82050 530556
rect 187602 530544 187608 530556
rect 187660 530544 187666 530596
rect 193030 530544 193036 530596
rect 193088 530584 193094 530596
rect 200206 530584 200212 530596
rect 193088 530556 200212 530584
rect 193088 530544 193094 530556
rect 200206 530544 200212 530556
rect 200264 530544 200270 530596
rect 207658 530544 207664 530596
rect 207716 530584 207722 530596
rect 222286 530584 222292 530596
rect 207716 530556 222292 530584
rect 207716 530544 207722 530556
rect 222286 530544 222292 530556
rect 222344 530544 222350 530596
rect 231210 530544 231216 530596
rect 231268 530584 231274 530596
rect 260926 530584 260932 530596
rect 231268 530556 260932 530584
rect 231268 530544 231274 530556
rect 260926 530544 260932 530556
rect 260984 530544 260990 530596
rect 204622 529184 204628 529236
rect 204680 529224 204686 529236
rect 238018 529224 238024 529236
rect 204680 529196 238024 529224
rect 204680 529184 204686 529196
rect 238018 529184 238024 529196
rect 238076 529184 238082 529236
rect 248506 529184 248512 529236
rect 248564 529224 248570 529236
rect 280246 529224 280252 529236
rect 248564 529196 280252 529224
rect 248564 529184 248570 529196
rect 280246 529184 280252 529196
rect 280304 529184 280310 529236
rect 226242 528572 226248 528624
rect 226300 528612 226306 528624
rect 229094 528612 229100 528624
rect 226300 528584 229100 528612
rect 226300 528572 226306 528584
rect 229094 528572 229100 528584
rect 229152 528572 229158 528624
rect 59262 528504 59268 528556
rect 59320 528544 59326 528556
rect 169754 528544 169760 528556
rect 59320 528516 169760 528544
rect 59320 528504 59326 528516
rect 169754 528504 169760 528516
rect 169812 528544 169818 528556
rect 170490 528544 170496 528556
rect 169812 528516 170496 528544
rect 169812 528504 169818 528516
rect 170490 528504 170496 528516
rect 170548 528504 170554 528556
rect 3418 528436 3424 528488
rect 3476 528476 3482 528488
rect 97994 528476 98000 528488
rect 3476 528448 98000 528476
rect 3476 528436 3482 528448
rect 97994 528436 98000 528448
rect 98052 528436 98058 528488
rect 193122 527892 193128 527944
rect 193180 527932 193186 527944
rect 205634 527932 205640 527944
rect 193180 527904 205640 527932
rect 193180 527892 193186 527904
rect 205634 527892 205640 527904
rect 205692 527892 205698 527944
rect 245654 527892 245660 527944
rect 245712 527932 245718 527944
rect 258258 527932 258264 527944
rect 245712 527904 258264 527932
rect 245712 527892 245718 527904
rect 258258 527892 258264 527904
rect 258316 527892 258322 527944
rect 201586 527824 201592 527876
rect 201644 527864 201650 527876
rect 248506 527864 248512 527876
rect 201644 527836 248512 527864
rect 201644 527824 201650 527836
rect 248506 527824 248512 527836
rect 248564 527824 248570 527876
rect 88334 527076 88340 527128
rect 88392 527116 88398 527128
rect 208486 527116 208492 527128
rect 88392 527088 208492 527116
rect 88392 527076 88398 527088
rect 208486 527076 208492 527088
rect 208544 527076 208550 527128
rect 243538 526464 243544 526516
rect 243596 526504 243602 526516
rect 254026 526504 254032 526516
rect 243596 526476 254032 526504
rect 243596 526464 243602 526476
rect 254026 526464 254032 526476
rect 254084 526464 254090 526516
rect 188982 526396 188988 526448
rect 189040 526436 189046 526448
rect 193306 526436 193312 526448
rect 189040 526408 193312 526436
rect 189040 526396 189046 526408
rect 193306 526396 193312 526408
rect 193364 526396 193370 526448
rect 202138 526396 202144 526448
rect 202196 526436 202202 526448
rect 227806 526436 227812 526448
rect 202196 526408 227812 526436
rect 202196 526396 202202 526408
rect 227806 526396 227812 526408
rect 227864 526396 227870 526448
rect 229830 526396 229836 526448
rect 229888 526436 229894 526448
rect 251266 526436 251272 526448
rect 229888 526408 251272 526436
rect 229888 526396 229894 526408
rect 251266 526396 251272 526408
rect 251324 526396 251330 526448
rect 131022 525104 131028 525156
rect 131080 525144 131086 525156
rect 182910 525144 182916 525156
rect 131080 525116 182916 525144
rect 131080 525104 131086 525116
rect 182910 525104 182916 525116
rect 182968 525104 182974 525156
rect 195974 525104 195980 525156
rect 196032 525144 196038 525156
rect 220078 525144 220084 525156
rect 196032 525116 220084 525144
rect 196032 525104 196038 525116
rect 220078 525104 220084 525116
rect 220136 525104 220142 525156
rect 234706 525104 234712 525156
rect 234764 525144 234770 525156
rect 254670 525144 254676 525156
rect 234764 525116 254676 525144
rect 234764 525104 234770 525116
rect 254670 525104 254676 525116
rect 254728 525104 254734 525156
rect 71866 525036 71872 525088
rect 71924 525076 71930 525088
rect 122834 525076 122840 525088
rect 71924 525048 122840 525076
rect 71924 525036 71930 525048
rect 122834 525036 122840 525048
rect 122892 525036 122898 525088
rect 172330 525036 172336 525088
rect 172388 525076 172394 525088
rect 239398 525076 239404 525088
rect 172388 525048 239404 525076
rect 172388 525036 172394 525048
rect 239398 525036 239404 525048
rect 239456 525036 239462 525088
rect 71038 523676 71044 523728
rect 71096 523716 71102 523728
rect 118694 523716 118700 523728
rect 71096 523688 118700 523716
rect 71096 523676 71102 523688
rect 118694 523676 118700 523688
rect 118752 523676 118758 523728
rect 199378 523676 199384 523728
rect 199436 523716 199442 523728
rect 208394 523716 208400 523728
rect 199436 523688 208400 523716
rect 199436 523676 199442 523688
rect 208394 523676 208400 523688
rect 208452 523676 208458 523728
rect 233326 523676 233332 523728
rect 233384 523716 233390 523728
rect 251266 523716 251272 523728
rect 233384 523688 251272 523716
rect 233384 523676 233390 523688
rect 251266 523676 251272 523688
rect 251324 523676 251330 523728
rect 63310 522928 63316 522980
rect 63368 522968 63374 522980
rect 162210 522968 162216 522980
rect 63368 522940 162216 522968
rect 63368 522928 63374 522940
rect 162210 522928 162216 522940
rect 162268 522928 162274 522980
rect 3418 522248 3424 522300
rect 3476 522288 3482 522300
rect 93118 522288 93124 522300
rect 3476 522260 93124 522288
rect 3476 522248 3482 522260
rect 93118 522248 93124 522260
rect 93176 522288 93182 522300
rect 94498 522288 94504 522300
rect 93176 522260 94504 522288
rect 93176 522248 93182 522260
rect 94498 522248 94504 522260
rect 94556 522248 94562 522300
rect 195238 522248 195244 522300
rect 195296 522288 195302 522300
rect 204438 522288 204444 522300
rect 195296 522260 204444 522288
rect 195296 522248 195302 522260
rect 204438 522248 204444 522260
rect 204496 522248 204502 522300
rect 144822 519528 144828 519580
rect 144880 519568 144886 519580
rect 244918 519568 244924 519580
rect 144880 519540 244924 519568
rect 144880 519528 144886 519540
rect 244918 519528 244924 519540
rect 244976 519528 244982 519580
rect 72418 518168 72424 518220
rect 72476 518208 72482 518220
rect 99374 518208 99380 518220
rect 72476 518180 99380 518208
rect 72476 518168 72482 518180
rect 99374 518168 99380 518180
rect 99432 518168 99438 518220
rect 141970 518168 141976 518220
rect 142028 518208 142034 518220
rect 216766 518208 216772 518220
rect 142028 518180 216772 518208
rect 142028 518168 142034 518180
rect 216766 518168 216772 518180
rect 216824 518168 216830 518220
rect 218698 518168 218704 518220
rect 218756 518208 218762 518220
rect 237466 518208 237472 518220
rect 218756 518180 237472 518208
rect 218756 518168 218762 518180
rect 237466 518168 237472 518180
rect 237524 518168 237530 518220
rect 65978 517216 65984 517268
rect 66036 517256 66042 517268
rect 69658 517256 69664 517268
rect 66036 517228 69664 517256
rect 66036 517216 66042 517228
rect 69658 517216 69664 517228
rect 69716 517216 69722 517268
rect 210418 516808 210424 516860
rect 210476 516848 210482 516860
rect 253934 516848 253940 516860
rect 210476 516820 253940 516848
rect 210476 516808 210482 516820
rect 253934 516808 253940 516820
rect 253992 516808 253998 516860
rect 158438 516740 158444 516792
rect 158496 516780 158502 516792
rect 238754 516780 238760 516792
rect 158496 516752 238760 516780
rect 158496 516740 158502 516752
rect 238754 516740 238760 516752
rect 238812 516740 238818 516792
rect 61930 515380 61936 515432
rect 61988 515420 61994 515432
rect 92566 515420 92572 515432
rect 61988 515392 92572 515420
rect 61988 515380 61994 515392
rect 92566 515380 92572 515392
rect 92624 515380 92630 515432
rect 181990 515380 181996 515432
rect 182048 515420 182054 515432
rect 216030 515420 216036 515432
rect 182048 515392 216036 515420
rect 182048 515380 182054 515392
rect 216030 515380 216036 515392
rect 216088 515380 216094 515432
rect 237558 515380 237564 515432
rect 237616 515420 237622 515432
rect 254578 515420 254584 515432
rect 237616 515392 254584 515420
rect 237616 515380 237622 515392
rect 254578 515380 254584 515392
rect 254636 515380 254642 515432
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 193122 514088 193128 514140
rect 193180 514128 193186 514140
rect 205726 514128 205732 514140
rect 193180 514100 205732 514128
rect 193180 514088 193186 514100
rect 205726 514088 205732 514100
rect 205784 514088 205790 514140
rect 145650 514020 145656 514072
rect 145708 514060 145714 514072
rect 234614 514060 234620 514072
rect 145708 514032 234620 514060
rect 145708 514020 145714 514032
rect 234614 514020 234620 514032
rect 234672 514020 234678 514072
rect 236086 513272 236092 513324
rect 236144 513312 236150 513324
rect 238110 513312 238116 513324
rect 236144 513284 238116 513312
rect 236144 513272 236150 513284
rect 238110 513272 238116 513284
rect 238168 513272 238174 513324
rect 184658 512592 184664 512644
rect 184716 512632 184722 512644
rect 246390 512632 246396 512644
rect 184716 512604 246396 512632
rect 184716 512592 184722 512604
rect 246390 512592 246396 512604
rect 246448 512592 246454 512644
rect 50982 511912 50988 511964
rect 51040 511952 51046 511964
rect 168834 511952 168840 511964
rect 51040 511924 168840 511952
rect 51040 511912 51046 511924
rect 168834 511912 168840 511924
rect 168892 511912 168898 511964
rect 168834 511232 168840 511284
rect 168892 511272 168898 511284
rect 169570 511272 169576 511284
rect 168892 511244 169576 511272
rect 168892 511232 168898 511244
rect 169570 511232 169576 511244
rect 169628 511272 169634 511284
rect 198090 511272 198096 511284
rect 169628 511244 198096 511272
rect 169628 511232 169634 511244
rect 198090 511232 198096 511244
rect 198148 511232 198154 511284
rect 165062 509872 165068 509924
rect 165120 509912 165126 509924
rect 214006 509912 214012 509924
rect 165120 509884 214012 509912
rect 165120 509872 165126 509884
rect 214006 509872 214012 509884
rect 214064 509872 214070 509924
rect 154482 508512 154488 508564
rect 154540 508552 154546 508564
rect 229830 508552 229836 508564
rect 154540 508524 229836 508552
rect 154540 508512 154546 508524
rect 229830 508512 229836 508524
rect 229888 508512 229894 508564
rect 139302 507084 139308 507136
rect 139360 507124 139366 507136
rect 267918 507124 267924 507136
rect 139360 507096 267924 507124
rect 139360 507084 139366 507096
rect 267918 507084 267924 507096
rect 267976 507084 267982 507136
rect 187510 505792 187516 505844
rect 187568 505832 187574 505844
rect 214558 505832 214564 505844
rect 187568 505804 214564 505832
rect 187568 505792 187574 505804
rect 214558 505792 214564 505804
rect 214616 505792 214622 505844
rect 136542 505724 136548 505776
rect 136600 505764 136606 505776
rect 219434 505764 219440 505776
rect 136600 505736 219440 505764
rect 136600 505724 136606 505736
rect 219434 505724 219440 505736
rect 219492 505724 219498 505776
rect 186958 504432 186964 504484
rect 187016 504472 187022 504484
rect 244458 504472 244464 504484
rect 187016 504444 244464 504472
rect 187016 504432 187022 504444
rect 244458 504432 244464 504444
rect 244516 504432 244522 504484
rect 143350 504364 143356 504416
rect 143408 504404 143414 504416
rect 231946 504404 231952 504416
rect 143408 504376 231952 504404
rect 143408 504364 143414 504376
rect 231946 504364 231952 504376
rect 232004 504364 232010 504416
rect 189718 503004 189724 503056
rect 189776 503044 189782 503056
rect 215938 503044 215944 503056
rect 189776 503016 215944 503044
rect 189776 503004 189782 503016
rect 215938 503004 215944 503016
rect 215996 503004 216002 503056
rect 205082 502936 205088 502988
rect 205140 502976 205146 502988
rect 240226 502976 240232 502988
rect 205140 502948 240232 502976
rect 205140 502936 205146 502948
rect 240226 502936 240232 502948
rect 240284 502936 240290 502988
rect 76006 502256 76012 502308
rect 76064 502296 76070 502308
rect 77202 502296 77208 502308
rect 76064 502268 77208 502296
rect 76064 502256 76070 502268
rect 77202 502256 77208 502268
rect 77260 502256 77266 502308
rect 212626 501712 212632 501764
rect 212684 501752 212690 501764
rect 213270 501752 213276 501764
rect 212684 501724 213276 501752
rect 212684 501712 212690 501724
rect 213270 501712 213276 501724
rect 213328 501712 213334 501764
rect 188430 501644 188436 501696
rect 188488 501684 188494 501696
rect 262398 501684 262404 501696
rect 188488 501656 262404 501684
rect 188488 501644 188494 501656
rect 262398 501644 262404 501656
rect 262456 501644 262462 501696
rect 77202 501576 77208 501628
rect 77260 501616 77266 501628
rect 212626 501616 212632 501628
rect 77260 501588 212632 501616
rect 77260 501576 77266 501588
rect 212626 501576 212632 501588
rect 212684 501576 212690 501628
rect 142062 500216 142068 500268
rect 142120 500256 142126 500268
rect 250438 500256 250444 500268
rect 142120 500228 250444 500256
rect 142120 500216 142126 500228
rect 250438 500216 250444 500228
rect 250496 500216 250502 500268
rect 155678 498788 155684 498840
rect 155736 498828 155742 498840
rect 229738 498828 229744 498840
rect 155736 498800 229744 498828
rect 155736 498788 155742 498800
rect 229738 498788 229744 498800
rect 229796 498788 229802 498840
rect 242894 498788 242900 498840
rect 242952 498828 242958 498840
rect 291378 498828 291384 498840
rect 242952 498800 291384 498828
rect 242952 498788 242958 498800
rect 291378 498788 291384 498800
rect 291436 498788 291442 498840
rect 192570 497428 192576 497480
rect 192628 497468 192634 497480
rect 203518 497468 203524 497480
rect 192628 497440 203524 497468
rect 192628 497428 192634 497440
rect 203518 497428 203524 497440
rect 203576 497428 203582 497480
rect 220814 497428 220820 497480
rect 220872 497468 220878 497480
rect 256786 497468 256792 497480
rect 220872 497440 256792 497468
rect 220872 497428 220878 497440
rect 256786 497428 256792 497440
rect 256844 497428 256850 497480
rect 162670 496068 162676 496120
rect 162728 496108 162734 496120
rect 254118 496108 254124 496120
rect 162728 496080 254124 496108
rect 162728 496068 162734 496080
rect 254118 496068 254124 496080
rect 254176 496068 254182 496120
rect 244366 495456 244372 495508
rect 244424 495496 244430 495508
rect 298094 495496 298100 495508
rect 244424 495468 298100 495496
rect 244424 495456 244430 495468
rect 298094 495456 298100 495468
rect 298152 495456 298158 495508
rect 127618 494708 127624 494760
rect 127676 494748 127682 494760
rect 244366 494748 244372 494760
rect 127676 494720 244372 494748
rect 127676 494708 127682 494720
rect 244366 494708 244372 494720
rect 244424 494708 244430 494760
rect 242894 493960 242900 494012
rect 242952 494000 242958 494012
rect 243538 494000 243544 494012
rect 242952 493972 243544 494000
rect 242952 493960 242958 493972
rect 243538 493960 243544 493972
rect 243596 493960 243602 494012
rect 246298 493348 246304 493400
rect 246356 493388 246362 493400
rect 251818 493388 251824 493400
rect 246356 493360 251824 493388
rect 246356 493348 246362 493360
rect 251818 493348 251824 493360
rect 251876 493348 251882 493400
rect 163958 493280 163964 493332
rect 164016 493320 164022 493332
rect 206370 493320 206376 493332
rect 164016 493292 206376 493320
rect 164016 493280 164022 493292
rect 206370 493280 206376 493292
rect 206428 493280 206434 493332
rect 223482 493280 223488 493332
rect 223540 493320 223546 493332
rect 253382 493320 253388 493332
rect 223540 493292 253388 493320
rect 223540 493280 223546 493292
rect 253382 493280 253388 493292
rect 253440 493280 253446 493332
rect 132402 492668 132408 492720
rect 132460 492708 132466 492720
rect 242894 492708 242900 492720
rect 132460 492680 242900 492708
rect 132460 492668 132466 492680
rect 242894 492668 242900 492680
rect 242952 492668 242958 492720
rect 196618 491988 196624 492040
rect 196676 492028 196682 492040
rect 218698 492028 218704 492040
rect 196676 492000 218704 492028
rect 196676 491988 196682 492000
rect 218698 491988 218704 492000
rect 218756 491988 218762 492040
rect 171870 491920 171876 491972
rect 171928 491960 171934 491972
rect 213178 491960 213184 491972
rect 171928 491932 213184 491960
rect 171928 491920 171934 491932
rect 213178 491920 213184 491932
rect 213236 491920 213242 491972
rect 222102 491920 222108 491972
rect 222160 491960 222166 491972
rect 247126 491960 247132 491972
rect 222160 491932 247132 491960
rect 222160 491920 222166 491932
rect 247126 491920 247132 491932
rect 247184 491920 247190 491972
rect 239398 491308 239404 491360
rect 239456 491348 239462 491360
rect 241422 491348 241428 491360
rect 239456 491320 241428 491348
rect 239456 491308 239462 491320
rect 241422 491308 241428 491320
rect 241480 491308 241486 491360
rect 198090 490628 198096 490680
rect 198148 490668 198154 490680
rect 215938 490668 215944 490680
rect 198148 490640 215944 490668
rect 198148 490628 198154 490640
rect 215938 490628 215944 490640
rect 215996 490628 216002 490680
rect 176102 490560 176108 490612
rect 176160 490600 176166 490612
rect 200298 490600 200304 490612
rect 176160 490572 200304 490600
rect 176160 490560 176166 490572
rect 200298 490560 200304 490572
rect 200356 490560 200362 490612
rect 142890 488520 142896 488572
rect 142948 488560 142954 488572
rect 143442 488560 143448 488572
rect 142948 488532 143448 488560
rect 142948 488520 142954 488532
rect 143442 488520 143448 488532
rect 143500 488560 143506 488572
rect 232590 488560 232596 488572
rect 143500 488532 232596 488560
rect 143500 488520 143506 488532
rect 232590 488520 232596 488532
rect 232648 488520 232654 488572
rect 104250 488452 104256 488504
rect 104308 488492 104314 488504
rect 198826 488492 198832 488504
rect 104308 488464 198832 488492
rect 104308 488452 104314 488464
rect 198826 488452 198832 488464
rect 198884 488452 198890 488504
rect 226978 488180 226984 488232
rect 227036 488220 227042 488232
rect 229094 488220 229100 488232
rect 227036 488192 229100 488220
rect 227036 488180 227042 488192
rect 229094 488180 229100 488192
rect 229152 488180 229158 488232
rect 198826 487840 198832 487892
rect 198884 487880 198890 487892
rect 227070 487880 227076 487892
rect 198884 487852 227076 487880
rect 198884 487840 198890 487852
rect 227070 487840 227076 487852
rect 227128 487840 227134 487892
rect 174998 487772 175004 487824
rect 175056 487812 175062 487824
rect 198734 487812 198740 487824
rect 175056 487784 198740 487812
rect 175056 487772 175062 487784
rect 198734 487772 198740 487784
rect 198792 487772 198798 487824
rect 199470 487772 199476 487824
rect 199528 487812 199534 487824
rect 241606 487812 241612 487824
rect 199528 487784 241612 487812
rect 199528 487772 199534 487784
rect 241606 487772 241612 487784
rect 241664 487772 241670 487824
rect 104250 487160 104256 487212
rect 104308 487200 104314 487212
rect 104802 487200 104808 487212
rect 104308 487172 104808 487200
rect 104308 487160 104314 487172
rect 104802 487160 104808 487172
rect 104860 487160 104866 487212
rect 160002 486412 160008 486464
rect 160060 486452 160066 486464
rect 174538 486452 174544 486464
rect 160060 486424 174544 486452
rect 160060 486412 160066 486424
rect 174538 486412 174544 486424
rect 174596 486412 174602 486464
rect 179414 485732 179420 485784
rect 179472 485772 179478 485784
rect 180518 485772 180524 485784
rect 179472 485744 180524 485772
rect 179472 485732 179478 485744
rect 180518 485732 180524 485744
rect 180576 485772 180582 485784
rect 580166 485772 580172 485784
rect 180576 485744 580172 485772
rect 180576 485732 180582 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 153102 485052 153108 485104
rect 153160 485092 153166 485104
rect 179414 485092 179420 485104
rect 153160 485064 179420 485092
rect 153160 485052 153166 485064
rect 179414 485052 179420 485064
rect 179472 485052 179478 485104
rect 144730 484372 144736 484424
rect 144788 484412 144794 484424
rect 241422 484412 241428 484424
rect 144788 484384 241428 484412
rect 144788 484372 144794 484384
rect 241422 484372 241428 484384
rect 241480 484412 241486 484424
rect 252554 484412 252560 484424
rect 241480 484384 252560 484412
rect 241480 484372 241486 484384
rect 252554 484372 252560 484384
rect 252612 484372 252618 484424
rect 93946 483624 93952 483676
rect 94004 483664 94010 483676
rect 94590 483664 94596 483676
rect 94004 483636 94596 483664
rect 94004 483624 94010 483636
rect 94590 483624 94596 483636
rect 94648 483664 94654 483676
rect 209866 483664 209872 483676
rect 94648 483636 209872 483664
rect 94648 483624 94654 483636
rect 209866 483624 209872 483636
rect 209924 483664 209930 483676
rect 210602 483664 210608 483676
rect 209924 483636 210608 483664
rect 209924 483624 209930 483636
rect 210602 483624 210608 483636
rect 210660 483624 210666 483676
rect 226150 482944 226156 482996
rect 226208 482984 226214 482996
rect 226334 482984 226340 482996
rect 226208 482956 226340 482984
rect 226208 482944 226214 482956
rect 226334 482944 226340 482956
rect 226392 482944 226398 482996
rect 226426 481652 226432 481704
rect 226484 481692 226490 481704
rect 245562 481692 245568 481704
rect 226484 481664 245568 481692
rect 226484 481652 226490 481664
rect 245562 481652 245568 481664
rect 245620 481692 245626 481704
rect 248414 481692 248420 481704
rect 245620 481664 248420 481692
rect 245620 481652 245626 481664
rect 248414 481652 248420 481664
rect 248472 481652 248478 481704
rect 192478 480904 192484 480956
rect 192536 480944 192542 480956
rect 215294 480944 215300 480956
rect 192536 480916 215300 480944
rect 192536 480904 192542 480916
rect 215294 480904 215300 480916
rect 215352 480904 215358 480956
rect 146938 480224 146944 480276
rect 146996 480264 147002 480276
rect 240778 480264 240784 480276
rect 146996 480236 240784 480264
rect 146996 480224 147002 480236
rect 240778 480224 240784 480236
rect 240836 480224 240842 480276
rect 175090 479544 175096 479596
rect 175148 479584 175154 479596
rect 202138 479584 202144 479596
rect 175148 479556 202144 479584
rect 175148 479544 175154 479556
rect 202138 479544 202144 479556
rect 202196 479544 202202 479596
rect 210602 479544 210608 479596
rect 210660 479584 210666 479596
rect 227806 479584 227812 479596
rect 210660 479556 227812 479584
rect 210660 479544 210666 479556
rect 227806 479544 227812 479556
rect 227864 479544 227870 479596
rect 233234 479544 233240 479596
rect 233292 479584 233298 479596
rect 252554 479584 252560 479596
rect 233292 479556 252560 479584
rect 233292 479544 233298 479556
rect 252554 479544 252560 479556
rect 252612 479544 252618 479596
rect 111058 479476 111064 479528
rect 111116 479516 111122 479528
rect 251266 479516 251272 479528
rect 111116 479488 251272 479516
rect 111116 479476 111122 479488
rect 251266 479476 251272 479488
rect 251324 479476 251330 479528
rect 110414 478864 110420 478916
rect 110472 478904 110478 478916
rect 111058 478904 111064 478916
rect 110472 478876 111064 478904
rect 110472 478864 110478 478876
rect 111058 478864 111064 478876
rect 111116 478864 111122 478916
rect 251266 478864 251272 478916
rect 251324 478904 251330 478916
rect 251910 478904 251916 478916
rect 251324 478876 251916 478904
rect 251324 478864 251330 478876
rect 251910 478864 251916 478876
rect 251968 478864 251974 478916
rect 168098 478184 168104 478236
rect 168156 478224 168162 478236
rect 211154 478224 211160 478236
rect 168156 478196 211160 478224
rect 168156 478184 168162 478196
rect 211154 478184 211160 478196
rect 211212 478184 211218 478236
rect 35158 478116 35164 478168
rect 35216 478156 35222 478168
rect 43438 478156 43444 478168
rect 35216 478128 43444 478156
rect 35216 478116 35222 478128
rect 43438 478116 43444 478128
rect 43496 478116 43502 478168
rect 126238 478116 126244 478168
rect 126296 478156 126302 478168
rect 208486 478156 208492 478168
rect 126296 478128 208492 478156
rect 126296 478116 126302 478128
rect 208486 478116 208492 478128
rect 208544 478156 208550 478168
rect 277670 478156 277676 478168
rect 208544 478128 277676 478156
rect 208544 478116 208550 478128
rect 277670 478116 277676 478128
rect 277728 478116 277734 478168
rect 218146 476824 218152 476876
rect 218204 476864 218210 476876
rect 250438 476864 250444 476876
rect 218204 476836 250444 476864
rect 218204 476824 218210 476836
rect 250438 476824 250444 476836
rect 250496 476824 250502 476876
rect 85482 476756 85488 476808
rect 85540 476796 85546 476808
rect 94130 476796 94136 476808
rect 85540 476768 94136 476796
rect 85540 476756 85546 476768
rect 94130 476756 94136 476768
rect 94188 476756 94194 476808
rect 102134 476756 102140 476808
rect 102192 476796 102198 476808
rect 102778 476796 102784 476808
rect 102192 476768 102784 476796
rect 102192 476756 102198 476768
rect 102778 476756 102784 476768
rect 102836 476796 102842 476808
rect 259638 476796 259644 476808
rect 102836 476768 259644 476796
rect 102836 476756 102842 476768
rect 259638 476756 259644 476768
rect 259696 476756 259702 476808
rect 3326 475328 3332 475380
rect 3384 475368 3390 475380
rect 35158 475368 35164 475380
rect 3384 475340 35164 475368
rect 3384 475328 3390 475340
rect 35158 475328 35164 475340
rect 35216 475328 35222 475380
rect 133138 475192 133144 475244
rect 133196 475232 133202 475244
rect 133690 475232 133696 475244
rect 133196 475204 133696 475232
rect 133196 475192 133202 475204
rect 133690 475192 133696 475204
rect 133748 475192 133754 475244
rect 106918 474784 106924 474836
rect 106976 474824 106982 474836
rect 241698 474824 241704 474836
rect 106976 474796 241704 474824
rect 106976 474784 106982 474796
rect 241698 474784 241704 474796
rect 241756 474824 241762 474836
rect 242158 474824 242164 474836
rect 241756 474796 242164 474824
rect 241756 474784 241762 474796
rect 242158 474784 242164 474796
rect 242216 474784 242222 474836
rect 133690 474716 133696 474768
rect 133748 474756 133754 474768
rect 291286 474756 291292 474768
rect 133748 474728 291292 474756
rect 133748 474716 133754 474728
rect 291286 474716 291292 474728
rect 291344 474716 291350 474768
rect 240134 473968 240140 474020
rect 240192 474008 240198 474020
rect 256878 474008 256884 474020
rect 240192 473980 256884 474008
rect 240192 473968 240198 473980
rect 256878 473968 256884 473980
rect 256936 473968 256942 474020
rect 133230 473356 133236 473408
rect 133288 473396 133294 473408
rect 270586 473396 270592 473408
rect 133288 473368 270592 473396
rect 133288 473356 133294 473368
rect 270586 473356 270592 473368
rect 270644 473356 270650 473408
rect 79962 472608 79968 472660
rect 80020 472648 80026 472660
rect 101398 472648 101404 472660
rect 80020 472620 101404 472648
rect 80020 472608 80026 472620
rect 101398 472608 101404 472620
rect 101456 472608 101462 472660
rect 148318 472064 148324 472116
rect 148376 472104 148382 472116
rect 229094 472104 229100 472116
rect 148376 472076 229100 472104
rect 148376 472064 148382 472076
rect 229094 472064 229100 472076
rect 229152 472104 229158 472116
rect 284478 472104 284484 472116
rect 229152 472076 284484 472104
rect 229152 472064 229158 472076
rect 284478 472064 284484 472076
rect 284536 472064 284542 472116
rect 105538 471996 105544 472048
rect 105596 472036 105602 472048
rect 258074 472036 258080 472048
rect 105596 472008 258080 472036
rect 105596 471996 105602 472008
rect 258074 471996 258080 472008
rect 258132 471996 258138 472048
rect 216766 471316 216772 471368
rect 216824 471356 216830 471368
rect 265066 471356 265072 471368
rect 216824 471328 265072 471356
rect 216824 471316 216830 471328
rect 265066 471316 265072 471328
rect 265124 471316 265130 471368
rect 79318 471248 79324 471300
rect 79376 471288 79382 471300
rect 91186 471288 91192 471300
rect 79376 471260 91192 471288
rect 79376 471248 79382 471260
rect 91186 471248 91192 471260
rect 91244 471248 91250 471300
rect 111058 471248 111064 471300
rect 111116 471288 111122 471300
rect 158714 471288 158720 471300
rect 111116 471260 158720 471288
rect 111116 471248 111122 471260
rect 158714 471248 158720 471260
rect 158772 471248 158778 471300
rect 166810 471248 166816 471300
rect 166868 471288 166874 471300
rect 169478 471288 169484 471300
rect 166868 471260 169484 471288
rect 166868 471248 166874 471260
rect 169478 471248 169484 471260
rect 169536 471288 169542 471300
rect 255498 471288 255504 471300
rect 169536 471260 255504 471288
rect 169536 471248 169542 471260
rect 255498 471248 255504 471260
rect 255556 471248 255562 471300
rect 116578 469820 116584 469872
rect 116636 469860 116642 469872
rect 150158 469860 150164 469872
rect 116636 469832 150164 469860
rect 116636 469820 116642 469832
rect 150158 469820 150164 469832
rect 150216 469860 150222 469872
rect 281626 469860 281632 469872
rect 150216 469832 281632 469860
rect 150216 469820 150222 469832
rect 281626 469820 281632 469832
rect 281684 469820 281690 469872
rect 90358 469208 90364 469260
rect 90416 469248 90422 469260
rect 91002 469248 91008 469260
rect 90416 469220 91008 469248
rect 90416 469208 90422 469220
rect 91002 469208 91008 469220
rect 91060 469248 91066 469260
rect 187050 469248 187056 469260
rect 91060 469220 187056 469248
rect 91060 469208 91066 469220
rect 187050 469208 187056 469220
rect 187108 469208 187114 469260
rect 187602 469208 187608 469260
rect 187660 469248 187666 469260
rect 253474 469248 253480 469260
rect 187660 469220 253480 469248
rect 187660 469208 187666 469220
rect 253474 469208 253480 469220
rect 253532 469208 253538 469260
rect 180518 468528 180524 468580
rect 180576 468568 180582 468580
rect 213914 468568 213920 468580
rect 180576 468540 213920 468568
rect 180576 468528 180582 468540
rect 213914 468528 213920 468540
rect 213972 468528 213978 468580
rect 245562 468528 245568 468580
rect 245620 468568 245626 468580
rect 265710 468568 265716 468580
rect 245620 468540 265716 468568
rect 245620 468528 245626 468540
rect 265710 468528 265716 468540
rect 265768 468528 265774 468580
rect 114462 468460 114468 468512
rect 114520 468500 114526 468512
rect 258258 468500 258264 468512
rect 114520 468472 258264 468500
rect 114520 468460 114526 468472
rect 258258 468460 258264 468472
rect 258316 468460 258322 468512
rect 113818 467848 113824 467900
rect 113876 467888 113882 467900
rect 114462 467888 114468 467900
rect 113876 467860 114468 467888
rect 113876 467848 113882 467860
rect 114462 467848 114468 467860
rect 114520 467848 114526 467900
rect 149698 466488 149704 466540
rect 149756 466528 149762 466540
rect 181530 466528 181536 466540
rect 149756 466500 181536 466528
rect 149756 466488 149762 466500
rect 181530 466488 181536 466500
rect 181588 466528 181594 466540
rect 182082 466528 182088 466540
rect 181588 466500 182088 466528
rect 181588 466488 181594 466500
rect 182082 466488 182088 466500
rect 182140 466488 182146 466540
rect 227714 466488 227720 466540
rect 227772 466528 227778 466540
rect 289998 466528 290004 466540
rect 227772 466500 290004 466528
rect 227772 466488 227778 466500
rect 289998 466488 290004 466500
rect 290056 466488 290062 466540
rect 175918 466420 175924 466472
rect 175976 466460 175982 466472
rect 248414 466460 248420 466472
rect 175976 466432 248420 466460
rect 175976 466420 175982 466432
rect 248414 466420 248420 466432
rect 248472 466420 248478 466472
rect 182082 465672 182088 465724
rect 182140 465712 182146 465724
rect 215294 465712 215300 465724
rect 182140 465684 215300 465712
rect 182140 465672 182146 465684
rect 215294 465672 215300 465684
rect 215352 465672 215358 465724
rect 223574 465672 223580 465724
rect 223632 465712 223638 465724
rect 246942 465712 246948 465724
rect 223632 465684 246948 465712
rect 223632 465672 223638 465684
rect 246942 465672 246948 465684
rect 247000 465712 247006 465724
rect 262858 465712 262864 465724
rect 247000 465684 262864 465712
rect 247000 465672 247006 465684
rect 262858 465672 262864 465684
rect 262916 465672 262922 465724
rect 94498 465536 94504 465588
rect 94556 465576 94562 465588
rect 95142 465576 95148 465588
rect 94556 465548 95148 465576
rect 94556 465536 94562 465548
rect 95142 465536 95148 465548
rect 95200 465536 95206 465588
rect 95142 465060 95148 465112
rect 95200 465100 95206 465112
rect 217410 465100 217416 465112
rect 95200 465072 217416 465100
rect 95200 465060 95206 465072
rect 217410 465060 217416 465072
rect 217468 465060 217474 465112
rect 235994 465060 236000 465112
rect 236052 465100 236058 465112
rect 271966 465100 271972 465112
rect 236052 465072 271972 465100
rect 236052 465060 236058 465072
rect 271966 465060 271972 465072
rect 272024 465100 272030 465112
rect 272518 465100 272524 465112
rect 272024 465072 272524 465100
rect 272024 465060 272030 465072
rect 272518 465060 272524 465072
rect 272576 465060 272582 465112
rect 162302 464992 162308 465044
rect 162360 465032 162366 465044
rect 162762 465032 162768 465044
rect 162360 465004 162768 465032
rect 162360 464992 162366 465004
rect 162762 464992 162768 465004
rect 162820 465032 162826 465044
rect 187694 465032 187700 465044
rect 162820 465004 187700 465032
rect 162820 464992 162826 465004
rect 187694 464992 187700 465004
rect 187752 464992 187758 465044
rect 241422 464380 241428 464432
rect 241480 464420 241486 464432
rect 259638 464420 259644 464432
rect 241480 464392 259644 464420
rect 241480 464380 241486 464392
rect 259638 464380 259644 464392
rect 259696 464380 259702 464432
rect 98638 464312 98644 464364
rect 98696 464352 98702 464364
rect 162762 464352 162768 464364
rect 98696 464324 162768 464352
rect 98696 464312 98702 464324
rect 162762 464312 162768 464324
rect 162820 464312 162826 464364
rect 193030 464312 193036 464364
rect 193088 464352 193094 464364
rect 212534 464352 212540 464364
rect 193088 464324 212540 464352
rect 193088 464312 193094 464324
rect 212534 464312 212540 464324
rect 212592 464312 212598 464364
rect 227070 464312 227076 464364
rect 227128 464352 227134 464364
rect 245654 464352 245660 464364
rect 227128 464324 245660 464352
rect 227128 464312 227134 464324
rect 245654 464312 245660 464324
rect 245712 464312 245718 464364
rect 279418 464312 279424 464364
rect 279476 464352 279482 464364
rect 289814 464352 289820 464364
rect 279476 464324 289820 464352
rect 279476 464312 279482 464324
rect 289814 464312 289820 464324
rect 289872 464312 289878 464364
rect 159358 463700 159364 463752
rect 159416 463740 159422 463752
rect 197354 463740 197360 463752
rect 159416 463712 197360 463740
rect 159416 463700 159422 463712
rect 197354 463700 197360 463712
rect 197412 463700 197418 463752
rect 205542 462952 205548 463004
rect 205600 462992 205606 463004
rect 270494 462992 270500 463004
rect 205600 462964 270500 462992
rect 205600 462952 205606 462964
rect 270494 462952 270500 462964
rect 270552 462952 270558 463004
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 17218 462380 17224 462392
rect 3292 462352 17224 462380
rect 3292 462340 3298 462352
rect 17218 462340 17224 462352
rect 17276 462340 17282 462392
rect 112438 462340 112444 462392
rect 112496 462380 112502 462392
rect 249058 462380 249064 462392
rect 112496 462352 249064 462380
rect 112496 462340 112502 462352
rect 249058 462340 249064 462352
rect 249116 462340 249122 462392
rect 137738 461592 137744 461644
rect 137796 461632 137802 461644
rect 152550 461632 152556 461644
rect 137796 461604 152556 461632
rect 137796 461592 137802 461604
rect 152550 461592 152556 461604
rect 152608 461592 152614 461644
rect 213822 461592 213828 461644
rect 213880 461632 213886 461644
rect 278774 461632 278780 461644
rect 213880 461604 278780 461632
rect 213880 461592 213886 461604
rect 278774 461592 278780 461604
rect 278832 461592 278838 461644
rect 201494 461456 201500 461508
rect 201552 461496 201558 461508
rect 202138 461496 202144 461508
rect 201552 461468 202144 461496
rect 201552 461456 201558 461468
rect 202138 461456 202144 461468
rect 202196 461456 202202 461508
rect 185670 461320 185676 461372
rect 185728 461360 185734 461372
rect 186130 461360 186136 461372
rect 185728 461332 186136 461360
rect 185728 461320 185734 461332
rect 186130 461320 186136 461332
rect 186188 461320 186194 461372
rect 174538 460980 174544 461032
rect 174596 461020 174602 461032
rect 201494 461020 201500 461032
rect 174596 460992 201500 461020
rect 174596 460980 174602 460992
rect 201494 460980 201500 460992
rect 201552 460980 201558 461032
rect 61930 460912 61936 460964
rect 61988 460952 61994 460964
rect 74534 460952 74540 460964
rect 61988 460924 74540 460952
rect 61988 460912 61994 460924
rect 74534 460912 74540 460924
rect 74592 460912 74598 460964
rect 186130 460912 186136 460964
rect 186188 460952 186194 460964
rect 259730 460952 259736 460964
rect 186188 460924 259736 460952
rect 186188 460912 186194 460924
rect 259730 460912 259736 460924
rect 259788 460912 259794 460964
rect 85574 460844 85580 460896
rect 85632 460884 85638 460896
rect 105538 460884 105544 460896
rect 85632 460856 105544 460884
rect 85632 460844 85638 460856
rect 105538 460844 105544 460856
rect 105596 460844 105602 460896
rect 62022 460164 62028 460216
rect 62080 460204 62086 460216
rect 85666 460204 85672 460216
rect 62080 460176 85672 460204
rect 62080 460164 62086 460176
rect 85666 460164 85672 460176
rect 85724 460164 85730 460216
rect 217410 460164 217416 460216
rect 217468 460204 217474 460216
rect 233142 460204 233148 460216
rect 217468 460176 233148 460204
rect 217468 460164 217474 460176
rect 233142 460164 233148 460176
rect 233200 460164 233206 460216
rect 104894 459892 104900 459944
rect 104952 459932 104958 459944
rect 105538 459932 105544 459944
rect 104952 459904 105544 459932
rect 104952 459892 104958 459904
rect 105538 459892 105544 459904
rect 105596 459892 105602 459944
rect 137830 459620 137836 459672
rect 137888 459660 137894 459672
rect 213270 459660 213276 459672
rect 137888 459632 213276 459660
rect 137888 459620 137894 459632
rect 213270 459620 213276 459632
rect 213328 459660 213334 459672
rect 213822 459660 213828 459672
rect 213328 459632 213828 459660
rect 213328 459620 213334 459632
rect 213822 459620 213828 459632
rect 213880 459620 213886 459672
rect 215294 459620 215300 459672
rect 215352 459660 215358 459672
rect 216030 459660 216036 459672
rect 215352 459632 216036 459660
rect 215352 459620 215358 459632
rect 216030 459620 216036 459632
rect 216088 459620 216094 459672
rect 153838 459552 153844 459604
rect 153896 459592 153902 459604
rect 252554 459592 252560 459604
rect 153896 459564 252560 459592
rect 153896 459552 153902 459564
rect 252554 459552 252560 459564
rect 252612 459592 252618 459604
rect 253566 459592 253572 459604
rect 252612 459564 253572 459592
rect 252612 459552 252618 459564
rect 253566 459552 253572 459564
rect 253624 459552 253630 459604
rect 68278 458804 68284 458856
rect 68336 458844 68342 458856
rect 90358 458844 90364 458856
rect 68336 458816 90364 458844
rect 68336 458804 68342 458816
rect 90358 458804 90364 458816
rect 90416 458804 90422 458856
rect 96522 458804 96528 458856
rect 96580 458844 96586 458856
rect 142890 458844 142896 458856
rect 96580 458816 142896 458844
rect 96580 458804 96586 458816
rect 142890 458804 142896 458816
rect 142948 458804 142954 458856
rect 169478 458804 169484 458856
rect 169536 458844 169542 458856
rect 176010 458844 176016 458856
rect 169536 458816 176016 458844
rect 169536 458804 169542 458816
rect 176010 458804 176016 458816
rect 176068 458804 176074 458856
rect 241514 458804 241520 458856
rect 241572 458844 241578 458856
rect 254302 458844 254308 458856
rect 241572 458816 254308 458844
rect 241572 458804 241578 458816
rect 254302 458804 254308 458816
rect 254360 458804 254366 458856
rect 254670 458804 254676 458856
rect 254728 458844 254734 458856
rect 270494 458844 270500 458856
rect 254728 458816 270500 458844
rect 254728 458804 254734 458816
rect 270494 458804 270500 458816
rect 270552 458804 270558 458856
rect 204530 458600 204536 458652
rect 204588 458640 204594 458652
rect 205542 458640 205548 458652
rect 204588 458612 205548 458640
rect 204588 458600 204594 458612
rect 205542 458600 205548 458612
rect 205600 458600 205606 458652
rect 52178 458260 52184 458312
rect 52236 458300 52242 458312
rect 149790 458300 149796 458312
rect 52236 458272 149796 458300
rect 52236 458260 52242 458272
rect 149790 458260 149796 458272
rect 149848 458260 149854 458312
rect 178678 458260 178684 458312
rect 178736 458300 178742 458312
rect 204530 458300 204536 458312
rect 178736 458272 204536 458300
rect 178736 458260 178742 458272
rect 204530 458260 204536 458272
rect 204588 458260 204594 458312
rect 142982 458192 142988 458244
rect 143040 458232 143046 458244
rect 247402 458232 247408 458244
rect 143040 458204 247408 458232
rect 143040 458192 143046 458204
rect 247402 458192 247408 458204
rect 247460 458232 247466 458244
rect 247460 458204 248414 458232
rect 247460 458192 247466 458204
rect 248386 458164 248414 458204
rect 277578 458164 277584 458176
rect 248386 458136 277584 458164
rect 277578 458124 277584 458136
rect 277636 458124 277642 458176
rect 214558 457512 214564 457564
rect 214616 457552 214622 457564
rect 234430 457552 234436 457564
rect 214616 457524 234436 457552
rect 214616 457512 214622 457524
rect 234430 457512 234436 457524
rect 234488 457512 234494 457564
rect 162762 457444 162768 457496
rect 162820 457484 162826 457496
rect 173710 457484 173716 457496
rect 162820 457456 173716 457484
rect 162820 457444 162826 457456
rect 173710 457444 173716 457456
rect 173768 457484 173774 457496
rect 218882 457484 218888 457496
rect 173768 457456 218888 457484
rect 173768 457444 173774 457456
rect 218882 457444 218888 457456
rect 218940 457444 218946 457496
rect 70302 456764 70308 456816
rect 70360 456804 70366 456816
rect 194594 456804 194600 456816
rect 70360 456776 194600 456804
rect 70360 456764 70366 456776
rect 194594 456764 194600 456776
rect 194652 456804 194658 456816
rect 195054 456804 195060 456816
rect 194652 456776 195060 456804
rect 194652 456764 194658 456776
rect 195054 456764 195060 456776
rect 195112 456764 195118 456816
rect 225046 456764 225052 456816
rect 225104 456804 225110 456816
rect 226150 456804 226156 456816
rect 225104 456776 226156 456804
rect 225104 456764 225110 456776
rect 226150 456764 226156 456776
rect 226208 456804 226214 456816
rect 302326 456804 302332 456816
rect 226208 456776 302332 456804
rect 226208 456764 226214 456776
rect 302326 456764 302332 456776
rect 302384 456764 302390 456816
rect 288342 456016 288348 456068
rect 288400 456056 288406 456068
rect 580166 456056 580172 456068
rect 288400 456028 580172 456056
rect 288400 456016 288406 456028
rect 580166 456016 580172 456028
rect 580224 456016 580230 456068
rect 238754 455880 238760 455932
rect 238812 455920 238818 455932
rect 239398 455920 239404 455932
rect 238812 455892 239404 455920
rect 238812 455880 238818 455892
rect 239398 455880 239404 455892
rect 239456 455880 239462 455932
rect 48222 455472 48228 455524
rect 48280 455512 48286 455524
rect 144178 455512 144184 455524
rect 48280 455484 144184 455512
rect 48280 455472 48286 455484
rect 144178 455472 144184 455484
rect 144236 455472 144242 455524
rect 185578 455472 185584 455524
rect 185636 455512 185642 455524
rect 196066 455512 196072 455524
rect 185636 455484 196072 455512
rect 185636 455472 185642 455484
rect 196066 455472 196072 455484
rect 196124 455472 196130 455524
rect 239398 455472 239404 455524
rect 239456 455512 239462 455524
rect 277486 455512 277492 455524
rect 239456 455484 277492 455512
rect 239456 455472 239462 455484
rect 277486 455472 277492 455484
rect 277544 455472 277550 455524
rect 82722 455404 82728 455456
rect 82780 455444 82786 455456
rect 211154 455444 211160 455456
rect 82780 455416 211160 455444
rect 82780 455404 82786 455416
rect 211154 455404 211160 455416
rect 211212 455404 211218 455456
rect 220078 455404 220084 455456
rect 220136 455444 220142 455456
rect 269758 455444 269764 455456
rect 220136 455416 269764 455444
rect 220136 455404 220142 455416
rect 269758 455404 269764 455416
rect 269816 455404 269822 455456
rect 75178 455336 75184 455388
rect 75236 455376 75242 455388
rect 75822 455376 75828 455388
rect 75236 455348 75828 455376
rect 75236 455336 75242 455348
rect 75822 455336 75828 455348
rect 75880 455376 75886 455388
rect 185578 455376 185584 455388
rect 75880 455348 185584 455376
rect 75880 455336 75886 455348
rect 185578 455336 185584 455348
rect 185636 455336 185642 455388
rect 222562 455064 222568 455116
rect 222620 455104 222626 455116
rect 223482 455104 223488 455116
rect 222620 455076 223488 455104
rect 222620 455064 222626 455076
rect 223482 455064 223488 455076
rect 223540 455064 223546 455116
rect 243538 454656 243544 454708
rect 243596 454696 243602 454708
rect 258074 454696 258080 454708
rect 243596 454668 258080 454696
rect 243596 454656 243602 454668
rect 258074 454656 258080 454668
rect 258132 454696 258138 454708
rect 270862 454696 270868 454708
rect 258132 454668 270868 454696
rect 258132 454656 258138 454668
rect 270862 454656 270868 454668
rect 270920 454656 270926 454708
rect 189074 454112 189080 454164
rect 189132 454152 189138 454164
rect 189132 454124 195974 454152
rect 189132 454112 189138 454124
rect 187050 454044 187056 454096
rect 187108 454084 187114 454096
rect 193582 454084 193588 454096
rect 187108 454056 193588 454084
rect 187108 454044 187114 454056
rect 193582 454044 193588 454056
rect 193640 454044 193646 454096
rect 195946 454084 195974 454124
rect 209774 454084 209780 454096
rect 195946 454056 209780 454084
rect 209774 454044 209780 454056
rect 209832 454084 209838 454096
rect 210418 454084 210424 454096
rect 209832 454056 210424 454084
rect 209832 454044 209838 454056
rect 210418 454044 210424 454056
rect 210476 454044 210482 454096
rect 222562 454044 222568 454096
rect 222620 454084 222626 454096
rect 258074 454084 258080 454096
rect 222620 454056 258080 454084
rect 222620 454044 222626 454056
rect 258074 454044 258080 454056
rect 258132 454044 258138 454096
rect 202138 453976 202144 454028
rect 202196 454016 202202 454028
rect 207014 454016 207020 454028
rect 202196 453988 207020 454016
rect 202196 453976 202202 453988
rect 207014 453976 207020 453988
rect 207072 453976 207078 454028
rect 214558 453976 214564 454028
rect 214616 454016 214622 454028
rect 215938 454016 215944 454028
rect 214616 453988 215944 454016
rect 214616 453976 214622 453988
rect 215938 453976 215944 453988
rect 215996 453976 216002 454028
rect 227806 453976 227812 454028
rect 227864 454016 227870 454028
rect 228726 454016 228732 454028
rect 227864 453988 228732 454016
rect 227864 453976 227870 453988
rect 228726 453976 228732 453988
rect 228784 453976 228790 454028
rect 230750 453976 230756 454028
rect 230808 454016 230814 454028
rect 232590 454016 232596 454028
rect 230808 453988 232596 454016
rect 230808 453976 230814 453988
rect 232590 453976 232596 453988
rect 232648 453976 232654 454028
rect 248598 453976 248604 454028
rect 248656 454016 248662 454028
rect 249702 454016 249708 454028
rect 248656 453988 249708 454016
rect 248656 453976 248662 453988
rect 249702 453976 249708 453988
rect 249760 453976 249766 454028
rect 251542 453976 251548 454028
rect 251600 454016 251606 454028
rect 251910 454016 251916 454028
rect 251600 453988 251916 454016
rect 251600 453976 251606 453988
rect 251910 453976 251916 453988
rect 251968 453976 251974 454028
rect 249058 453908 249064 453960
rect 249116 453948 249122 453960
rect 253382 453948 253388 453960
rect 249116 453920 253388 453948
rect 249116 453908 249122 453920
rect 253382 453908 253388 453920
rect 253440 453908 253446 453960
rect 265710 453296 265716 453348
rect 265768 453336 265774 453348
rect 274910 453336 274916 453348
rect 265768 453308 274916 453336
rect 265768 453296 265774 453308
rect 274910 453296 274916 453308
rect 274968 453296 274974 453348
rect 221182 453160 221188 453212
rect 221240 453200 221246 453212
rect 223666 453200 223672 453212
rect 221240 453172 223672 453200
rect 221240 453160 221246 453172
rect 223666 453160 223672 453172
rect 223724 453160 223730 453212
rect 66070 453024 66076 453076
rect 66128 453064 66134 453076
rect 70486 453064 70492 453076
rect 66128 453036 70492 453064
rect 66128 453024 66134 453036
rect 70486 453024 70492 453036
rect 70544 453024 70550 453076
rect 180058 452684 180064 452736
rect 180116 452724 180122 452736
rect 180610 452724 180616 452736
rect 180116 452696 180616 452724
rect 180116 452684 180122 452696
rect 180610 452684 180616 452696
rect 180668 452724 180674 452736
rect 207934 452724 207940 452736
rect 180668 452696 207940 452724
rect 180668 452684 180674 452696
rect 207934 452684 207940 452696
rect 207992 452684 207998 452736
rect 236454 452684 236460 452736
rect 236512 452724 236518 452736
rect 244274 452724 244280 452736
rect 236512 452696 244280 452724
rect 236512 452684 236518 452696
rect 244274 452684 244280 452696
rect 244332 452684 244338 452736
rect 77662 452616 77668 452668
rect 77720 452656 77726 452668
rect 160830 452656 160836 452668
rect 77720 452628 160836 452656
rect 77720 452616 77726 452628
rect 160830 452616 160836 452628
rect 160888 452656 160894 452668
rect 200206 452656 200212 452668
rect 160888 452628 200212 452656
rect 160888 452616 160894 452628
rect 200206 452616 200212 452628
rect 200264 452616 200270 452668
rect 234430 452616 234436 452668
rect 234488 452656 234494 452668
rect 262398 452656 262404 452668
rect 234488 452628 262404 452656
rect 234488 452616 234494 452628
rect 262398 452616 262404 452628
rect 262456 452616 262462 452668
rect 199286 452548 199292 452600
rect 199344 452588 199350 452600
rect 199470 452588 199476 452600
rect 199344 452560 199476 452588
rect 199344 452548 199350 452560
rect 199470 452548 199476 452560
rect 199528 452548 199534 452600
rect 210510 451868 210516 451920
rect 210568 451908 210574 451920
rect 251082 451908 251088 451920
rect 210568 451880 251088 451908
rect 210568 451868 210574 451880
rect 251082 451868 251088 451880
rect 251140 451868 251146 451920
rect 176470 451324 176476 451376
rect 176528 451364 176534 451376
rect 199286 451364 199292 451376
rect 176528 451336 199292 451364
rect 176528 451324 176534 451336
rect 199286 451324 199292 451336
rect 199344 451324 199350 451376
rect 240134 451324 240140 451376
rect 240192 451364 240198 451376
rect 241422 451364 241428 451376
rect 240192 451336 241428 451364
rect 240192 451324 240198 451336
rect 241422 451324 241428 451336
rect 241480 451364 241486 451376
rect 257338 451364 257344 451376
rect 241480 451336 257344 451364
rect 241480 451324 241486 451336
rect 257338 451324 257344 451336
rect 257396 451324 257402 451376
rect 101398 451256 101404 451308
rect 101456 451296 101462 451308
rect 129090 451296 129096 451308
rect 101456 451268 129096 451296
rect 101456 451256 101462 451268
rect 129090 451256 129096 451268
rect 129148 451296 129154 451308
rect 241054 451296 241060 451308
rect 129148 451268 241060 451296
rect 129148 451256 129154 451268
rect 241054 451256 241060 451268
rect 241112 451256 241118 451308
rect 250622 451256 250628 451308
rect 250680 451296 250686 451308
rect 255222 451296 255228 451308
rect 250680 451268 255228 451296
rect 250680 451256 250686 451268
rect 255222 451256 255228 451268
rect 255280 451256 255286 451308
rect 288526 451256 288532 451308
rect 288584 451296 288590 451308
rect 582650 451296 582656 451308
rect 288584 451268 582656 451296
rect 288584 451256 288590 451268
rect 582650 451256 582656 451268
rect 582708 451256 582714 451308
rect 142154 450684 142160 450696
rect 122806 450656 142160 450684
rect 68922 450576 68928 450628
rect 68980 450616 68986 450628
rect 80054 450616 80060 450628
rect 68980 450588 80060 450616
rect 68980 450576 68986 450588
rect 80054 450576 80060 450588
rect 80112 450576 80118 450628
rect 95142 450576 95148 450628
rect 95200 450616 95206 450628
rect 96706 450616 96712 450628
rect 95200 450588 96712 450616
rect 95200 450576 95206 450588
rect 96706 450576 96712 450588
rect 96764 450576 96770 450628
rect 107930 450576 107936 450628
rect 107988 450616 107994 450628
rect 122806 450616 122834 450656
rect 142154 450644 142160 450656
rect 142212 450684 142218 450696
rect 142982 450684 142988 450696
rect 142212 450656 142988 450684
rect 142212 450644 142218 450656
rect 142982 450644 142988 450656
rect 143040 450644 143046 450696
rect 107988 450588 122834 450616
rect 107988 450576 107994 450588
rect 77294 450508 77300 450560
rect 77352 450548 77358 450560
rect 113818 450548 113824 450560
rect 77352 450520 113824 450548
rect 77352 450508 77358 450520
rect 113818 450508 113824 450520
rect 113876 450508 113882 450560
rect 154390 450508 154396 450560
rect 154448 450548 154454 450560
rect 154448 450520 238754 450548
rect 154448 450508 154454 450520
rect 238726 450480 238754 450520
rect 255222 450508 255228 450560
rect 255280 450548 255286 450560
rect 298278 450548 298284 450560
rect 255280 450520 298284 450548
rect 255280 450508 255286 450520
rect 298278 450508 298284 450520
rect 298336 450508 298342 450560
rect 251174 450480 251180 450492
rect 238726 450452 251180 450480
rect 251174 450440 251180 450452
rect 251232 450480 251238 450492
rect 259638 450480 259644 450492
rect 251232 450452 259644 450480
rect 251232 450440 251238 450452
rect 259638 450440 259644 450452
rect 259696 450440 259702 450492
rect 250438 450236 250444 450288
rect 250496 450276 250502 450288
rect 254118 450276 254124 450288
rect 250496 450248 254124 450276
rect 250496 450236 250502 450248
rect 254118 450236 254124 450248
rect 254176 450236 254182 450288
rect 166442 449896 166448 449948
rect 166500 449936 166506 449948
rect 167638 449936 167644 449948
rect 166500 449908 167644 449936
rect 166500 449896 166506 449908
rect 167638 449896 167644 449908
rect 167696 449896 167702 449948
rect 183370 449896 183376 449948
rect 183428 449936 183434 449948
rect 184934 449936 184940 449948
rect 183428 449908 184940 449936
rect 183428 449896 183434 449908
rect 184934 449896 184940 449908
rect 184992 449896 184998 449948
rect 186222 449896 186228 449948
rect 186280 449936 186286 449948
rect 205634 449936 205640 449948
rect 186280 449908 205640 449936
rect 186280 449896 186286 449908
rect 205634 449896 205640 449908
rect 205692 449896 205698 449948
rect 191926 449692 191932 449744
rect 191984 449732 191990 449744
rect 202322 449732 202328 449744
rect 191984 449704 202328 449732
rect 191984 449692 191990 449704
rect 202322 449692 202328 449704
rect 202380 449692 202386 449744
rect 251818 449692 251824 449744
rect 251876 449732 251882 449744
rect 253934 449732 253940 449744
rect 251876 449704 253940 449732
rect 251876 449692 251882 449704
rect 253934 449692 253940 449704
rect 253992 449692 253998 449744
rect 253474 449556 253480 449608
rect 253532 449596 253538 449608
rect 255682 449596 255688 449608
rect 253532 449568 255688 449596
rect 253532 449556 253538 449568
rect 255682 449556 255688 449568
rect 255740 449556 255746 449608
rect 254578 449216 254584 449268
rect 254636 449256 254642 449268
rect 265066 449256 265072 449268
rect 254636 449228 265072 449256
rect 254636 449216 254642 449228
rect 265066 449216 265072 449228
rect 265124 449216 265130 449268
rect 147766 449148 147772 449200
rect 147824 449188 147830 449200
rect 148870 449188 148876 449200
rect 147824 449160 148876 449188
rect 147824 449148 147830 449160
rect 148870 449148 148876 449160
rect 148928 449188 148934 449200
rect 188338 449188 188344 449200
rect 148928 449160 188344 449188
rect 148928 449148 148934 449160
rect 188338 449148 188344 449160
rect 188396 449148 188402 449200
rect 255590 449148 255596 449200
rect 255648 449188 255654 449200
rect 276014 449188 276020 449200
rect 255648 449160 276020 449188
rect 255648 449148 255654 449160
rect 276014 449148 276020 449160
rect 276072 449148 276078 449200
rect 70854 448604 70860 448656
rect 70912 448644 70918 448656
rect 147766 448644 147772 448656
rect 70912 448616 147772 448644
rect 70912 448604 70918 448616
rect 147766 448604 147772 448616
rect 147824 448604 147830 448656
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 40678 448576 40684 448588
rect 3200 448548 40684 448576
rect 3200 448536 3206 448548
rect 40678 448536 40684 448548
rect 40736 448536 40742 448588
rect 63218 448536 63224 448588
rect 63276 448576 63282 448588
rect 166258 448576 166264 448588
rect 63276 448548 166264 448576
rect 63276 448536 63282 448548
rect 166258 448536 166264 448548
rect 166316 448536 166322 448588
rect 166442 448468 166448 448520
rect 166500 448508 166506 448520
rect 190454 448508 190460 448520
rect 166500 448480 190460 448508
rect 166500 448468 166506 448480
rect 190454 448468 190460 448480
rect 190512 448468 190518 448520
rect 191834 448400 191840 448452
rect 191892 448440 191898 448452
rect 193398 448440 193404 448452
rect 191892 448412 193404 448440
rect 191892 448400 191898 448412
rect 193398 448400 193404 448412
rect 193456 448400 193462 448452
rect 73154 447788 73160 447840
rect 73212 447828 73218 447840
rect 77662 447828 77668 447840
rect 73212 447800 77668 447828
rect 73212 447788 73218 447800
rect 77662 447788 77668 447800
rect 77720 447788 77726 447840
rect 131758 447788 131764 447840
rect 131816 447828 131822 447840
rect 154390 447828 154396 447840
rect 131816 447800 154396 447828
rect 131816 447788 131822 447800
rect 154390 447788 154396 447800
rect 154448 447788 154454 447840
rect 254486 447448 254492 447500
rect 254544 447488 254550 447500
rect 258718 447488 258724 447500
rect 254544 447460 258724 447488
rect 254544 447448 254550 447460
rect 258718 447448 258724 447460
rect 258776 447448 258782 447500
rect 166994 447040 167000 447092
rect 167052 447080 167058 447092
rect 168190 447080 168196 447092
rect 167052 447052 168196 447080
rect 167052 447040 167058 447052
rect 168190 447040 168196 447052
rect 168248 447080 168254 447092
rect 191558 447080 191564 447092
rect 168248 447052 191564 447080
rect 168248 447040 168254 447052
rect 191558 447040 191564 447052
rect 191616 447040 191622 447092
rect 255498 447040 255504 447092
rect 255556 447080 255562 447092
rect 277578 447080 277584 447092
rect 255556 447052 277584 447080
rect 255556 447040 255562 447052
rect 277578 447040 277584 447052
rect 277636 447080 277642 447092
rect 283006 447080 283012 447092
rect 277636 447052 283012 447080
rect 277636 447040 277642 447052
rect 283006 447040 283012 447052
rect 283064 447040 283070 447092
rect 95234 446428 95240 446480
rect 95292 446468 95298 446480
rect 148318 446468 148324 446480
rect 95292 446440 148324 446468
rect 95292 446428 95298 446440
rect 148318 446428 148324 446440
rect 148376 446428 148382 446480
rect 71130 446360 71136 446412
rect 71188 446400 71194 446412
rect 166994 446400 167000 446412
rect 71188 446372 167000 446400
rect 71188 446360 71194 446372
rect 166994 446360 167000 446372
rect 167052 446360 167058 446412
rect 67634 445680 67640 445732
rect 67692 445720 67698 445732
rect 70854 445720 70860 445732
rect 67692 445692 70860 445720
rect 67692 445680 67698 445692
rect 70854 445680 70860 445692
rect 70912 445680 70918 445732
rect 137830 445680 137836 445732
rect 137888 445720 137894 445732
rect 138014 445720 138020 445732
rect 137888 445692 138020 445720
rect 137888 445680 137894 445692
rect 138014 445680 138020 445692
rect 138072 445680 138078 445732
rect 158714 445680 158720 445732
rect 158772 445720 158778 445732
rect 159358 445720 159364 445732
rect 158772 445692 159364 445720
rect 158772 445680 158778 445692
rect 159358 445680 159364 445692
rect 159416 445680 159422 445732
rect 77110 445000 77116 445052
rect 77168 445040 77174 445052
rect 86218 445040 86224 445052
rect 77168 445012 86224 445040
rect 77168 445000 77174 445012
rect 86218 445000 86224 445012
rect 86276 445000 86282 445052
rect 86862 445000 86868 445052
rect 86920 445040 86926 445052
rect 138014 445040 138020 445052
rect 86920 445012 138020 445040
rect 86920 445000 86926 445012
rect 138014 445000 138020 445012
rect 138072 445000 138078 445052
rect 153010 445000 153016 445052
rect 153068 445040 153074 445052
rect 190362 445040 190368 445052
rect 153068 445012 190368 445040
rect 153068 445000 153074 445012
rect 190362 445000 190368 445012
rect 190420 445040 190426 445052
rect 191558 445040 191564 445052
rect 190420 445012 191564 445040
rect 190420 445000 190426 445012
rect 191558 445000 191564 445012
rect 191616 445000 191622 445052
rect 83458 444456 83464 444508
rect 83516 444496 83522 444508
rect 86862 444496 86868 444508
rect 83516 444468 86868 444496
rect 83516 444456 83522 444468
rect 86862 444456 86868 444468
rect 86920 444456 86926 444508
rect 101398 444456 101404 444508
rect 101456 444496 101462 444508
rect 104158 444496 104164 444508
rect 101456 444468 104164 444496
rect 101456 444456 101462 444468
rect 104158 444456 104164 444468
rect 104216 444456 104222 444508
rect 70394 444388 70400 444440
rect 70452 444428 70458 444440
rect 158714 444428 158720 444440
rect 70452 444400 158720 444428
rect 70452 444388 70458 444400
rect 158714 444388 158720 444400
rect 158772 444388 158778 444440
rect 173158 444320 173164 444372
rect 173216 444360 173222 444372
rect 180058 444360 180064 444372
rect 173216 444332 180064 444360
rect 173216 444320 173222 444332
rect 180058 444320 180064 444332
rect 180116 444320 180122 444372
rect 255498 443640 255504 443692
rect 255556 443680 255562 443692
rect 260558 443680 260564 443692
rect 255556 443652 260564 443680
rect 255556 443640 255562 443652
rect 260558 443640 260564 443652
rect 260616 443640 260622 443692
rect 78674 443028 78680 443080
rect 78732 443068 78738 443080
rect 173158 443068 173164 443080
rect 78732 443040 173164 443068
rect 78732 443028 78738 443040
rect 173158 443028 173164 443040
rect 173216 443028 173222 443080
rect 66162 442960 66168 443012
rect 66220 443000 66226 443012
rect 193030 443000 193036 443012
rect 66220 442972 193036 443000
rect 66220 442960 66226 442972
rect 193030 442960 193036 442972
rect 193088 442960 193094 443012
rect 270586 443000 270592 443012
rect 269316 442972 270592 443000
rect 269316 442944 269344 442972
rect 270586 442960 270592 442972
rect 270644 442960 270650 443012
rect 77202 442892 77208 442944
rect 77260 442932 77266 442944
rect 83182 442932 83188 442944
rect 77260 442904 83188 442932
rect 77260 442892 77266 442904
rect 83182 442892 83188 442904
rect 83240 442892 83246 442944
rect 184750 442892 184756 442944
rect 184808 442932 184814 442944
rect 184934 442932 184940 442944
rect 184808 442904 184940 442932
rect 184808 442892 184814 442904
rect 184934 442892 184940 442904
rect 184992 442892 184998 442944
rect 269298 442892 269304 442944
rect 269356 442892 269362 442944
rect 262858 442280 262864 442332
rect 262916 442320 262922 442332
rect 272058 442320 272064 442332
rect 262916 442292 272064 442320
rect 262916 442280 262922 442292
rect 272058 442280 272064 442292
rect 272116 442280 272122 442332
rect 260558 442212 260564 442264
rect 260616 442252 260622 442264
rect 269298 442252 269304 442264
rect 260616 442224 269304 442252
rect 260616 442212 260622 442224
rect 269298 442212 269304 442224
rect 269356 442212 269362 442264
rect 88242 441668 88248 441720
rect 88300 441708 88306 441720
rect 184198 441708 184204 441720
rect 88300 441680 184204 441708
rect 88300 441668 88306 441680
rect 184198 441668 184204 441680
rect 184256 441668 184262 441720
rect 67726 441600 67732 441652
rect 67784 441640 67790 441652
rect 184750 441640 184756 441652
rect 67784 441612 184756 441640
rect 67784 441600 67790 441612
rect 184750 441600 184756 441612
rect 184808 441640 184814 441652
rect 191374 441640 191380 441652
rect 184808 441612 191380 441640
rect 184808 441600 184814 441612
rect 191374 441600 191380 441612
rect 191432 441600 191438 441652
rect 64690 440852 64696 440904
rect 64748 440892 64754 440904
rect 186038 440892 186044 440904
rect 64748 440864 186044 440892
rect 64748 440852 64754 440864
rect 186038 440852 186044 440864
rect 186096 440892 186102 440904
rect 190638 440892 190644 440904
rect 186096 440864 190644 440892
rect 186096 440852 186102 440864
rect 190638 440852 190644 440864
rect 190696 440852 190702 440904
rect 78582 440240 78588 440292
rect 78640 440280 78646 440292
rect 174538 440280 174544 440292
rect 78640 440252 174544 440280
rect 78640 440240 78646 440252
rect 174538 440240 174544 440252
rect 174596 440240 174602 440292
rect 155678 440172 155684 440224
rect 155736 440212 155742 440224
rect 191650 440212 191656 440224
rect 155736 440184 191656 440212
rect 155736 440172 155742 440184
rect 191650 440172 191656 440184
rect 191708 440172 191714 440224
rect 4798 439492 4804 439544
rect 4856 439532 4862 439544
rect 103790 439532 103796 439544
rect 4856 439504 103796 439532
rect 4856 439492 4862 439504
rect 103790 439492 103796 439504
rect 103848 439492 103854 439544
rect 177942 439492 177948 439544
rect 178000 439532 178006 439544
rect 185578 439532 185584 439544
rect 178000 439504 185584 439532
rect 178000 439492 178006 439504
rect 185578 439492 185584 439504
rect 185636 439492 185642 439544
rect 255498 439492 255504 439544
rect 255556 439532 255562 439544
rect 288618 439532 288624 439544
rect 255556 439504 288624 439532
rect 255556 439492 255562 439504
rect 288618 439492 288624 439504
rect 288676 439492 288682 439544
rect 104802 438948 104808 439000
rect 104860 438988 104866 439000
rect 107654 438988 107660 439000
rect 104860 438960 107660 438988
rect 104860 438948 104866 438960
rect 107654 438948 107660 438960
rect 107712 438948 107718 439000
rect 67358 438880 67364 438932
rect 67416 438920 67422 438932
rect 154022 438920 154028 438932
rect 67416 438892 154028 438920
rect 67416 438880 67422 438892
rect 154022 438880 154028 438892
rect 154080 438880 154086 438932
rect 103790 438812 103796 438864
rect 103848 438852 103854 438864
rect 104434 438852 104440 438864
rect 103848 438824 104440 438852
rect 103848 438812 103854 438824
rect 104434 438812 104440 438824
rect 104492 438852 104498 438864
rect 106918 438852 106924 438864
rect 104492 438824 106924 438852
rect 104492 438812 104498 438824
rect 106918 438812 106924 438824
rect 106976 438812 106982 438864
rect 178034 438132 178040 438184
rect 178092 438172 178098 438184
rect 179230 438172 179236 438184
rect 178092 438144 179236 438172
rect 178092 438132 178098 438144
rect 179230 438132 179236 438144
rect 179288 438172 179294 438184
rect 190638 438172 190644 438184
rect 179288 438144 190644 438172
rect 179288 438132 179294 438144
rect 190638 438132 190644 438144
rect 190696 438132 190702 438184
rect 255498 438132 255504 438184
rect 255556 438172 255562 438184
rect 281626 438172 281632 438184
rect 255556 438144 281632 438172
rect 255556 438132 255562 438144
rect 281626 438132 281632 438144
rect 281684 438132 281690 438184
rect 67266 437452 67272 437504
rect 67324 437492 67330 437504
rect 67542 437492 67548 437504
rect 67324 437464 67548 437492
rect 67324 437452 67330 437464
rect 67542 437452 67548 437464
rect 67600 437492 67606 437504
rect 147030 437492 147036 437504
rect 67600 437464 147036 437492
rect 67600 437452 67606 437464
rect 147030 437452 147036 437464
rect 147088 437452 147094 437504
rect 255498 437452 255504 437504
rect 255556 437492 255562 437504
rect 296806 437492 296812 437504
rect 255556 437464 296812 437492
rect 255556 437452 255562 437464
rect 296806 437452 296812 437464
rect 296864 437452 296870 437504
rect 102502 436772 102508 436824
rect 102560 436812 102566 436824
rect 111058 436812 111064 436824
rect 102560 436784 111064 436812
rect 102560 436772 102566 436784
rect 111058 436772 111064 436784
rect 111116 436772 111122 436824
rect 177942 436772 177948 436824
rect 178000 436812 178006 436824
rect 184658 436812 184664 436824
rect 178000 436784 184664 436812
rect 178000 436772 178006 436784
rect 184658 436772 184664 436784
rect 184716 436812 184722 436824
rect 191650 436812 191656 436824
rect 184716 436784 191656 436812
rect 184716 436772 184722 436784
rect 191650 436772 191656 436784
rect 191708 436772 191714 436824
rect 110782 436704 110788 436756
rect 110840 436744 110846 436756
rect 186314 436744 186320 436756
rect 110840 436716 186320 436744
rect 110840 436704 110846 436716
rect 186314 436704 186320 436716
rect 186372 436704 186378 436756
rect 255682 436704 255688 436756
rect 255740 436744 255746 436756
rect 285950 436744 285956 436756
rect 255740 436716 285956 436744
rect 255740 436704 255746 436716
rect 285950 436704 285956 436716
rect 286008 436704 286014 436756
rect 94038 436636 94044 436688
rect 94096 436676 94102 436688
rect 98638 436676 98644 436688
rect 94096 436648 98644 436676
rect 94096 436636 94102 436648
rect 98638 436636 98644 436648
rect 98696 436636 98702 436688
rect 78214 436364 78220 436416
rect 78272 436404 78278 436416
rect 79318 436404 79324 436416
rect 78272 436376 79324 436404
rect 78272 436364 78278 436376
rect 79318 436364 79324 436376
rect 79376 436364 79382 436416
rect 59262 436160 59268 436212
rect 59320 436200 59326 436212
rect 69658 436200 69664 436212
rect 59320 436172 69664 436200
rect 59320 436160 59326 436172
rect 69658 436160 69664 436172
rect 69716 436200 69722 436212
rect 70026 436200 70032 436212
rect 69716 436172 70032 436200
rect 69716 436160 69722 436172
rect 70026 436160 70032 436172
rect 70084 436160 70090 436212
rect 81158 436160 81164 436212
rect 81216 436200 81222 436212
rect 88978 436200 88984 436212
rect 81216 436172 88984 436200
rect 81216 436160 81222 436172
rect 88978 436160 88984 436172
rect 89036 436160 89042 436212
rect 15838 436092 15844 436144
rect 15896 436132 15902 436144
rect 70854 436132 70860 436144
rect 15896 436104 70860 436132
rect 15896 436092 15902 436104
rect 70854 436092 70860 436104
rect 70912 436132 70918 436144
rect 75178 436132 75184 436144
rect 70912 436104 75184 436132
rect 70912 436092 70918 436104
rect 75178 436092 75184 436104
rect 75236 436092 75242 436144
rect 87322 436092 87328 436144
rect 87380 436132 87386 436144
rect 88242 436132 88248 436144
rect 87380 436104 88248 436132
rect 87380 436092 87386 436104
rect 88242 436092 88248 436104
rect 88300 436092 88306 436144
rect 148318 435344 148324 435396
rect 148376 435384 148382 435396
rect 185670 435384 185676 435396
rect 148376 435356 185676 435384
rect 148376 435344 148382 435356
rect 185670 435344 185676 435356
rect 185728 435344 185734 435396
rect 255498 435344 255504 435396
rect 255556 435384 255562 435396
rect 259730 435384 259736 435396
rect 255556 435356 259736 435384
rect 255556 435344 255562 435356
rect 259730 435344 259736 435356
rect 259788 435384 259794 435396
rect 276290 435384 276296 435396
rect 259788 435356 276296 435384
rect 259788 435344 259794 435356
rect 276290 435344 276296 435356
rect 276348 435344 276354 435396
rect 65886 434800 65892 434852
rect 65944 434840 65950 434852
rect 158806 434840 158812 434852
rect 65944 434812 158812 434840
rect 65944 434800 65950 434812
rect 158806 434800 158812 434812
rect 158864 434800 158870 434852
rect 3418 434732 3424 434784
rect 3476 434772 3482 434784
rect 112438 434772 112444 434784
rect 3476 434744 112444 434772
rect 3476 434732 3482 434744
rect 112438 434732 112444 434744
rect 112496 434732 112502 434784
rect 272518 434772 272524 434784
rect 272431 434744 272524 434772
rect 272518 434732 272524 434744
rect 272576 434772 272582 434784
rect 295518 434772 295524 434784
rect 272576 434744 295524 434772
rect 272576 434732 272582 434744
rect 295518 434732 295524 434744
rect 295576 434732 295582 434784
rect 67542 434664 67548 434716
rect 67600 434704 67606 434716
rect 71314 434704 71320 434716
rect 67600 434676 71320 434704
rect 67600 434664 67606 434676
rect 71314 434664 71320 434676
rect 71372 434664 71378 434716
rect 115750 434664 115756 434716
rect 115808 434704 115814 434716
rect 146938 434704 146944 434716
rect 115808 434676 146944 434704
rect 115808 434664 115814 434676
rect 146938 434664 146944 434676
rect 146996 434664 147002 434716
rect 187050 434664 187056 434716
rect 187108 434704 187114 434716
rect 189074 434704 189080 434716
rect 187108 434676 189080 434704
rect 187108 434664 187114 434676
rect 189074 434664 189080 434676
rect 189132 434664 189138 434716
rect 255498 434664 255504 434716
rect 255556 434704 255562 434716
rect 272536 434704 272564 434732
rect 255556 434676 272564 434704
rect 255556 434664 255562 434676
rect 68646 434052 68652 434104
rect 68704 434092 68710 434104
rect 71774 434092 71780 434104
rect 68704 434064 71780 434092
rect 68704 434052 68710 434064
rect 71774 434052 71780 434064
rect 71832 434092 71838 434104
rect 72694 434092 72700 434104
rect 71832 434064 72700 434092
rect 71832 434052 71838 434064
rect 72694 434052 72700 434064
rect 72752 434052 72758 434104
rect 53742 433984 53748 434036
rect 53800 434024 53806 434036
rect 61746 434024 61752 434036
rect 53800 433996 61752 434024
rect 53800 433984 53806 433996
rect 61746 433984 61752 433996
rect 61804 434024 61810 434036
rect 66806 434024 66812 434036
rect 61804 433996 66812 434024
rect 61804 433984 61810 433996
rect 66806 433984 66812 433996
rect 66864 433984 66870 434036
rect 72602 433984 72608 434036
rect 72660 434024 72666 434036
rect 132494 434024 132500 434036
rect 72660 433996 132500 434024
rect 72660 433984 72666 433996
rect 132494 433984 132500 433996
rect 132552 433984 132558 434036
rect 73982 433644 73988 433696
rect 74040 433644 74046 433696
rect 74000 433276 74028 433644
rect 64846 433248 74028 433276
rect 52362 432624 52368 432676
rect 52420 432664 52426 432676
rect 64846 432664 64874 433248
rect 115842 433236 115848 433288
rect 115900 433276 115906 433288
rect 115900 433248 142154 433276
rect 115900 433236 115906 433248
rect 142126 433208 142154 433248
rect 150250 433236 150256 433288
rect 150308 433276 150314 433288
rect 150526 433276 150532 433288
rect 150308 433248 150532 433276
rect 150308 433236 150314 433248
rect 150526 433236 150532 433248
rect 150584 433236 150590 433288
rect 151078 433208 151084 433220
rect 142126 433180 151084 433208
rect 151078 433168 151084 433180
rect 151136 433168 151142 433220
rect 52420 432636 64874 432664
rect 52420 432624 52426 432636
rect 255958 432624 255964 432676
rect 256016 432664 256022 432676
rect 256878 432664 256884 432676
rect 256016 432636 256884 432664
rect 256016 432624 256022 432636
rect 256878 432624 256884 432636
rect 256936 432664 256942 432676
rect 266630 432664 266636 432676
rect 256936 432636 266636 432664
rect 256936 432624 256942 432636
rect 266630 432624 266636 432636
rect 266688 432624 266694 432676
rect 53650 432556 53656 432608
rect 53708 432596 53714 432608
rect 145650 432596 145656 432608
rect 53708 432568 145656 432596
rect 53708 432556 53714 432568
rect 145650 432556 145656 432568
rect 145708 432556 145714 432608
rect 258718 432556 258724 432608
rect 258776 432596 258782 432608
rect 271966 432596 271972 432608
rect 258776 432568 271972 432596
rect 258776 432556 258782 432568
rect 271966 432556 271972 432568
rect 272024 432556 272030 432608
rect 191650 431984 191656 431996
rect 178512 431956 191656 431984
rect 115566 431876 115572 431928
rect 115624 431916 115630 431928
rect 126238 431916 126244 431928
rect 115624 431888 126244 431916
rect 115624 431876 115630 431888
rect 126238 431876 126244 431888
rect 126296 431876 126302 431928
rect 155770 431876 155776 431928
rect 155828 431916 155834 431928
rect 178034 431916 178040 431928
rect 155828 431888 178040 431916
rect 155828 431876 155834 431888
rect 178034 431876 178040 431888
rect 178092 431916 178098 431928
rect 178512 431916 178540 431956
rect 191650 431944 191656 431956
rect 191708 431944 191714 431996
rect 178092 431888 178540 431916
rect 178092 431876 178098 431888
rect 112898 431196 112904 431248
rect 112956 431236 112962 431248
rect 124858 431236 124864 431248
rect 112956 431208 124864 431236
rect 112956 431196 112962 431208
rect 124858 431196 124864 431208
rect 124916 431196 124922 431248
rect 154022 431196 154028 431248
rect 154080 431236 154086 431248
rect 170490 431236 170496 431248
rect 154080 431208 170496 431236
rect 154080 431196 154086 431208
rect 170490 431196 170496 431208
rect 170548 431236 170554 431248
rect 191742 431236 191748 431248
rect 170548 431208 191748 431236
rect 170548 431196 170554 431208
rect 191742 431196 191748 431208
rect 191800 431196 191806 431248
rect 255406 431196 255412 431248
rect 255464 431236 255470 431248
rect 289906 431236 289912 431248
rect 255464 431208 289912 431236
rect 255464 431196 255470 431208
rect 289906 431196 289912 431208
rect 289964 431196 289970 431248
rect 65794 430652 65800 430704
rect 65852 430692 65858 430704
rect 66070 430692 66076 430704
rect 65852 430664 66076 430692
rect 65852 430652 65858 430664
rect 66070 430652 66076 430664
rect 66128 430652 66134 430704
rect 63310 430584 63316 430636
rect 63368 430624 63374 430636
rect 67542 430624 67548 430636
rect 63368 430596 67548 430624
rect 63368 430584 63374 430596
rect 67542 430584 67548 430596
rect 67600 430584 67606 430636
rect 115750 430516 115756 430568
rect 115808 430556 115814 430568
rect 133230 430556 133236 430568
rect 115808 430528 133236 430556
rect 115808 430516 115814 430528
rect 133230 430516 133236 430528
rect 133288 430516 133294 430568
rect 166350 430516 166356 430568
rect 166408 430556 166414 430568
rect 191006 430556 191012 430568
rect 166408 430528 191012 430556
rect 166408 430516 166414 430528
rect 191006 430516 191012 430528
rect 191064 430516 191070 430568
rect 139302 429836 139308 429888
rect 139360 429876 139366 429888
rect 155310 429876 155316 429888
rect 139360 429848 155316 429876
rect 139360 429836 139366 429848
rect 155310 429836 155316 429848
rect 155368 429836 155374 429888
rect 60550 429224 60556 429276
rect 60608 429264 60614 429276
rect 66070 429264 66076 429276
rect 60608 429236 66076 429264
rect 60608 429224 60614 429236
rect 66070 429224 66076 429236
rect 66128 429264 66134 429276
rect 66622 429264 66628 429276
rect 66128 429236 66628 429264
rect 66128 429224 66134 429236
rect 66622 429224 66628 429236
rect 66680 429224 66686 429276
rect 115842 429088 115848 429140
rect 115900 429128 115906 429140
rect 151262 429128 151268 429140
rect 115900 429100 151268 429128
rect 115900 429088 115906 429100
rect 151262 429088 151268 429100
rect 151320 429088 151326 429140
rect 152918 429088 152924 429140
rect 152976 429128 152982 429140
rect 190822 429128 190828 429140
rect 152976 429100 190828 429128
rect 152976 429088 152982 429100
rect 190822 429088 190828 429100
rect 190880 429088 190886 429140
rect 176654 427728 176660 427780
rect 176712 427768 176718 427780
rect 190822 427768 190828 427780
rect 176712 427740 190828 427768
rect 176712 427728 176718 427740
rect 190822 427728 190828 427740
rect 190880 427728 190886 427780
rect 119338 427048 119344 427100
rect 119396 427088 119402 427100
rect 133138 427088 133144 427100
rect 119396 427060 133144 427088
rect 119396 427048 119402 427060
rect 133138 427048 133144 427060
rect 133196 427048 133202 427100
rect 151630 427048 151636 427100
rect 151688 427088 151694 427100
rect 176654 427088 176660 427100
rect 151688 427060 176660 427088
rect 151688 427048 151694 427060
rect 176654 427048 176660 427060
rect 176712 427048 176718 427100
rect 285766 427048 285772 427100
rect 285824 427088 285830 427100
rect 291286 427088 291292 427100
rect 285824 427060 291292 427088
rect 285824 427048 285830 427060
rect 291286 427048 291292 427060
rect 291344 427088 291350 427100
rect 582558 427088 582564 427100
rect 291344 427060 582564 427088
rect 291344 427048 291350 427060
rect 582558 427048 582564 427060
rect 582616 427048 582622 427100
rect 64690 426436 64696 426488
rect 64748 426476 64754 426488
rect 66806 426476 66812 426488
rect 64748 426448 66812 426476
rect 64748 426436 64754 426448
rect 66806 426436 66812 426448
rect 66864 426436 66870 426488
rect 255406 426436 255412 426488
rect 255464 426476 255470 426488
rect 285766 426476 285772 426488
rect 255464 426448 285772 426476
rect 255464 426436 255470 426448
rect 285766 426436 285772 426448
rect 285824 426436 285830 426488
rect 115842 426368 115848 426420
rect 115900 426408 115906 426420
rect 124214 426408 124220 426420
rect 115900 426380 124220 426408
rect 115900 426368 115906 426380
rect 124214 426368 124220 426380
rect 124272 426368 124278 426420
rect 255498 426368 255504 426420
rect 255556 426408 255562 426420
rect 273530 426408 273536 426420
rect 255556 426380 273536 426408
rect 255556 426368 255562 426380
rect 273530 426368 273536 426380
rect 273588 426368 273594 426420
rect 41322 425688 41328 425740
rect 41380 425728 41386 425740
rect 65794 425728 65800 425740
rect 41380 425700 65800 425728
rect 41380 425688 41386 425700
rect 65794 425688 65800 425700
rect 65852 425728 65858 425740
rect 66622 425728 66628 425740
rect 65852 425700 66628 425728
rect 65852 425688 65858 425700
rect 66622 425688 66628 425700
rect 66680 425688 66686 425740
rect 173802 425688 173808 425740
rect 173860 425728 173866 425740
rect 191742 425728 191748 425740
rect 173860 425700 191748 425728
rect 173860 425688 173866 425700
rect 191742 425688 191748 425700
rect 191800 425688 191806 425740
rect 273530 425688 273536 425740
rect 273588 425728 273594 425740
rect 283190 425728 283196 425740
rect 273588 425700 283196 425728
rect 273588 425688 273594 425700
rect 283190 425688 283196 425700
rect 283248 425688 283254 425740
rect 115842 425008 115848 425060
rect 115900 425048 115906 425060
rect 155218 425048 155224 425060
rect 115900 425020 155224 425048
rect 115900 425008 115906 425020
rect 155218 425008 155224 425020
rect 155276 425008 155282 425060
rect 175182 424328 175188 424380
rect 175240 424368 175246 424380
rect 186130 424368 186136 424380
rect 175240 424340 186136 424368
rect 175240 424328 175246 424340
rect 186130 424328 186136 424340
rect 186188 424368 186194 424380
rect 191742 424368 191748 424380
rect 186188 424340 191748 424368
rect 186188 424328 186194 424340
rect 191742 424328 191748 424340
rect 191800 424328 191806 424380
rect 53742 423648 53748 423700
rect 53800 423688 53806 423700
rect 66806 423688 66812 423700
rect 53800 423660 66812 423688
rect 53800 423648 53806 423660
rect 66806 423648 66812 423660
rect 66864 423648 66870 423700
rect 115842 423580 115848 423632
rect 115900 423620 115906 423632
rect 118694 423620 118700 423632
rect 115900 423592 118700 423620
rect 115900 423580 115906 423592
rect 118694 423580 118700 423592
rect 118752 423620 118758 423632
rect 148318 423620 148324 423632
rect 118752 423592 148324 423620
rect 118752 423580 118758 423592
rect 148318 423580 148324 423592
rect 148376 423580 148382 423632
rect 155862 423580 155868 423632
rect 155920 423620 155926 423632
rect 158806 423620 158812 423632
rect 155920 423592 158812 423620
rect 155920 423580 155926 423592
rect 158806 423580 158812 423592
rect 158864 423620 158870 423632
rect 191006 423620 191012 423632
rect 158864 423592 191012 423620
rect 158864 423580 158870 423592
rect 191006 423580 191012 423592
rect 191064 423580 191070 423632
rect 50982 422288 50988 422340
rect 51040 422328 51046 422340
rect 66254 422328 66260 422340
rect 51040 422300 66260 422328
rect 51040 422288 51046 422300
rect 66254 422288 66260 422300
rect 66312 422288 66318 422340
rect 255498 422288 255504 422340
rect 255556 422328 255562 422340
rect 281810 422328 281816 422340
rect 255556 422300 281816 422328
rect 255556 422288 255562 422300
rect 281810 422288 281816 422300
rect 281868 422288 281874 422340
rect 64598 421064 64604 421116
rect 64656 421104 64662 421116
rect 67174 421104 67180 421116
rect 64656 421076 67180 421104
rect 64656 421064 64662 421076
rect 67174 421064 67180 421076
rect 67232 421064 67238 421116
rect 48130 420928 48136 420980
rect 48188 420968 48194 420980
rect 66898 420968 66904 420980
rect 48188 420940 66904 420968
rect 48188 420928 48194 420940
rect 66898 420928 66904 420940
rect 66956 420928 66962 420980
rect 143442 420928 143448 420980
rect 143500 420968 143506 420980
rect 192478 420968 192484 420980
rect 143500 420940 192484 420968
rect 143500 420928 143506 420940
rect 192478 420928 192484 420940
rect 192536 420928 192542 420980
rect 255498 420928 255504 420980
rect 255556 420968 255562 420980
rect 298370 420968 298376 420980
rect 255556 420940 298376 420968
rect 255556 420928 255562 420940
rect 298370 420928 298376 420940
rect 298428 420928 298434 420980
rect 155586 420860 155592 420912
rect 155644 420900 155650 420912
rect 191742 420900 191748 420912
rect 155644 420872 191748 420900
rect 155644 420860 155650 420872
rect 191742 420860 191748 420872
rect 191800 420860 191806 420912
rect 263778 420180 263784 420232
rect 263836 420220 263842 420232
rect 264882 420220 264888 420232
rect 263836 420192 264888 420220
rect 263836 420180 263842 420192
rect 264882 420180 264888 420192
rect 264940 420220 264946 420232
rect 298094 420220 298100 420232
rect 264940 420192 298100 420220
rect 264940 420180 264946 420192
rect 298094 420180 298100 420192
rect 298152 420180 298158 420232
rect 255498 419500 255504 419552
rect 255556 419540 255562 419552
rect 263778 419540 263784 419552
rect 255556 419512 263784 419540
rect 255556 419500 255562 419512
rect 263778 419500 263784 419512
rect 263836 419500 263842 419552
rect 149790 419432 149796 419484
rect 149848 419472 149854 419484
rect 191742 419472 191748 419484
rect 149848 419444 191748 419472
rect 149848 419432 149854 419444
rect 191742 419432 191748 419444
rect 191800 419432 191806 419484
rect 255406 419432 255412 419484
rect 255464 419472 255470 419484
rect 285674 419472 285680 419484
rect 255464 419444 285680 419472
rect 255464 419432 255470 419444
rect 285674 419432 285680 419444
rect 285732 419472 285738 419484
rect 287422 419472 287428 419484
rect 285732 419444 287428 419472
rect 285732 419432 285738 419444
rect 287422 419432 287428 419444
rect 287480 419472 287486 419484
rect 582374 419472 582380 419484
rect 287480 419444 582380 419472
rect 287480 419432 287486 419444
rect 582374 419432 582380 419444
rect 582432 419432 582438 419484
rect 115842 419364 115848 419416
rect 115900 419404 115906 419416
rect 153838 419404 153844 419416
rect 115900 419376 153844 419404
rect 115900 419364 115906 419376
rect 153838 419364 153844 419376
rect 153896 419364 153902 419416
rect 176562 418752 176568 418804
rect 176620 418792 176626 418804
rect 187694 418792 187700 418804
rect 176620 418764 187700 418792
rect 176620 418752 176626 418764
rect 187694 418752 187700 418764
rect 187752 418752 187758 418804
rect 61654 418208 61660 418260
rect 61712 418248 61718 418260
rect 63218 418248 63224 418260
rect 61712 418220 63224 418248
rect 61712 418208 61718 418220
rect 63218 418208 63224 418220
rect 63276 418248 63282 418260
rect 66622 418248 66628 418260
rect 63276 418220 66628 418248
rect 63276 418208 63282 418220
rect 66622 418208 66628 418220
rect 66680 418208 66686 418260
rect 61930 418072 61936 418124
rect 61988 418112 61994 418124
rect 66990 418112 66996 418124
rect 61988 418084 66996 418112
rect 61988 418072 61994 418084
rect 66990 418072 66996 418084
rect 67048 418072 67054 418124
rect 281442 418072 281448 418124
rect 281500 418112 281506 418124
rect 582466 418112 582472 418124
rect 281500 418084 582472 418112
rect 281500 418072 281506 418084
rect 582466 418072 582472 418084
rect 582524 418072 582530 418124
rect 148870 417392 148876 417444
rect 148928 417432 148934 417444
rect 166350 417432 166356 417444
rect 148928 417404 166356 417432
rect 148928 417392 148934 417404
rect 166350 417392 166356 417404
rect 166408 417392 166414 417444
rect 255406 417392 255412 417444
rect 255464 417432 255470 417444
rect 280430 417432 280436 417444
rect 255464 417404 280436 417432
rect 255464 417392 255470 417404
rect 280430 417392 280436 417404
rect 280488 417432 280494 417444
rect 281442 417432 281448 417444
rect 280488 417404 281448 417432
rect 280488 417392 280494 417404
rect 281442 417392 281448 417404
rect 281500 417392 281506 417444
rect 118694 417188 118700 417240
rect 118752 417228 118758 417240
rect 119338 417228 119344 417240
rect 118752 417200 119344 417228
rect 118752 417188 118758 417200
rect 119338 417188 119344 417200
rect 119396 417188 119402 417240
rect 115842 416780 115848 416832
rect 115900 416820 115906 416832
rect 118694 416820 118700 416832
rect 115900 416792 118700 416820
rect 115900 416780 115906 416792
rect 118694 416780 118700 416792
rect 118752 416780 118758 416832
rect 126238 416780 126244 416832
rect 126296 416820 126302 416832
rect 154390 416820 154396 416832
rect 126296 416792 154396 416820
rect 126296 416780 126302 416792
rect 154390 416780 154396 416792
rect 154448 416780 154454 416832
rect 166350 416780 166356 416832
rect 166408 416820 166414 416832
rect 166718 416820 166724 416832
rect 166408 416792 166724 416820
rect 166408 416780 166414 416792
rect 166718 416780 166724 416792
rect 166776 416820 166782 416832
rect 191742 416820 191748 416832
rect 166776 416792 191748 416820
rect 166776 416780 166782 416792
rect 191742 416780 191748 416792
rect 191800 416780 191806 416832
rect 255406 416780 255412 416832
rect 255464 416820 255470 416832
rect 265158 416820 265164 416832
rect 255464 416792 265164 416820
rect 255464 416780 255470 416792
rect 265158 416780 265164 416792
rect 265216 416780 265222 416832
rect 149054 416100 149060 416152
rect 149112 416140 149118 416152
rect 150250 416140 150256 416152
rect 149112 416112 150256 416140
rect 149112 416100 149118 416112
rect 150250 416100 150256 416112
rect 150308 416140 150314 416152
rect 169754 416140 169760 416152
rect 150308 416112 169760 416140
rect 150308 416100 150314 416112
rect 169754 416100 169760 416112
rect 169812 416100 169818 416152
rect 50890 416032 50896 416084
rect 50948 416072 50954 416084
rect 56410 416072 56416 416084
rect 50948 416044 56416 416072
rect 50948 416032 50954 416044
rect 56410 416032 56416 416044
rect 56468 416072 56474 416084
rect 66806 416072 66812 416084
rect 56468 416044 66812 416072
rect 56468 416032 56474 416044
rect 66806 416032 66812 416044
rect 66864 416032 66870 416084
rect 120074 416032 120080 416084
rect 120132 416072 120138 416084
rect 151170 416072 151176 416084
rect 120132 416044 151176 416072
rect 120132 416032 120138 416044
rect 151170 416032 151176 416044
rect 151228 416032 151234 416084
rect 153102 416032 153108 416084
rect 153160 416072 153166 416084
rect 190638 416072 190644 416084
rect 153160 416044 190644 416072
rect 153160 416032 153166 416044
rect 190638 416032 190644 416044
rect 190696 416032 190702 416084
rect 115842 415420 115848 415472
rect 115900 415460 115906 415472
rect 120074 415460 120080 415472
rect 115900 415432 120080 415460
rect 115900 415420 115906 415432
rect 120074 415420 120080 415432
rect 120132 415420 120138 415472
rect 122190 415420 122196 415472
rect 122248 415460 122254 415472
rect 149054 415460 149060 415472
rect 122248 415432 149060 415460
rect 122248 415420 122254 415432
rect 149054 415420 149060 415432
rect 149112 415420 149118 415472
rect 144178 415352 144184 415404
rect 144236 415392 144242 415404
rect 191466 415392 191472 415404
rect 144236 415364 191472 415392
rect 144236 415352 144242 415364
rect 191466 415352 191472 415364
rect 191524 415352 191530 415404
rect 184842 415284 184848 415336
rect 184900 415324 184906 415336
rect 188338 415324 188344 415336
rect 184900 415296 188344 415324
rect 184900 415284 184906 415296
rect 188338 415284 188344 415296
rect 188396 415284 188402 415336
rect 115842 414672 115848 414724
rect 115900 414712 115906 414724
rect 122742 414712 122748 414724
rect 115900 414684 122748 414712
rect 115900 414672 115906 414684
rect 122742 414672 122748 414684
rect 122800 414712 122806 414724
rect 125686 414712 125692 414724
rect 122800 414684 125692 414712
rect 122800 414672 122806 414684
rect 125686 414672 125692 414684
rect 125744 414672 125750 414724
rect 55030 413992 55036 414044
rect 55088 414032 55094 414044
rect 66806 414032 66812 414044
rect 55088 414004 66812 414032
rect 55088 413992 55094 414004
rect 66806 413992 66812 414004
rect 66864 413992 66870 414044
rect 115750 413924 115756 413976
rect 115808 413964 115814 413976
rect 127618 413964 127624 413976
rect 115808 413936 127624 413964
rect 115808 413924 115814 413936
rect 127618 413924 127624 413936
rect 127676 413924 127682 413976
rect 255406 413788 255412 413840
rect 255464 413828 255470 413840
rect 259638 413828 259644 413840
rect 255464 413800 259644 413828
rect 255464 413788 255470 413800
rect 259638 413788 259644 413800
rect 259696 413788 259702 413840
rect 114738 413584 114744 413636
rect 114796 413624 114802 413636
rect 117314 413624 117320 413636
rect 114796 413596 117320 413624
rect 114796 413584 114802 413596
rect 117314 413584 117320 413596
rect 117372 413584 117378 413636
rect 55122 413244 55128 413296
rect 55180 413284 55186 413296
rect 66622 413284 66628 413296
rect 55180 413256 66628 413284
rect 55180 413244 55186 413256
rect 66622 413244 66628 413256
rect 66680 413244 66686 413296
rect 184842 412632 184848 412684
rect 184900 412672 184906 412684
rect 191742 412672 191748 412684
rect 184900 412644 191748 412672
rect 184900 412632 184906 412644
rect 191742 412632 191748 412644
rect 191800 412632 191806 412684
rect 255406 412428 255412 412480
rect 255464 412468 255470 412480
rect 258258 412468 258264 412480
rect 255464 412440 258264 412468
rect 255464 412428 255470 412440
rect 258258 412428 258264 412440
rect 258316 412428 258322 412480
rect 115014 411884 115020 411936
rect 115072 411924 115078 411936
rect 122834 411924 122840 411936
rect 115072 411896 122840 411924
rect 115072 411884 115078 411896
rect 122834 411884 122840 411896
rect 122892 411924 122898 411936
rect 123478 411924 123484 411936
rect 122892 411896 123484 411924
rect 122892 411884 122898 411896
rect 123478 411884 123484 411896
rect 123536 411884 123542 411936
rect 147030 411884 147036 411936
rect 147088 411924 147094 411936
rect 158806 411924 158812 411936
rect 147088 411896 158812 411924
rect 147088 411884 147094 411896
rect 158806 411884 158812 411896
rect 158864 411884 158870 411936
rect 260098 411884 260104 411936
rect 260156 411924 260162 411936
rect 288710 411924 288716 411936
rect 260156 411896 288716 411924
rect 260156 411884 260162 411896
rect 288710 411884 288716 411896
rect 288768 411884 288774 411936
rect 61930 411272 61936 411324
rect 61988 411312 61994 411324
rect 66898 411312 66904 411324
rect 61988 411284 66904 411312
rect 61988 411272 61994 411284
rect 66898 411272 66904 411284
rect 66956 411272 66962 411324
rect 158806 411272 158812 411324
rect 158864 411312 158870 411324
rect 159358 411312 159364 411324
rect 158864 411284 159364 411312
rect 158864 411272 158870 411284
rect 159358 411272 159364 411284
rect 159416 411312 159422 411324
rect 192846 411312 192852 411324
rect 159416 411284 192852 411312
rect 159416 411272 159422 411284
rect 192846 411272 192852 411284
rect 192904 411272 192910 411324
rect 52178 411204 52184 411256
rect 52236 411244 52242 411256
rect 66806 411244 66812 411256
rect 52236 411216 66812 411244
rect 52236 411204 52242 411216
rect 66806 411204 66812 411216
rect 66864 411204 66870 411256
rect 115566 411204 115572 411256
rect 115624 411244 115630 411256
rect 122190 411244 122196 411256
rect 115624 411216 122196 411244
rect 115624 411204 115630 411216
rect 122190 411204 122196 411216
rect 122248 411204 122254 411256
rect 44082 410524 44088 410576
rect 44140 410564 44146 410576
rect 52178 410564 52184 410576
rect 44140 410536 52184 410564
rect 44140 410524 44146 410536
rect 52178 410524 52184 410536
rect 52236 410524 52242 410576
rect 177850 410524 177856 410576
rect 177908 410564 177914 410576
rect 190454 410564 190460 410576
rect 177908 410536 190460 410564
rect 177908 410524 177914 410536
rect 190454 410524 190460 410536
rect 190512 410524 190518 410576
rect 187510 410388 187516 410440
rect 187568 410428 187574 410440
rect 189074 410428 189080 410440
rect 187568 410400 189080 410428
rect 187568 410388 187574 410400
rect 189074 410388 189080 410400
rect 189132 410388 189138 410440
rect 2774 410184 2780 410236
rect 2832 410224 2838 410236
rect 4798 410224 4804 410236
rect 2832 410196 4804 410224
rect 2832 410184 2838 410196
rect 4798 410184 4804 410196
rect 4856 410184 4862 410236
rect 121454 409844 121460 409896
rect 121512 409884 121518 409896
rect 155770 409884 155776 409896
rect 121512 409856 155776 409884
rect 121512 409844 121518 409856
rect 155770 409844 155776 409856
rect 155828 409884 155834 409896
rect 160094 409884 160100 409896
rect 155828 409856 160100 409884
rect 155828 409844 155834 409856
rect 160094 409844 160100 409856
rect 160152 409844 160158 409896
rect 115842 409776 115848 409828
rect 115900 409816 115906 409828
rect 126238 409816 126244 409828
rect 115900 409788 126244 409816
rect 115900 409776 115906 409788
rect 126238 409776 126244 409788
rect 126296 409776 126302 409828
rect 49602 408484 49608 408536
rect 49660 408524 49666 408536
rect 66806 408524 66812 408536
rect 49660 408496 66812 408524
rect 49660 408484 49666 408496
rect 66806 408484 66812 408496
rect 66864 408484 66870 408536
rect 115842 408484 115848 408536
rect 115900 408524 115906 408536
rect 151170 408524 151176 408536
rect 115900 408496 151176 408524
rect 115900 408484 115906 408496
rect 151170 408484 151176 408496
rect 151228 408484 151234 408536
rect 191742 408524 191748 408536
rect 186332 408496 191748 408524
rect 186332 408468 186360 408496
rect 191742 408484 191748 408496
rect 191800 408484 191806 408536
rect 255406 408484 255412 408536
rect 255464 408524 255470 408536
rect 270770 408524 270776 408536
rect 255464 408496 270776 408524
rect 255464 408484 255470 408496
rect 270770 408484 270776 408496
rect 270828 408524 270834 408536
rect 276106 408524 276112 408536
rect 270828 408496 276112 408524
rect 270828 408484 270834 408496
rect 276106 408484 276112 408496
rect 276164 408484 276170 408536
rect 39850 408416 39856 408468
rect 39908 408456 39914 408468
rect 48222 408456 48228 408468
rect 39908 408428 48228 408456
rect 39908 408416 39914 408428
rect 48222 408416 48228 408428
rect 48280 408456 48286 408468
rect 66898 408456 66904 408468
rect 48280 408428 66904 408456
rect 48280 408416 48286 408428
rect 66898 408416 66904 408428
rect 66956 408416 66962 408468
rect 140682 408416 140688 408468
rect 140740 408456 140746 408468
rect 186314 408456 186320 408468
rect 140740 408428 186320 408456
rect 140740 408416 140746 408428
rect 186314 408416 186320 408428
rect 186372 408416 186378 408468
rect 255406 407804 255412 407856
rect 255464 407844 255470 407856
rect 259638 407844 259644 407856
rect 255464 407816 259644 407844
rect 255464 407804 255470 407816
rect 259638 407804 259644 407816
rect 259696 407844 259702 407856
rect 265066 407844 265072 407856
rect 259696 407816 265072 407844
rect 259696 407804 259702 407816
rect 265066 407804 265072 407816
rect 265124 407804 265130 407856
rect 159910 407736 159916 407788
rect 159968 407776 159974 407788
rect 166994 407776 167000 407788
rect 159968 407748 167000 407776
rect 159968 407736 159974 407748
rect 166994 407736 167000 407748
rect 167052 407736 167058 407788
rect 255498 407736 255504 407788
rect 255556 407776 255562 407788
rect 273530 407776 273536 407788
rect 255556 407748 273536 407776
rect 255556 407736 255562 407748
rect 273530 407736 273536 407748
rect 273588 407736 273594 407788
rect 166994 407124 167000 407176
rect 167052 407164 167058 407176
rect 191650 407164 191656 407176
rect 167052 407136 191656 407164
rect 167052 407124 167058 407136
rect 191650 407124 191656 407136
rect 191708 407124 191714 407176
rect 113082 407056 113088 407108
rect 113140 407096 113146 407108
rect 131758 407096 131764 407108
rect 113140 407068 131764 407096
rect 113140 407056 113146 407068
rect 131758 407056 131764 407068
rect 131816 407056 131822 407108
rect 57882 406376 57888 406428
rect 57940 406416 57946 406428
rect 64782 406416 64788 406428
rect 57940 406388 64788 406416
rect 57940 406376 57946 406388
rect 64782 406376 64788 406388
rect 64840 406416 64846 406428
rect 66806 406416 66812 406428
rect 64840 406388 66812 406416
rect 64840 406376 64846 406388
rect 66806 406376 66812 406388
rect 66864 406376 66870 406428
rect 154482 406376 154488 406428
rect 154540 406416 154546 406428
rect 191742 406416 191748 406428
rect 154540 406388 191748 406416
rect 154540 406376 154546 406388
rect 191742 406376 191748 406388
rect 191800 406376 191806 406428
rect 255498 405696 255504 405748
rect 255556 405736 255562 405748
rect 276106 405736 276112 405748
rect 255556 405708 276112 405736
rect 255556 405696 255562 405708
rect 276106 405696 276112 405708
rect 276164 405696 276170 405748
rect 115842 405628 115848 405680
rect 115900 405668 115906 405680
rect 121454 405668 121460 405680
rect 115900 405640 121460 405668
rect 115900 405628 115906 405640
rect 121454 405628 121460 405640
rect 121512 405628 121518 405680
rect 152918 405628 152924 405680
rect 152976 405668 152982 405680
rect 154482 405668 154488 405680
rect 152976 405640 154488 405668
rect 152976 405628 152982 405640
rect 154482 405628 154488 405640
rect 154540 405628 154546 405680
rect 153838 404444 153844 404456
rect 142126 404416 153844 404444
rect 63218 404336 63224 404388
rect 63276 404376 63282 404388
rect 66806 404376 66812 404388
rect 63276 404348 66812 404376
rect 63276 404336 63282 404348
rect 66806 404336 66812 404348
rect 66864 404336 66870 404388
rect 115842 404336 115848 404388
rect 115900 404376 115906 404388
rect 142126 404376 142154 404416
rect 153838 404404 153844 404416
rect 153896 404404 153902 404456
rect 115900 404348 142154 404376
rect 115900 404336 115906 404348
rect 162210 404336 162216 404388
rect 162268 404376 162274 404388
rect 162578 404376 162584 404388
rect 162268 404348 162584 404376
rect 162268 404336 162274 404348
rect 162578 404336 162584 404348
rect 162636 404376 162642 404388
rect 177482 404376 177488 404388
rect 162636 404348 177488 404376
rect 162636 404336 162642 404348
rect 177482 404336 177488 404348
rect 177540 404336 177546 404388
rect 164050 404268 164056 404320
rect 164108 404308 164114 404320
rect 169754 404308 169760 404320
rect 164108 404280 169760 404308
rect 164108 404268 164114 404280
rect 169754 404268 169760 404280
rect 169812 404268 169818 404320
rect 53650 403588 53656 403640
rect 53708 403628 53714 403640
rect 67634 403628 67640 403640
rect 53708 403600 67640 403628
rect 53708 403588 53714 403600
rect 67634 403588 67640 403600
rect 67692 403588 67698 403640
rect 119982 403588 119988 403640
rect 120040 403628 120046 403640
rect 162578 403628 162584 403640
rect 120040 403600 162584 403628
rect 120040 403588 120046 403600
rect 162578 403588 162584 403600
rect 162636 403588 162642 403640
rect 172422 403588 172428 403640
rect 172480 403628 172486 403640
rect 182910 403628 182916 403640
rect 172480 403600 182916 403628
rect 172480 403588 172486 403600
rect 182910 403588 182916 403600
rect 182968 403588 182974 403640
rect 115842 402976 115848 403028
rect 115900 403016 115906 403028
rect 148318 403016 148324 403028
rect 115900 402988 148324 403016
rect 115900 402976 115906 402988
rect 148318 402976 148324 402988
rect 148376 402976 148382 403028
rect 169754 402976 169760 403028
rect 169812 403016 169818 403028
rect 191742 403016 191748 403028
rect 169812 402988 191748 403016
rect 169812 402976 169818 402988
rect 191742 402976 191748 402988
rect 191800 402976 191806 403028
rect 256878 402976 256884 403028
rect 256936 403016 256942 403028
rect 291286 403016 291292 403028
rect 256936 402988 291292 403016
rect 256936 402976 256942 402988
rect 291286 402976 291292 402988
rect 291344 402976 291350 403028
rect 255314 402908 255320 402960
rect 255372 402948 255378 402960
rect 287146 402948 287152 402960
rect 255372 402920 287152 402948
rect 255372 402908 255378 402920
rect 287146 402908 287152 402920
rect 287204 402908 287210 402960
rect 185578 401820 185584 401872
rect 185636 401860 185642 401872
rect 193122 401860 193128 401872
rect 185636 401832 193128 401860
rect 185636 401820 185642 401832
rect 193122 401820 193128 401832
rect 193180 401820 193186 401872
rect 116578 401616 116584 401668
rect 116636 401656 116642 401668
rect 181438 401656 181444 401668
rect 116636 401628 181444 401656
rect 116636 401616 116642 401628
rect 181438 401616 181444 401628
rect 181496 401616 181502 401668
rect 186038 401004 186044 401056
rect 186096 401044 186102 401056
rect 186958 401044 186964 401056
rect 186096 401016 186964 401044
rect 186096 401004 186102 401016
rect 186958 401004 186964 401016
rect 187016 401004 187022 401056
rect 118878 400868 118884 400920
rect 118936 400908 118942 400920
rect 143534 400908 143540 400920
rect 118936 400880 143540 400908
rect 118936 400868 118942 400880
rect 143534 400868 143540 400880
rect 143592 400868 143598 400920
rect 172054 400868 172060 400920
rect 172112 400908 172118 400920
rect 191558 400908 191564 400920
rect 172112 400880 191564 400908
rect 172112 400868 172118 400880
rect 191558 400868 191564 400880
rect 191616 400868 191622 400920
rect 115566 400664 115572 400716
rect 115624 400704 115630 400716
rect 119982 400704 119988 400716
rect 115624 400676 119988 400704
rect 115624 400664 115630 400676
rect 119982 400664 119988 400676
rect 120040 400664 120046 400716
rect 115750 400528 115756 400580
rect 115808 400568 115814 400580
rect 122190 400568 122196 400580
rect 115808 400540 122196 400568
rect 115808 400528 115814 400540
rect 122190 400528 122196 400540
rect 122248 400528 122254 400580
rect 59078 400188 59084 400240
rect 59136 400228 59142 400240
rect 66806 400228 66812 400240
rect 59136 400200 66812 400228
rect 59136 400188 59142 400200
rect 66806 400188 66812 400200
rect 66864 400188 66870 400240
rect 123662 400188 123668 400240
rect 123720 400228 123726 400240
rect 186038 400228 186044 400240
rect 123720 400200 186044 400228
rect 123720 400188 123726 400200
rect 186038 400188 186044 400200
rect 186096 400188 186102 400240
rect 255406 400188 255412 400240
rect 255464 400228 255470 400240
rect 280430 400228 280436 400240
rect 255464 400200 280436 400228
rect 255464 400188 255470 400200
rect 280430 400188 280436 400200
rect 280488 400188 280494 400240
rect 148962 399440 148968 399492
rect 149020 399480 149026 399492
rect 181530 399480 181536 399492
rect 149020 399452 181536 399480
rect 149020 399440 149026 399452
rect 181530 399440 181536 399452
rect 181588 399440 181594 399492
rect 115842 398896 115848 398948
rect 115900 398936 115906 398948
rect 137278 398936 137284 398948
rect 115900 398908 137284 398936
rect 115900 398896 115906 398908
rect 137278 398896 137284 398908
rect 137336 398896 137342 398948
rect 53650 398828 53656 398880
rect 53708 398868 53714 398880
rect 66806 398868 66812 398880
rect 53708 398840 66812 398868
rect 53708 398828 53714 398840
rect 66806 398828 66812 398840
rect 66864 398828 66870 398880
rect 128998 398828 129004 398880
rect 129056 398868 129062 398880
rect 190270 398868 190276 398880
rect 129056 398840 190276 398868
rect 129056 398828 129062 398840
rect 190270 398828 190276 398840
rect 190328 398868 190334 398880
rect 191742 398868 191748 398880
rect 190328 398840 191748 398868
rect 190328 398828 190334 398840
rect 191742 398828 191748 398840
rect 191800 398828 191806 398880
rect 255406 398828 255412 398880
rect 255464 398868 255470 398880
rect 255464 398840 267734 398868
rect 255464 398828 255470 398840
rect 60642 398760 60648 398812
rect 60700 398800 60706 398812
rect 65886 398800 65892 398812
rect 60700 398772 65892 398800
rect 60700 398760 60706 398772
rect 65886 398760 65892 398772
rect 65944 398800 65950 398812
rect 66530 398800 66536 398812
rect 65944 398772 66536 398800
rect 65944 398760 65950 398772
rect 66530 398760 66536 398772
rect 66588 398760 66594 398812
rect 267706 398800 267734 398840
rect 268378 398800 268384 398812
rect 267706 398772 268384 398800
rect 268378 398760 268384 398772
rect 268436 398800 268442 398812
rect 274818 398800 274824 398812
rect 268436 398772 274824 398800
rect 268436 398760 268442 398772
rect 274818 398760 274824 398772
rect 274876 398760 274882 398812
rect 115842 398284 115848 398336
rect 115900 398324 115906 398336
rect 116026 398324 116032 398336
rect 115900 398296 116032 398324
rect 115900 398284 115906 398296
rect 116026 398284 116032 398296
rect 116084 398324 116090 398336
rect 118878 398324 118884 398336
rect 116084 398296 118884 398324
rect 116084 398284 116090 398296
rect 118878 398284 118884 398296
rect 118936 398284 118942 398336
rect 255406 398216 255412 398268
rect 255464 398256 255470 398268
rect 258902 398256 258908 398268
rect 255464 398228 258908 398256
rect 255464 398216 255470 398228
rect 258902 398216 258908 398228
rect 258960 398216 258966 398268
rect 118878 398148 118884 398200
rect 118936 398188 118942 398200
rect 147490 398188 147496 398200
rect 118936 398160 147496 398188
rect 118936 398148 118942 398160
rect 147490 398148 147496 398160
rect 147548 398188 147554 398200
rect 173250 398188 173256 398200
rect 147548 398160 173256 398188
rect 147548 398148 147554 398160
rect 173250 398148 173256 398160
rect 173308 398148 173314 398200
rect 174998 398148 175004 398200
rect 175056 398188 175062 398200
rect 180150 398188 180156 398200
rect 175056 398160 180156 398188
rect 175056 398148 175062 398160
rect 180150 398148 180156 398160
rect 180208 398148 180214 398200
rect 145650 398080 145656 398132
rect 145708 398120 145714 398132
rect 145708 398092 180794 398120
rect 145708 398080 145714 398092
rect 180766 398052 180794 398092
rect 188890 398080 188896 398132
rect 188948 398120 188954 398132
rect 189718 398120 189724 398132
rect 188948 398092 189724 398120
rect 188948 398080 188954 398092
rect 189718 398080 189724 398092
rect 189776 398080 189782 398132
rect 191742 398120 191748 398132
rect 190426 398092 191748 398120
rect 183554 398052 183560 398064
rect 180766 398024 183560 398052
rect 183554 398012 183560 398024
rect 183612 398052 183618 398064
rect 190426 398052 190454 398092
rect 191742 398080 191748 398092
rect 191800 398080 191806 398132
rect 265618 398080 265624 398132
rect 265676 398120 265682 398132
rect 275002 398120 275008 398132
rect 265676 398092 275008 398120
rect 265676 398080 265682 398092
rect 275002 398080 275008 398092
rect 275060 398080 275066 398132
rect 183612 398024 190454 398052
rect 183612 398012 183618 398024
rect 36538 397468 36544 397520
rect 36596 397508 36602 397520
rect 67082 397508 67088 397520
rect 36596 397480 67088 397508
rect 36596 397468 36602 397480
rect 67082 397468 67088 397480
rect 67140 397468 67146 397520
rect 163498 397400 163504 397452
rect 163556 397440 163562 397452
rect 163958 397440 163964 397452
rect 163556 397412 163964 397440
rect 163556 397400 163562 397412
rect 163958 397400 163964 397412
rect 164016 397400 164022 397452
rect 140038 396720 140044 396772
rect 140096 396760 140102 396772
rect 180518 396760 180524 396772
rect 140096 396732 180524 396760
rect 140096 396720 140102 396732
rect 180518 396720 180524 396732
rect 180576 396760 180582 396772
rect 187142 396760 187148 396772
rect 180576 396732 187148 396760
rect 180576 396720 180582 396732
rect 187142 396720 187148 396732
rect 187200 396720 187206 396772
rect 115106 396516 115112 396568
rect 115164 396556 115170 396568
rect 118878 396556 118884 396568
rect 115164 396528 118884 396556
rect 115164 396516 115170 396528
rect 118878 396516 118884 396528
rect 118936 396516 118942 396568
rect 115566 396040 115572 396092
rect 115624 396080 115630 396092
rect 122098 396080 122104 396092
rect 115624 396052 122104 396080
rect 115624 396040 115630 396052
rect 122098 396040 122104 396052
rect 122156 396040 122162 396092
rect 163498 396040 163504 396092
rect 163556 396080 163562 396092
rect 192478 396080 192484 396092
rect 163556 396052 192484 396080
rect 163556 396040 163562 396052
rect 192478 396040 192484 396052
rect 192536 396040 192542 396092
rect 57698 395292 57704 395344
rect 57756 395332 57762 395344
rect 67266 395332 67272 395344
rect 57756 395304 67272 395332
rect 57756 395292 57762 395304
rect 67266 395292 67272 395304
rect 67324 395292 67330 395344
rect 168282 395292 168288 395344
rect 168340 395332 168346 395344
rect 176102 395332 176108 395344
rect 168340 395304 176108 395332
rect 168340 395292 168346 395304
rect 176102 395292 176108 395304
rect 176160 395292 176166 395344
rect 164050 394952 164056 395004
rect 164108 394992 164114 395004
rect 164970 394992 164976 395004
rect 164108 394964 164976 394992
rect 164108 394952 164114 394964
rect 164970 394952 164976 394964
rect 165028 394952 165034 395004
rect 115842 394748 115848 394800
rect 115900 394788 115906 394800
rect 151078 394788 151084 394800
rect 115900 394760 151084 394788
rect 115900 394748 115906 394760
rect 151078 394748 151084 394760
rect 151136 394748 151142 394800
rect 157978 394720 157984 394732
rect 115952 394692 157984 394720
rect 115842 394612 115848 394664
rect 115900 394652 115906 394664
rect 115952 394652 115980 394692
rect 157978 394680 157984 394692
rect 158036 394680 158042 394732
rect 161474 394680 161480 394732
rect 161532 394720 161538 394732
rect 162670 394720 162676 394732
rect 161532 394692 162676 394720
rect 161532 394680 161538 394692
rect 162670 394680 162676 394692
rect 162728 394720 162734 394732
rect 191834 394720 191840 394732
rect 162728 394692 191840 394720
rect 162728 394680 162734 394692
rect 191834 394680 191840 394692
rect 191892 394680 191898 394732
rect 115900 394624 115980 394652
rect 115900 394612 115906 394624
rect 155310 394612 155316 394664
rect 155368 394652 155374 394664
rect 155954 394652 155960 394664
rect 155368 394624 155960 394652
rect 155368 394612 155374 394624
rect 155954 394612 155960 394624
rect 156012 394612 156018 394664
rect 117222 393932 117228 393984
rect 117280 393972 117286 393984
rect 136634 393972 136640 393984
rect 117280 393944 136640 393972
rect 117280 393932 117286 393944
rect 136634 393932 136640 393944
rect 136692 393932 136698 393984
rect 61838 393388 61844 393440
rect 61896 393428 61902 393440
rect 65978 393428 65984 393440
rect 61896 393400 65984 393428
rect 61896 393388 61902 393400
rect 65978 393388 65984 393400
rect 66036 393388 66042 393440
rect 177390 393320 177396 393372
rect 177448 393360 177454 393372
rect 191006 393360 191012 393372
rect 177448 393332 191012 393360
rect 177448 393320 177454 393332
rect 191006 393320 191012 393332
rect 191064 393320 191070 393372
rect 255498 393320 255504 393372
rect 255556 393360 255562 393372
rect 278958 393360 278964 393372
rect 255556 393332 278964 393360
rect 255556 393320 255562 393332
rect 278958 393320 278964 393332
rect 279016 393320 279022 393372
rect 160094 393252 160100 393304
rect 160152 393292 160158 393304
rect 161382 393292 161388 393304
rect 160152 393264 161388 393292
rect 160152 393252 160158 393264
rect 161382 393252 161388 393264
rect 161440 393292 161446 393304
rect 191926 393292 191932 393304
rect 161440 393264 191932 393292
rect 161440 393252 161446 393264
rect 191926 393252 191932 393264
rect 191984 393252 191990 393304
rect 148410 392640 148416 392692
rect 148468 392680 148474 392692
rect 161474 392680 161480 392692
rect 148468 392652 161480 392680
rect 148468 392640 148474 392652
rect 161474 392640 161480 392652
rect 161532 392640 161538 392692
rect 144178 392572 144184 392624
rect 144236 392612 144242 392624
rect 160094 392612 160100 392624
rect 144236 392584 160100 392612
rect 144236 392572 144242 392584
rect 160094 392572 160100 392584
rect 160152 392572 160158 392624
rect 253658 392572 253664 392624
rect 253716 392612 253722 392624
rect 279418 392612 279424 392624
rect 253716 392584 279424 392612
rect 253716 392572 253722 392584
rect 279418 392572 279424 392584
rect 279476 392572 279482 392624
rect 115934 392300 115940 392352
rect 115992 392340 115998 392352
rect 117222 392340 117228 392352
rect 115992 392312 117228 392340
rect 115992 392300 115998 392312
rect 117222 392300 117228 392312
rect 117280 392300 117286 392352
rect 57698 391960 57704 392012
rect 57756 392000 57762 392012
rect 66806 392000 66812 392012
rect 57756 391972 66812 392000
rect 57756 391960 57762 391972
rect 66806 391960 66812 391972
rect 66864 391960 66870 392012
rect 115842 391960 115848 392012
rect 115900 392000 115906 392012
rect 145650 392000 145656 392012
rect 115900 391972 145656 392000
rect 115900 391960 115906 391972
rect 145650 391960 145656 391972
rect 145708 391960 145714 392012
rect 162210 391960 162216 392012
rect 162268 392000 162274 392012
rect 171870 392000 171876 392012
rect 162268 391972 171876 392000
rect 162268 391960 162274 391972
rect 171870 391960 171876 391972
rect 171928 392000 171934 392012
rect 172422 392000 172428 392012
rect 171928 391972 172428 392000
rect 171928 391960 171934 391972
rect 172422 391960 172428 391972
rect 172480 391960 172486 392012
rect 254302 391960 254308 392012
rect 254360 392000 254366 392012
rect 255314 392000 255320 392012
rect 254360 391972 255320 392000
rect 254360 391960 254366 391972
rect 255314 391960 255320 391972
rect 255372 391960 255378 392012
rect 78646 391496 82814 391524
rect 78646 391456 78674 391496
rect 77266 391428 78674 391456
rect 82786 391456 82814 391496
rect 82786 391428 85574 391456
rect 35158 391280 35164 391332
rect 35216 391320 35222 391332
rect 68554 391320 68560 391332
rect 35216 391292 68560 391320
rect 35216 391280 35222 391292
rect 68554 391280 68560 391292
rect 68612 391280 68618 391332
rect 4798 391212 4804 391264
rect 4856 391252 4862 391264
rect 77266 391252 77294 391428
rect 85546 391388 85574 391428
rect 85546 391360 86954 391388
rect 4856 391224 77294 391252
rect 86926 391252 86954 391360
rect 93826 391360 106366 391388
rect 93826 391252 93854 391360
rect 86926 391224 93854 391252
rect 99208 391292 99374 391320
rect 4856 391212 4862 391224
rect 86926 391156 93854 391184
rect 68554 391076 68560 391128
rect 68612 391116 68618 391128
rect 86926 391116 86954 391156
rect 68612 391088 86954 391116
rect 68612 391076 68618 391088
rect 93826 390980 93854 391156
rect 93946 390980 93952 390992
rect 93826 390952 93952 390980
rect 93946 390940 93952 390952
rect 94004 390940 94010 390992
rect 94958 390940 94964 390992
rect 95016 390980 95022 390992
rect 99208 390980 99236 391292
rect 99346 391252 99374 391292
rect 99346 391224 106274 391252
rect 95016 390952 99236 390980
rect 95016 390940 95022 390952
rect 106246 390912 106274 391224
rect 106338 390980 106366 391360
rect 112714 391280 112720 391332
rect 112772 391320 112778 391332
rect 116578 391320 116584 391332
rect 112772 391292 116584 391320
rect 112772 391280 112778 391292
rect 116578 391280 116584 391292
rect 116636 391280 116642 391332
rect 253566 391280 253572 391332
rect 253624 391320 253630 391332
rect 295334 391320 295340 391332
rect 253624 391292 295340 391320
rect 253624 391280 253630 391292
rect 295334 391280 295340 391292
rect 295392 391280 295398 391332
rect 173618 391212 173624 391264
rect 173676 391252 173682 391264
rect 173676 391224 180794 391252
rect 173676 391212 173682 391224
rect 107286 390980 107292 390992
rect 106338 390952 107292 390980
rect 107286 390940 107292 390952
rect 107344 390940 107350 390992
rect 180766 390980 180794 391224
rect 264238 391212 264244 391264
rect 264296 391252 264302 391264
rect 280338 391252 280344 391264
rect 264296 391224 280344 391252
rect 264296 391212 264302 391224
rect 280338 391212 280344 391224
rect 280396 391212 280402 391264
rect 286318 391212 286324 391264
rect 286376 391252 286382 391264
rect 292574 391252 292580 391264
rect 286376 391224 292580 391252
rect 286376 391212 286382 391224
rect 292574 391212 292580 391224
rect 292632 391252 292638 391264
rect 580258 391252 580264 391264
rect 292632 391224 580264 391252
rect 292632 391212 292638 391224
rect 580258 391212 580264 391224
rect 580316 391212 580322 391264
rect 194134 390980 194140 390992
rect 180766 390952 194140 390980
rect 194134 390940 194140 390952
rect 194192 390940 194198 390992
rect 112714 390912 112720 390924
rect 106246 390884 112720 390912
rect 112714 390872 112720 390884
rect 112772 390872 112778 390924
rect 191834 390872 191840 390924
rect 191892 390912 191898 390924
rect 195974 390912 195980 390924
rect 191892 390884 195980 390912
rect 191892 390872 191898 390884
rect 195974 390872 195980 390884
rect 196032 390872 196038 390924
rect 171962 390600 171968 390652
rect 172020 390640 172026 390652
rect 173618 390640 173624 390652
rect 172020 390612 173624 390640
rect 172020 390600 172026 390612
rect 173618 390600 173624 390612
rect 173676 390600 173682 390652
rect 158438 390532 158444 390584
rect 158496 390572 158502 390584
rect 163590 390572 163596 390584
rect 158496 390544 163596 390572
rect 158496 390532 158502 390544
rect 163590 390532 163596 390544
rect 163648 390572 163654 390584
rect 191742 390572 191748 390584
rect 163648 390544 191748 390572
rect 163648 390532 163654 390544
rect 191742 390532 191748 390544
rect 191800 390532 191806 390584
rect 251818 390532 251824 390584
rect 251876 390572 251882 390584
rect 259638 390572 259644 390584
rect 251876 390544 259644 390572
rect 251876 390532 251882 390544
rect 259638 390532 259644 390544
rect 259696 390532 259702 390584
rect 67634 390124 67640 390176
rect 67692 390164 67698 390176
rect 68784 390164 68790 390176
rect 67692 390136 68790 390164
rect 67692 390124 67698 390136
rect 68784 390124 68790 390136
rect 68842 390124 68848 390176
rect 154482 389852 154488 389904
rect 154540 389892 154546 389904
rect 164878 389892 164884 389904
rect 154540 389864 164884 389892
rect 154540 389852 154546 389864
rect 164878 389852 164884 389864
rect 164936 389852 164942 389904
rect 160094 389784 160100 389836
rect 160152 389824 160158 389836
rect 160738 389824 160744 389836
rect 160152 389796 160744 389824
rect 160152 389784 160158 389796
rect 160738 389784 160744 389796
rect 160796 389824 160802 389836
rect 186406 389824 186412 389836
rect 160796 389796 186412 389824
rect 160796 389784 160802 389796
rect 186406 389784 186412 389796
rect 186464 389784 186470 389836
rect 40678 389240 40684 389292
rect 40736 389280 40742 389292
rect 100754 389280 100760 389292
rect 40736 389252 100760 389280
rect 40736 389240 40742 389252
rect 100754 389240 100760 389252
rect 100812 389240 100818 389292
rect 110782 389240 110788 389292
rect 110840 389280 110846 389292
rect 141418 389280 141424 389292
rect 110840 389252 141424 389280
rect 110840 389240 110846 389252
rect 141418 389240 141424 389252
rect 141476 389240 141482 389292
rect 187142 389240 187148 389292
rect 187200 389280 187206 389292
rect 215294 389280 215300 389292
rect 187200 389252 215300 389280
rect 187200 389240 187206 389252
rect 215294 389240 215300 389252
rect 215352 389240 215358 389292
rect 238754 389240 238760 389292
rect 238812 389280 238818 389292
rect 239030 389280 239036 389292
rect 238812 389252 239036 389280
rect 238812 389240 238818 389252
rect 239030 389240 239036 389252
rect 239088 389280 239094 389292
rect 260098 389280 260104 389292
rect 239088 389252 260104 389280
rect 239088 389240 239094 389252
rect 260098 389240 260104 389252
rect 260156 389240 260162 389292
rect 17218 389172 17224 389224
rect 17276 389212 17282 389224
rect 81710 389212 81716 389224
rect 17276 389184 81716 389212
rect 17276 389172 17282 389184
rect 81710 389172 81716 389184
rect 81768 389172 81774 389224
rect 98914 389172 98920 389224
rect 98972 389212 98978 389224
rect 160094 389212 160100 389224
rect 98972 389184 160100 389212
rect 98972 389172 98978 389184
rect 160094 389172 160100 389184
rect 160152 389172 160158 389224
rect 178862 389172 178868 389224
rect 178920 389212 178926 389224
rect 200206 389212 200212 389224
rect 178920 389184 200212 389212
rect 178920 389172 178926 389184
rect 200206 389172 200212 389184
rect 200264 389172 200270 389224
rect 201586 389172 201592 389224
rect 201644 389212 201650 389224
rect 267826 389212 267832 389224
rect 201644 389184 267832 389212
rect 201644 389172 201650 389184
rect 267826 389172 267832 389184
rect 267884 389172 267890 389224
rect 169018 389104 169024 389156
rect 169076 389144 169082 389156
rect 169478 389144 169484 389156
rect 169076 389116 169484 389144
rect 169076 389104 169082 389116
rect 169478 389104 169484 389116
rect 169536 389144 169542 389156
rect 205910 389144 205916 389156
rect 169536 389116 205916 389144
rect 169536 389104 169542 389116
rect 205910 389104 205916 389116
rect 205968 389104 205974 389156
rect 253382 389104 253388 389156
rect 253440 389144 253446 389156
rect 276198 389144 276204 389156
rect 253440 389116 276204 389144
rect 253440 389104 253446 389116
rect 276198 389104 276204 389116
rect 276256 389104 276262 389156
rect 172422 389036 172428 389088
rect 172480 389076 172486 389088
rect 202966 389076 202972 389088
rect 172480 389048 202972 389076
rect 172480 389036 172486 389048
rect 202966 389036 202972 389048
rect 203024 389036 203030 389088
rect 250714 389036 250720 389088
rect 250772 389076 250778 389088
rect 253658 389076 253664 389088
rect 250772 389048 253664 389076
rect 250772 389036 250778 389048
rect 253658 389036 253664 389048
rect 253716 389036 253722 389088
rect 164878 388560 164884 388612
rect 164936 388600 164942 388612
rect 171778 388600 171784 388612
rect 164936 388572 171784 388600
rect 164936 388560 164942 388572
rect 171778 388560 171784 388572
rect 171836 388560 171842 388612
rect 59170 388424 59176 388476
rect 59228 388464 59234 388476
rect 59228 388436 64874 388464
rect 59228 388424 59234 388436
rect 64846 388396 64874 388436
rect 67358 388424 67364 388476
rect 67416 388464 67422 388476
rect 71038 388464 71044 388476
rect 67416 388436 71044 388464
rect 67416 388424 67422 388436
rect 71038 388424 71044 388436
rect 71096 388424 71102 388476
rect 82722 388424 82728 388476
rect 82780 388464 82786 388476
rect 108390 388464 108396 388476
rect 82780 388436 108396 388464
rect 82780 388424 82786 388436
rect 108390 388424 108396 388436
rect 108448 388424 108454 388476
rect 233326 388424 233332 388476
rect 233384 388464 233390 388476
rect 245838 388464 245844 388476
rect 233384 388436 245844 388464
rect 233384 388424 233390 388436
rect 245838 388424 245844 388436
rect 245896 388424 245902 388476
rect 247678 388424 247684 388476
rect 247736 388464 247742 388476
rect 251358 388464 251364 388476
rect 247736 388436 251364 388464
rect 247736 388424 247742 388436
rect 251358 388424 251364 388436
rect 251416 388424 251422 388476
rect 262858 388424 262864 388476
rect 262916 388464 262922 388476
rect 291378 388464 291384 388476
rect 262916 388436 291384 388464
rect 262916 388424 262922 388436
rect 291378 388424 291384 388436
rect 291436 388424 291442 388476
rect 71682 388396 71688 388408
rect 64846 388368 71688 388396
rect 71682 388356 71688 388368
rect 71740 388356 71746 388408
rect 238110 388356 238116 388408
rect 238168 388396 238174 388408
rect 239398 388396 239404 388408
rect 238168 388368 239404 388396
rect 238168 388356 238174 388368
rect 239398 388356 239404 388368
rect 239456 388356 239462 388408
rect 71682 387948 71688 388000
rect 71740 387988 71746 388000
rect 72510 387988 72516 388000
rect 71740 387960 72516 387988
rect 71740 387948 71746 387960
rect 72510 387948 72516 387960
rect 72568 387948 72574 388000
rect 83182 387880 83188 387932
rect 83240 387920 83246 387932
rect 84102 387920 84108 387932
rect 83240 387892 84108 387920
rect 83240 387880 83246 387892
rect 84102 387880 84108 387892
rect 84160 387880 84166 387932
rect 70854 387812 70860 387864
rect 70912 387852 70918 387864
rect 72510 387852 72516 387864
rect 70912 387824 72516 387852
rect 70912 387812 70918 387824
rect 72510 387812 72516 387824
rect 72568 387812 72574 387864
rect 77202 387812 77208 387864
rect 77260 387852 77266 387864
rect 78030 387852 78036 387864
rect 77260 387824 78036 387852
rect 77260 387812 77266 387824
rect 78030 387812 78036 387824
rect 78088 387812 78094 387864
rect 123570 387852 123576 387864
rect 122806 387824 123576 387852
rect 88242 387744 88248 387796
rect 88300 387784 88306 387796
rect 92014 387784 92020 387796
rect 88300 387756 92020 387784
rect 88300 387744 88306 387756
rect 92014 387744 92020 387756
rect 92072 387744 92078 387796
rect 93394 387744 93400 387796
rect 93452 387784 93458 387796
rect 122806 387784 122834 387824
rect 123570 387812 123576 387824
rect 123628 387852 123634 387864
rect 125594 387852 125600 387864
rect 123628 387824 125600 387852
rect 123628 387812 123634 387824
rect 125594 387812 125600 387824
rect 125652 387812 125658 387864
rect 166626 387812 166632 387864
rect 166684 387852 166690 387864
rect 167638 387852 167644 387864
rect 166684 387824 167644 387852
rect 166684 387812 166690 387824
rect 167638 387812 167644 387824
rect 167696 387812 167702 387864
rect 220170 387812 220176 387864
rect 220228 387852 220234 387864
rect 221918 387852 221924 387864
rect 220228 387824 221924 387852
rect 220228 387812 220234 387824
rect 221918 387812 221924 387824
rect 221976 387812 221982 387864
rect 227622 387812 227628 387864
rect 227680 387852 227686 387864
rect 228358 387852 228364 387864
rect 227680 387824 228364 387852
rect 227680 387812 227686 387824
rect 228358 387812 228364 387824
rect 228416 387812 228422 387864
rect 232498 387812 232504 387864
rect 232556 387852 232562 387864
rect 234246 387852 234252 387864
rect 232556 387824 234252 387852
rect 232556 387812 232562 387824
rect 234246 387812 234252 387824
rect 234304 387812 234310 387864
rect 244918 387812 244924 387864
rect 244976 387852 244982 387864
rect 245654 387852 245660 387864
rect 244976 387824 245660 387852
rect 244976 387812 244982 387824
rect 245654 387812 245660 387824
rect 245712 387812 245718 387864
rect 252002 387812 252008 387864
rect 252060 387852 252066 387864
rect 253382 387852 253388 387864
rect 252060 387824 253388 387852
rect 252060 387812 252066 387824
rect 253382 387812 253388 387824
rect 253440 387812 253446 387864
rect 93452 387756 122834 387784
rect 93452 387744 93458 387756
rect 188338 387744 188344 387796
rect 188396 387784 188402 387796
rect 218698 387784 218704 387796
rect 188396 387756 218704 387784
rect 188396 387744 188402 387756
rect 218698 387744 218704 387756
rect 218756 387744 218762 387796
rect 225782 387744 225788 387796
rect 225840 387784 225846 387796
rect 260926 387784 260932 387796
rect 225840 387756 260932 387784
rect 225840 387744 225846 387756
rect 260926 387744 260932 387756
rect 260984 387744 260990 387796
rect 186774 387676 186780 387728
rect 186832 387716 186838 387728
rect 211614 387716 211620 387728
rect 186832 387688 211620 387716
rect 186832 387676 186838 387688
rect 211614 387676 211620 387688
rect 211672 387676 211678 387728
rect 242894 387676 242900 387728
rect 242952 387716 242958 387728
rect 266538 387716 266544 387728
rect 242952 387688 266544 387716
rect 242952 387676 242958 387688
rect 266538 387676 266544 387688
rect 266596 387716 266602 387728
rect 266722 387716 266728 387728
rect 266596 387688 266728 387716
rect 266596 387676 266602 387688
rect 266722 387676 266728 387688
rect 266780 387676 266786 387728
rect 219986 387268 219992 387320
rect 220044 387308 220050 387320
rect 225782 387308 225788 387320
rect 220044 387280 225788 387308
rect 220044 387268 220050 387280
rect 225782 387268 225788 387280
rect 225840 387268 225846 387320
rect 240962 387200 240968 387252
rect 241020 387240 241026 387252
rect 242894 387240 242900 387252
rect 241020 387212 242900 387240
rect 241020 387200 241026 387212
rect 242894 387200 242900 387212
rect 242952 387200 242958 387252
rect 100386 387064 100392 387116
rect 100444 387104 100450 387116
rect 100444 387076 109632 387104
rect 100444 387064 100450 387076
rect 69014 386996 69020 387048
rect 69072 387036 69078 387048
rect 69750 387036 69756 387048
rect 69072 387008 69756 387036
rect 69072 386996 69078 387008
rect 69750 386996 69756 387008
rect 69808 386996 69814 387048
rect 78674 386996 78680 387048
rect 78732 387036 78738 387048
rect 79502 387036 79508 387048
rect 78732 387008 79508 387036
rect 78732 386996 78738 387008
rect 79502 386996 79508 387008
rect 79560 386996 79566 387048
rect 93854 386996 93860 387048
rect 93912 387036 93918 387048
rect 94130 387036 94136 387048
rect 93912 387008 94136 387036
rect 93912 386996 93918 387008
rect 94130 386996 94136 387008
rect 94188 386996 94194 387048
rect 102134 386996 102140 387048
rect 102192 387036 102198 387048
rect 102502 387036 102508 387048
rect 102192 387008 102508 387036
rect 102192 386996 102198 387008
rect 102502 386996 102508 387008
rect 102560 386996 102566 387048
rect 109034 386996 109040 387048
rect 109092 387036 109098 387048
rect 109494 387036 109500 387048
rect 109092 387008 109500 387036
rect 109092 386996 109098 387008
rect 109494 386996 109500 387008
rect 109552 386996 109558 387048
rect 109604 387036 109632 387076
rect 110690 387064 110696 387116
rect 110748 387104 110754 387116
rect 188614 387104 188620 387116
rect 110748 387076 188620 387104
rect 110748 387064 110754 387076
rect 188614 387064 188620 387076
rect 188672 387064 188678 387116
rect 266722 387064 266728 387116
rect 266780 387104 266786 387116
rect 272242 387104 272248 387116
rect 266780 387076 272248 387104
rect 266780 387064 266786 387076
rect 272242 387064 272248 387076
rect 272300 387064 272306 387116
rect 281442 387064 281448 387116
rect 281500 387104 281506 387116
rect 582374 387104 582380 387116
rect 281500 387076 582380 387104
rect 281500 387064 281506 387076
rect 582374 387064 582380 387076
rect 582432 387064 582438 387116
rect 111058 387036 111064 387048
rect 109604 387008 111064 387036
rect 111058 386996 111064 387008
rect 111116 386996 111122 387048
rect 155218 386452 155224 386504
rect 155276 386492 155282 386504
rect 163498 386492 163504 386504
rect 155276 386464 163504 386492
rect 155276 386452 155282 386464
rect 163498 386452 163504 386464
rect 163556 386452 163562 386504
rect 84930 386316 84936 386368
rect 84988 386356 84994 386368
rect 140038 386356 140044 386368
rect 84988 386328 140044 386356
rect 84988 386316 84994 386328
rect 140038 386316 140044 386328
rect 140096 386316 140102 386368
rect 186406 386316 186412 386368
rect 186464 386356 186470 386368
rect 232498 386356 232504 386368
rect 186464 386328 232504 386356
rect 186464 386316 186470 386328
rect 232498 386316 232504 386328
rect 232556 386316 232562 386368
rect 245838 386316 245844 386368
rect 245896 386356 245902 386368
rect 246942 386356 246948 386368
rect 245896 386328 246948 386356
rect 245896 386316 245902 386328
rect 246942 386316 246948 386328
rect 247000 386356 247006 386368
rect 262858 386356 262864 386368
rect 247000 386328 262864 386356
rect 247000 386316 247006 386328
rect 262858 386316 262864 386328
rect 262916 386316 262922 386368
rect 39942 386248 39948 386300
rect 40000 386288 40006 386300
rect 88426 386288 88432 386300
rect 40000 386260 88432 386288
rect 40000 386248 40006 386260
rect 88426 386248 88432 386260
rect 88484 386288 88490 386300
rect 89254 386288 89260 386300
rect 88484 386260 89260 386288
rect 88484 386248 88490 386260
rect 89254 386248 89260 386260
rect 89312 386248 89318 386300
rect 107746 386248 107752 386300
rect 107804 386288 107810 386300
rect 134610 386288 134616 386300
rect 107804 386260 134616 386288
rect 107804 386248 107810 386260
rect 134610 386248 134616 386260
rect 134668 386288 134674 386300
rect 135162 386288 135168 386300
rect 134668 386260 135168 386288
rect 134668 386248 134674 386260
rect 135162 386248 135168 386260
rect 135220 386248 135226 386300
rect 195422 386248 195428 386300
rect 195480 386288 195486 386300
rect 197354 386288 197360 386300
rect 195480 386260 197360 386288
rect 195480 386248 195486 386260
rect 197354 386248 197360 386260
rect 197412 386248 197418 386300
rect 217318 386248 217324 386300
rect 217376 386288 217382 386300
rect 218238 386288 218244 386300
rect 217376 386260 218244 386288
rect 217376 386248 217382 386260
rect 218238 386248 218244 386260
rect 218296 386248 218302 386300
rect 239490 386248 239496 386300
rect 239548 386288 239554 386300
rect 253566 386288 253572 386300
rect 239548 386260 253572 386288
rect 239548 386248 239554 386260
rect 253566 386248 253572 386260
rect 253624 386248 253630 386300
rect 135162 385704 135168 385756
rect 135220 385744 135226 385756
rect 163498 385744 163504 385756
rect 135220 385716 163504 385744
rect 135220 385704 135226 385716
rect 163498 385704 163504 385716
rect 163556 385704 163562 385756
rect 139394 385636 139400 385688
rect 139452 385676 139458 385688
rect 189718 385676 189724 385688
rect 139452 385648 189724 385676
rect 139452 385636 139458 385648
rect 189718 385636 189724 385648
rect 189776 385636 189782 385688
rect 129734 384956 129740 385008
rect 129792 384996 129798 385008
rect 130930 384996 130936 385008
rect 129792 384968 130936 384996
rect 129792 384956 129798 384968
rect 130930 384956 130936 384968
rect 130988 384996 130994 385008
rect 230566 384996 230572 385008
rect 130988 384968 230572 384996
rect 130988 384956 130994 384968
rect 230566 384956 230572 384968
rect 230624 384996 230630 385008
rect 231486 384996 231492 385008
rect 230624 384968 231492 384996
rect 230624 384956 230630 384968
rect 231486 384956 231492 384968
rect 231544 384956 231550 385008
rect 242158 384956 242164 385008
rect 242216 384996 242222 385008
rect 271874 384996 271880 385008
rect 242216 384968 271880 384996
rect 242216 384956 242222 384968
rect 271874 384956 271880 384968
rect 271932 384956 271938 385008
rect 96890 384276 96896 384328
rect 96948 384316 96954 384328
rect 116578 384316 116584 384328
rect 96948 384288 116584 384316
rect 96948 384276 96954 384288
rect 116578 384276 116584 384288
rect 116636 384316 116642 384328
rect 129734 384316 129740 384328
rect 116636 384288 129740 384316
rect 116636 384276 116642 384288
rect 129734 384276 129740 384288
rect 129792 384276 129798 384328
rect 3510 383664 3516 383716
rect 3568 383704 3574 383716
rect 113450 383704 113456 383716
rect 3568 383676 113456 383704
rect 3568 383664 3574 383676
rect 113450 383664 113456 383676
rect 113508 383664 113514 383716
rect 228358 383664 228364 383716
rect 228416 383704 228422 383716
rect 280338 383704 280344 383716
rect 228416 383676 280344 383704
rect 228416 383664 228422 383676
rect 280338 383664 280344 383676
rect 280396 383664 280402 383716
rect 111058 383596 111064 383648
rect 111116 383636 111122 383648
rect 135898 383636 135904 383648
rect 111116 383608 135904 383636
rect 111116 383596 111122 383608
rect 135898 383596 135904 383608
rect 135956 383596 135962 383648
rect 177482 383596 177488 383648
rect 177540 383636 177546 383648
rect 256878 383636 256884 383648
rect 177540 383608 256884 383636
rect 177540 383596 177546 383608
rect 256878 383596 256884 383608
rect 256936 383596 256942 383648
rect 87046 383324 87052 383376
rect 87104 383364 87110 383376
rect 91278 383364 91284 383376
rect 87104 383336 91284 383364
rect 87104 383324 87110 383336
rect 91278 383324 91284 383336
rect 91336 383324 91342 383376
rect 135898 382984 135904 383036
rect 135956 383024 135962 383036
rect 174262 383024 174268 383036
rect 135956 382996 174268 383024
rect 135956 382984 135962 382996
rect 174262 382984 174268 382996
rect 174320 382984 174326 383036
rect 65978 382916 65984 382968
rect 66036 382956 66042 382968
rect 75178 382956 75184 382968
rect 66036 382928 75184 382956
rect 66036 382916 66042 382928
rect 75178 382916 75184 382928
rect 75236 382916 75242 382968
rect 78766 382916 78772 382968
rect 78824 382956 78830 382968
rect 97258 382956 97264 382968
rect 78824 382928 97264 382956
rect 78824 382916 78830 382928
rect 97258 382916 97264 382928
rect 97316 382916 97322 382968
rect 97442 382916 97448 382968
rect 97500 382956 97506 382968
rect 118694 382956 118700 382968
rect 97500 382928 118700 382956
rect 97500 382916 97506 382928
rect 118694 382916 118700 382928
rect 118752 382956 118758 382968
rect 231854 382956 231860 382968
rect 118752 382928 231860 382956
rect 118752 382916 118758 382928
rect 231854 382916 231860 382928
rect 231912 382956 231918 382968
rect 281718 382956 281724 382968
rect 231912 382928 281724 382956
rect 231912 382916 231918 382928
rect 281718 382916 281724 382928
rect 281776 382916 281782 382968
rect 182082 382168 182088 382220
rect 182140 382208 182146 382220
rect 229094 382208 229100 382220
rect 182140 382180 229100 382208
rect 182140 382168 182146 382180
rect 229094 382168 229100 382180
rect 229152 382168 229158 382220
rect 181438 381692 181444 381744
rect 181496 381732 181502 381744
rect 182082 381732 182088 381744
rect 181496 381704 182088 381732
rect 181496 381692 181502 381704
rect 182082 381692 182088 381704
rect 182140 381692 182146 381744
rect 102042 381556 102048 381608
rect 102100 381596 102106 381608
rect 113358 381596 113364 381608
rect 102100 381568 113364 381596
rect 102100 381556 102106 381568
rect 113358 381556 113364 381568
rect 113416 381556 113422 381608
rect 214558 381556 214564 381608
rect 214616 381596 214622 381608
rect 238754 381596 238760 381608
rect 214616 381568 238760 381596
rect 214616 381556 214622 381568
rect 238754 381556 238760 381568
rect 238812 381556 238818 381608
rect 77478 381488 77484 381540
rect 77536 381528 77542 381540
rect 161382 381528 161388 381540
rect 77536 381500 161388 381528
rect 77536 381488 77542 381500
rect 161382 381488 161388 381500
rect 161440 381528 161446 381540
rect 169018 381528 169024 381540
rect 161440 381500 169024 381528
rect 161440 381488 161446 381500
rect 169018 381488 169024 381500
rect 169076 381488 169082 381540
rect 230566 381488 230572 381540
rect 230624 381528 230630 381540
rect 277670 381528 277676 381540
rect 230624 381500 277676 381528
rect 230624 381488 230630 381500
rect 277670 381488 277676 381500
rect 277728 381488 277734 381540
rect 75270 380808 75276 380860
rect 75328 380848 75334 380860
rect 161474 380848 161480 380860
rect 75328 380820 161480 380848
rect 75328 380808 75334 380820
rect 161474 380808 161480 380820
rect 161532 380848 161538 380860
rect 162210 380848 162216 380860
rect 161532 380820 162216 380848
rect 161532 380808 161538 380820
rect 162210 380808 162216 380820
rect 162268 380808 162274 380860
rect 188614 380808 188620 380860
rect 188672 380848 188678 380860
rect 188982 380848 188988 380860
rect 188672 380820 188988 380848
rect 188672 380808 188678 380820
rect 188982 380808 188988 380820
rect 189040 380848 189046 380860
rect 250714 380848 250720 380860
rect 189040 380820 250720 380848
rect 189040 380808 189046 380820
rect 250714 380808 250720 380820
rect 250772 380808 250778 380860
rect 109126 380128 109132 380180
rect 109184 380168 109190 380180
rect 128998 380168 129004 380180
rect 109184 380140 129004 380168
rect 109184 380128 109190 380140
rect 128998 380128 129004 380140
rect 129056 380128 129062 380180
rect 141418 380128 141424 380180
rect 141476 380168 141482 380180
rect 187694 380168 187700 380180
rect 141476 380140 187700 380168
rect 141476 380128 141482 380140
rect 187694 380128 187700 380140
rect 187752 380128 187758 380180
rect 190270 380128 190276 380180
rect 190328 380168 190334 380180
rect 265066 380168 265072 380180
rect 190328 380140 265072 380168
rect 190328 380128 190334 380140
rect 265066 380128 265072 380140
rect 265124 380168 265130 380180
rect 273346 380168 273352 380180
rect 265124 380140 273352 380168
rect 265124 380128 265130 380140
rect 273346 380128 273352 380140
rect 273404 380128 273410 380180
rect 82814 379448 82820 379500
rect 82872 379488 82878 379500
rect 164878 379488 164884 379500
rect 82872 379460 164884 379488
rect 82872 379448 82878 379460
rect 164878 379448 164884 379460
rect 164936 379448 164942 379500
rect 189166 379448 189172 379500
rect 189224 379488 189230 379500
rect 273530 379488 273536 379500
rect 189224 379460 273536 379488
rect 189224 379448 189230 379460
rect 273530 379448 273536 379460
rect 273588 379448 273594 379500
rect 187694 379380 187700 379432
rect 187752 379420 187758 379432
rect 247678 379420 247684 379432
rect 187752 379392 247684 379420
rect 187752 379380 187758 379392
rect 247678 379380 247684 379392
rect 247736 379380 247742 379432
rect 273346 379244 273352 379296
rect 273404 379284 273410 379296
rect 273530 379284 273536 379296
rect 273404 379256 273536 379284
rect 273404 379244 273410 379256
rect 273530 379244 273536 379256
rect 273588 379244 273594 379296
rect 104894 378768 104900 378820
rect 104952 378808 104958 378820
rect 153930 378808 153936 378820
rect 104952 378780 153936 378808
rect 104952 378768 104958 378780
rect 153930 378768 153936 378780
rect 153988 378768 153994 378820
rect 252462 378768 252468 378820
rect 252520 378808 252526 378820
rect 266538 378808 266544 378820
rect 252520 378780 266544 378808
rect 252520 378768 252526 378780
rect 266538 378768 266544 378780
rect 266596 378768 266602 378820
rect 72510 378088 72516 378140
rect 72568 378128 72574 378140
rect 148410 378128 148416 378140
rect 72568 378100 148416 378128
rect 72568 378088 72574 378100
rect 148410 378088 148416 378100
rect 148468 378088 148474 378140
rect 161290 378088 161296 378140
rect 161348 378128 161354 378140
rect 223574 378128 223580 378140
rect 161348 378100 223580 378128
rect 161348 378088 161354 378100
rect 223574 378088 223580 378100
rect 223632 378128 223638 378140
rect 224218 378128 224224 378140
rect 223632 378100 224224 378128
rect 223632 378088 223638 378100
rect 224218 378088 224224 378100
rect 224276 378088 224282 378140
rect 236638 378088 236644 378140
rect 236696 378128 236702 378140
rect 264238 378128 264244 378140
rect 236696 378100 264244 378128
rect 236696 378088 236702 378100
rect 264238 378088 264244 378100
rect 264296 378088 264302 378140
rect 93946 377408 93952 377460
rect 94004 377448 94010 377460
rect 120718 377448 120724 377460
rect 94004 377420 120724 377448
rect 94004 377408 94010 377420
rect 120718 377408 120724 377420
rect 120776 377448 120782 377460
rect 228358 377448 228364 377460
rect 120776 377420 228364 377448
rect 120776 377408 120782 377420
rect 228358 377408 228364 377420
rect 228416 377408 228422 377460
rect 151170 376660 151176 376712
rect 151228 376700 151234 376712
rect 247126 376700 247132 376712
rect 151228 376672 247132 376700
rect 151228 376660 151234 376672
rect 247126 376660 247132 376672
rect 247184 376660 247190 376712
rect 77202 376592 77208 376644
rect 77260 376632 77266 376644
rect 154482 376632 154488 376644
rect 77260 376604 154488 376632
rect 77260 376592 77266 376604
rect 154482 376592 154488 376604
rect 154540 376592 154546 376644
rect 75914 376048 75920 376100
rect 75972 376088 75978 376100
rect 77202 376088 77208 376100
rect 75972 376060 77208 376088
rect 75972 376048 75978 376060
rect 77202 376048 77208 376060
rect 77260 376048 77266 376100
rect 46750 375980 46756 376032
rect 46808 376020 46814 376032
rect 78674 376020 78680 376032
rect 46808 375992 78680 376020
rect 46808 375980 46814 375992
rect 78674 375980 78680 375992
rect 78732 375980 78738 376032
rect 108850 375980 108856 376032
rect 108908 376020 108914 376032
rect 116026 376020 116032 376032
rect 108908 375992 116032 376020
rect 108908 375980 108914 375992
rect 116026 375980 116032 375992
rect 116084 375980 116090 376032
rect 65886 375300 65892 375352
rect 65944 375340 65950 375352
rect 171870 375340 171876 375352
rect 65944 375312 171876 375340
rect 65944 375300 65950 375312
rect 171870 375300 171876 375312
rect 171928 375340 171934 375352
rect 172054 375340 172060 375352
rect 171928 375312 172060 375340
rect 171928 375300 171934 375312
rect 172054 375300 172060 375312
rect 172112 375300 172118 375352
rect 174262 375300 174268 375352
rect 174320 375340 174326 375352
rect 235994 375340 236000 375352
rect 174320 375312 236000 375340
rect 174320 375300 174326 375312
rect 235994 375300 236000 375312
rect 236052 375340 236058 375352
rect 236638 375340 236644 375352
rect 236052 375312 236644 375340
rect 236052 375300 236058 375312
rect 236638 375300 236644 375312
rect 236696 375300 236702 375352
rect 279418 375300 279424 375352
rect 279476 375340 279482 375352
rect 281534 375340 281540 375352
rect 279476 375312 281540 375340
rect 279476 375300 279482 375312
rect 281534 375300 281540 375312
rect 281592 375300 281598 375352
rect 236638 374688 236644 374740
rect 236696 374728 236702 374740
rect 291378 374728 291384 374740
rect 236696 374700 291384 374728
rect 236696 374688 236702 374700
rect 291378 374688 291384 374700
rect 291436 374688 291442 374740
rect 88334 374620 88340 374672
rect 88392 374660 88398 374672
rect 141510 374660 141516 374672
rect 88392 374632 141516 374660
rect 88392 374620 88398 374632
rect 141510 374620 141516 374632
rect 141568 374660 141574 374672
rect 142246 374660 142252 374672
rect 141568 374632 142252 374660
rect 141568 374620 141574 374632
rect 142246 374620 142252 374632
rect 142304 374620 142310 374672
rect 148318 374620 148324 374672
rect 148376 374660 148382 374672
rect 241514 374660 241520 374672
rect 148376 374632 241520 374660
rect 148376 374620 148382 374632
rect 241514 374620 241520 374632
rect 241572 374660 241578 374672
rect 251818 374660 251824 374672
rect 241572 374632 251824 374660
rect 241572 374620 241578 374632
rect 251818 374620 251824 374632
rect 251876 374620 251882 374672
rect 163498 373940 163504 373992
rect 163556 373980 163562 373992
rect 245746 373980 245752 373992
rect 163556 373952 245752 373980
rect 163556 373940 163562 373952
rect 245746 373940 245752 373952
rect 245804 373940 245810 373992
rect 77202 373328 77208 373380
rect 77260 373368 77266 373380
rect 84286 373368 84292 373380
rect 77260 373340 84292 373368
rect 77260 373328 77266 373340
rect 84286 373328 84292 373340
rect 84344 373328 84350 373380
rect 107562 373328 107568 373380
rect 107620 373368 107626 373380
rect 115934 373368 115940 373380
rect 107620 373340 115940 373368
rect 107620 373328 107626 373340
rect 115934 373328 115940 373340
rect 115992 373328 115998 373380
rect 153930 373328 153936 373380
rect 153988 373368 153994 373380
rect 186406 373368 186412 373380
rect 153988 373340 186412 373368
rect 153988 373328 153994 373340
rect 186406 373328 186412 373340
rect 186464 373328 186470 373380
rect 244918 373328 244924 373380
rect 244976 373368 244982 373380
rect 258718 373368 258724 373380
rect 244976 373340 258724 373368
rect 244976 373328 244982 373340
rect 258718 373328 258724 373340
rect 258776 373328 258782 373380
rect 74534 373260 74540 373312
rect 74592 373300 74598 373312
rect 157334 373300 157340 373312
rect 74592 373272 157340 373300
rect 74592 373260 74598 373272
rect 157334 373260 157340 373272
rect 157392 373260 157398 373312
rect 191098 373260 191104 373312
rect 191156 373300 191162 373312
rect 203518 373300 203524 373312
rect 191156 373272 203524 373300
rect 191156 373260 191162 373272
rect 203518 373260 203524 373272
rect 203576 373260 203582 373312
rect 251910 373260 251916 373312
rect 251968 373300 251974 373312
rect 266630 373300 266636 373312
rect 251968 373272 266636 373300
rect 251968 373260 251974 373272
rect 266630 373260 266636 373272
rect 266688 373260 266694 373312
rect 117958 372580 117964 372632
rect 118016 372620 118022 372632
rect 147490 372620 147496 372632
rect 118016 372592 147496 372620
rect 118016 372580 118022 372592
rect 147490 372580 147496 372592
rect 147548 372620 147554 372632
rect 147674 372620 147680 372632
rect 147548 372592 147680 372620
rect 147548 372580 147554 372592
rect 147674 372580 147680 372592
rect 147732 372580 147738 372632
rect 245746 372580 245752 372632
rect 245804 372620 245810 372632
rect 246298 372620 246304 372632
rect 245804 372592 246304 372620
rect 245804 372580 245810 372592
rect 246298 372580 246304 372592
rect 246356 372580 246362 372632
rect 179046 372512 179052 372564
rect 179104 372552 179110 372564
rect 227714 372552 227720 372564
rect 179104 372524 227720 372552
rect 179104 372512 179110 372524
rect 227714 372512 227720 372524
rect 227772 372512 227778 372564
rect 84102 372444 84108 372496
rect 84160 372484 84166 372496
rect 180058 372484 180064 372496
rect 84160 372456 180064 372484
rect 84160 372444 84166 372456
rect 180058 372444 180064 372456
rect 180116 372444 180122 372496
rect 182910 372444 182916 372496
rect 182968 372484 182974 372496
rect 222194 372484 222200 372496
rect 182968 372456 222200 372484
rect 182968 372444 182974 372456
rect 222194 372444 222200 372456
rect 222252 372444 222258 372496
rect 48222 371832 48228 371884
rect 48280 371872 48286 371884
rect 75914 371872 75920 371884
rect 48280 371844 75920 371872
rect 48280 371832 48286 371844
rect 75914 371832 75920 371844
rect 75972 371832 75978 371884
rect 249702 371832 249708 371884
rect 249760 371872 249766 371884
rect 269390 371872 269396 371884
rect 249760 371844 269396 371872
rect 249760 371832 249766 371844
rect 269390 371832 269396 371844
rect 269448 371832 269454 371884
rect 179414 371764 179420 371816
rect 179472 371804 179478 371816
rect 180058 371804 180064 371816
rect 179472 371776 180064 371804
rect 179472 371764 179478 371776
rect 180058 371764 180064 371776
rect 180116 371764 180122 371816
rect 222194 371220 222200 371272
rect 222252 371260 222258 371272
rect 222838 371260 222844 371272
rect 222252 371232 222844 371260
rect 222252 371220 222258 371232
rect 222838 371220 222844 371232
rect 222896 371220 222902 371272
rect 227714 371220 227720 371272
rect 227772 371260 227778 371272
rect 228450 371260 228456 371272
rect 227772 371232 228456 371260
rect 227772 371220 227778 371232
rect 228450 371220 228456 371232
rect 228508 371220 228514 371272
rect 270402 371220 270408 371272
rect 270460 371260 270466 371272
rect 274910 371260 274916 371272
rect 270460 371232 274916 371260
rect 270460 371220 270466 371232
rect 274910 371220 274916 371232
rect 274968 371220 274974 371272
rect 155678 371152 155684 371204
rect 155736 371192 155742 371204
rect 240134 371192 240140 371204
rect 155736 371164 240140 371192
rect 155736 371152 155742 371164
rect 240134 371152 240140 371164
rect 240192 371192 240198 371204
rect 240870 371192 240876 371204
rect 240192 371164 240876 371192
rect 240192 371152 240198 371164
rect 240870 371152 240876 371164
rect 240928 371152 240934 371204
rect 247034 371152 247040 371204
rect 247092 371192 247098 371204
rect 248322 371192 248328 371204
rect 247092 371164 248328 371192
rect 247092 371152 247098 371164
rect 248322 371152 248328 371164
rect 248380 371192 248386 371204
rect 295426 371192 295432 371204
rect 248380 371164 295432 371192
rect 248380 371152 248386 371164
rect 295426 371152 295432 371164
rect 295484 371152 295490 371204
rect 85574 371084 85580 371136
rect 85632 371124 85638 371136
rect 160738 371124 160744 371136
rect 85632 371096 160744 371124
rect 85632 371084 85638 371096
rect 160738 371084 160744 371096
rect 160796 371084 160802 371136
rect 170398 371084 170404 371136
rect 170456 371124 170462 371136
rect 234614 371124 234620 371136
rect 170456 371096 234620 371124
rect 170456 371084 170462 371096
rect 234614 371084 234620 371096
rect 234672 371084 234678 371136
rect 234614 370472 234620 370524
rect 234672 370512 234678 370524
rect 244918 370512 244924 370524
rect 234672 370484 244924 370512
rect 234672 370472 234678 370484
rect 244918 370472 244924 370484
rect 244976 370472 244982 370524
rect 160094 370268 160100 370320
rect 160152 370308 160158 370320
rect 160738 370308 160744 370320
rect 160152 370280 160744 370308
rect 160152 370268 160158 370280
rect 160738 370268 160744 370280
rect 160796 370268 160802 370320
rect 97258 369792 97264 369844
rect 97316 369832 97322 369844
rect 129734 369832 129740 369844
rect 97316 369804 129740 369832
rect 97316 369792 97322 369804
rect 129734 369792 129740 369804
rect 129792 369792 129798 369844
rect 187694 369792 187700 369844
rect 187752 369832 187758 369844
rect 242158 369832 242164 369844
rect 187752 369804 242164 369832
rect 187752 369792 187758 369804
rect 242158 369792 242164 369804
rect 242216 369792 242222 369844
rect 164878 369724 164884 369776
rect 164936 369764 164942 369776
rect 213914 369764 213920 369776
rect 164936 369736 213920 369764
rect 164936 369724 164942 369736
rect 213914 369724 213920 369736
rect 213972 369724 213978 369776
rect 129734 369180 129740 369232
rect 129792 369220 129798 369232
rect 130378 369220 130384 369232
rect 129792 369192 130384 369220
rect 129792 369180 129798 369192
rect 130378 369180 130384 369192
rect 130436 369220 130442 369232
rect 180058 369220 180064 369232
rect 130436 369192 180064 369220
rect 130436 369180 130442 369192
rect 180058 369180 180064 369192
rect 180116 369180 180122 369232
rect 71682 369112 71688 369164
rect 71740 369152 71746 369164
rect 163958 369152 163964 369164
rect 71740 369124 163964 369152
rect 71740 369112 71746 369124
rect 163958 369112 163964 369124
rect 164016 369152 164022 369164
rect 165062 369152 165068 369164
rect 164016 369124 165068 369152
rect 164016 369112 164022 369124
rect 165062 369112 165068 369124
rect 165120 369112 165126 369164
rect 234522 369112 234528 369164
rect 234580 369152 234586 369164
rect 259454 369152 259460 369164
rect 234580 369124 259460 369152
rect 234580 369112 234586 369124
rect 259454 369112 259460 369124
rect 259512 369112 259518 369164
rect 111058 368432 111064 368484
rect 111116 368472 111122 368484
rect 113266 368472 113272 368484
rect 111116 368444 113272 368472
rect 111116 368432 111122 368444
rect 113266 368432 113272 368444
rect 113324 368472 113330 368484
rect 276106 368472 276112 368484
rect 113324 368444 276112 368472
rect 113324 368432 113330 368444
rect 276106 368432 276112 368444
rect 276164 368432 276170 368484
rect 71038 368364 71044 368416
rect 71096 368404 71102 368416
rect 169754 368404 169760 368416
rect 71096 368376 169760 368404
rect 71096 368364 71102 368376
rect 169754 368364 169760 368376
rect 169812 368364 169818 368416
rect 228358 367752 228364 367804
rect 228416 367792 228422 367804
rect 263686 367792 263692 367804
rect 228416 367764 263692 367792
rect 228416 367752 228422 367764
rect 263686 367752 263692 367764
rect 263744 367752 263750 367804
rect 67726 367004 67732 367056
rect 67784 367044 67790 367056
rect 155954 367044 155960 367056
rect 67784 367016 155960 367044
rect 67784 367004 67790 367016
rect 155954 367004 155960 367016
rect 156012 367004 156018 367056
rect 157334 367004 157340 367056
rect 157392 367044 157398 367056
rect 158438 367044 158444 367056
rect 157392 367016 158444 367044
rect 157392 367004 157398 367016
rect 158438 367004 158444 367016
rect 158496 367044 158502 367056
rect 201494 367044 201500 367056
rect 158496 367016 201500 367044
rect 158496 367004 158502 367016
rect 201494 367004 201500 367016
rect 201552 367004 201558 367056
rect 75178 366936 75184 366988
rect 75236 366976 75242 366988
rect 137462 366976 137468 366988
rect 75236 366948 137468 366976
rect 75236 366936 75242 366948
rect 137462 366936 137468 366948
rect 137520 366936 137526 366988
rect 176102 366936 176108 366988
rect 176160 366976 176166 366988
rect 176746 366976 176752 366988
rect 176160 366948 176752 366976
rect 176160 366936 176166 366948
rect 176746 366936 176752 366948
rect 176804 366936 176810 366988
rect 176746 366324 176752 366376
rect 176804 366364 176810 366376
rect 254118 366364 254124 366376
rect 176804 366336 254124 366364
rect 176804 366324 176810 366336
rect 254118 366324 254124 366336
rect 254176 366324 254182 366376
rect 73246 365644 73252 365696
rect 73304 365684 73310 365696
rect 166994 365684 167000 365696
rect 73304 365656 167000 365684
rect 73304 365644 73310 365656
rect 166994 365644 167000 365656
rect 167052 365684 167058 365696
rect 167638 365684 167644 365696
rect 167052 365656 167644 365684
rect 167052 365644 167058 365656
rect 167638 365644 167644 365656
rect 167696 365644 167702 365696
rect 186406 365644 186412 365696
rect 186464 365684 186470 365696
rect 240962 365684 240968 365696
rect 186464 365656 240968 365684
rect 186464 365644 186470 365656
rect 240962 365644 240968 365656
rect 241020 365644 241026 365696
rect 248966 365644 248972 365696
rect 249024 365684 249030 365696
rect 249794 365684 249800 365696
rect 249024 365656 249800 365684
rect 249024 365644 249030 365656
rect 249794 365644 249800 365656
rect 249852 365644 249858 365696
rect 57698 365576 57704 365628
rect 57756 365616 57762 365628
rect 144178 365616 144184 365628
rect 57756 365588 144184 365616
rect 57756 365576 57762 365588
rect 144178 365576 144184 365588
rect 144236 365576 144242 365628
rect 163958 365576 163964 365628
rect 164016 365616 164022 365628
rect 196066 365616 196072 365628
rect 164016 365588 196072 365616
rect 164016 365576 164022 365588
rect 196066 365576 196072 365588
rect 196124 365576 196130 365628
rect 196066 365168 196072 365220
rect 196124 365208 196130 365220
rect 196618 365208 196624 365220
rect 196124 365180 196624 365208
rect 196124 365168 196130 365180
rect 196618 365168 196624 365180
rect 196676 365168 196682 365220
rect 242250 364964 242256 365016
rect 242308 365004 242314 365016
rect 284478 365004 284484 365016
rect 242308 364976 284484 365004
rect 242308 364964 242314 364976
rect 284478 364964 284484 364976
rect 284536 364964 284542 365016
rect 69106 364284 69112 364336
rect 69164 364324 69170 364336
rect 171134 364324 171140 364336
rect 69164 364296 171140 364324
rect 69164 364284 69170 364296
rect 171134 364284 171140 364296
rect 171192 364324 171198 364336
rect 171962 364324 171968 364336
rect 171192 364296 171968 364324
rect 171192 364284 171198 364296
rect 171962 364284 171968 364296
rect 172020 364284 172026 364336
rect 180058 364284 180064 364336
rect 180116 364324 180122 364336
rect 180610 364324 180616 364336
rect 180116 364296 180616 364324
rect 180116 364284 180122 364296
rect 180610 364284 180616 364296
rect 180668 364324 180674 364336
rect 207014 364324 207020 364336
rect 180668 364296 207020 364324
rect 180668 364284 180674 364296
rect 207014 364284 207020 364296
rect 207072 364284 207078 364336
rect 123570 364216 123576 364268
rect 123628 364256 123634 364268
rect 226334 364256 226340 364268
rect 123628 364228 226340 364256
rect 123628 364216 123634 364228
rect 226334 364216 226340 364228
rect 226392 364216 226398 364268
rect 228450 363672 228456 363724
rect 228508 363712 228514 363724
rect 251818 363712 251824 363724
rect 228508 363684 251824 363712
rect 228508 363672 228514 363684
rect 251818 363672 251824 363684
rect 251876 363672 251882 363724
rect 260098 363672 260104 363724
rect 260156 363712 260162 363724
rect 296714 363712 296720 363724
rect 260156 363684 296720 363712
rect 260156 363672 260162 363684
rect 296714 363672 296720 363684
rect 296772 363672 296778 363724
rect 226334 363604 226340 363656
rect 226392 363644 226398 363656
rect 266630 363644 266636 363656
rect 226392 363616 266636 363644
rect 226392 363604 226398 363616
rect 266630 363604 266636 363616
rect 266688 363604 266694 363656
rect 111794 362856 111800 362908
rect 111852 362896 111858 362908
rect 112530 362896 112536 362908
rect 111852 362868 112536 362896
rect 111852 362856 111858 362868
rect 112530 362856 112536 362868
rect 112588 362896 112594 362908
rect 252002 362896 252008 362908
rect 112588 362868 252008 362896
rect 112588 362856 112594 362868
rect 252002 362856 252008 362868
rect 252060 362856 252066 362908
rect 266630 362856 266636 362908
rect 266688 362896 266694 362908
rect 293954 362896 293960 362908
rect 266688 362868 293960 362896
rect 266688 362856 266694 362868
rect 293954 362856 293960 362868
rect 294012 362856 294018 362908
rect 93854 362176 93860 362228
rect 93912 362216 93918 362228
rect 110506 362216 110512 362228
rect 93912 362188 110512 362216
rect 93912 362176 93918 362188
rect 110506 362176 110512 362188
rect 110564 362176 110570 362228
rect 151078 362176 151084 362228
rect 151136 362216 151142 362228
rect 216674 362216 216680 362228
rect 151136 362188 216680 362216
rect 151136 362176 151142 362188
rect 216674 362176 216680 362188
rect 216732 362176 216738 362228
rect 249610 361564 249616 361616
rect 249668 361604 249674 361616
rect 274726 361604 274732 361616
rect 249668 361576 274732 361604
rect 249668 361564 249674 361576
rect 274726 361564 274732 361576
rect 274784 361564 274790 361616
rect 73154 361496 73160 361548
rect 73212 361536 73218 361548
rect 140774 361536 140780 361548
rect 73212 361508 140780 361536
rect 73212 361496 73218 361508
rect 140774 361496 140780 361508
rect 140832 361496 140838 361548
rect 153838 361496 153844 361548
rect 153896 361536 153902 361548
rect 270770 361536 270776 361548
rect 153896 361508 270776 361536
rect 153896 361496 153902 361508
rect 270770 361496 270776 361508
rect 270828 361496 270834 361548
rect 140774 360816 140780 360868
rect 140832 360856 140838 360868
rect 142062 360856 142068 360868
rect 140832 360828 142068 360856
rect 140832 360816 140838 360828
rect 142062 360816 142068 360828
rect 142120 360856 142126 360868
rect 168374 360856 168380 360868
rect 142120 360828 168380 360856
rect 142120 360816 142126 360828
rect 168374 360816 168380 360828
rect 168432 360816 168438 360868
rect 69014 360136 69020 360188
rect 69072 360176 69078 360188
rect 69658 360176 69664 360188
rect 69072 360148 69664 360176
rect 69072 360136 69078 360148
rect 69658 360136 69664 360148
rect 69716 360176 69722 360188
rect 197354 360176 197360 360188
rect 69716 360148 197360 360176
rect 69716 360136 69722 360148
rect 197354 360136 197360 360148
rect 197412 360136 197418 360188
rect 168374 360068 168380 360120
rect 168432 360108 168438 360120
rect 169478 360108 169484 360120
rect 168432 360080 169484 360108
rect 168432 360068 168438 360080
rect 169478 360068 169484 360080
rect 169536 360108 169542 360120
rect 178862 360108 178868 360120
rect 169536 360080 178868 360108
rect 169536 360068 169542 360080
rect 178862 360068 178868 360080
rect 178920 360068 178926 360120
rect 206278 359456 206284 359508
rect 206336 359496 206342 359508
rect 260834 359496 260840 359508
rect 206336 359468 260840 359496
rect 206336 359456 206342 359468
rect 260834 359456 260840 359468
rect 260892 359456 260898 359508
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 36538 358748 36544 358760
rect 3384 358720 36544 358748
rect 3384 358708 3390 358720
rect 36538 358708 36544 358720
rect 36596 358708 36602 358760
rect 145650 358708 145656 358760
rect 145708 358748 145714 358760
rect 255314 358748 255320 358760
rect 145708 358720 255320 358748
rect 145708 358708 145714 358720
rect 255314 358708 255320 358720
rect 255372 358708 255378 358760
rect 100754 358028 100760 358080
rect 100812 358068 100818 358080
rect 122834 358068 122840 358080
rect 100812 358040 122840 358068
rect 100812 358028 100818 358040
rect 122834 358028 122840 358040
rect 122892 358068 122898 358080
rect 123754 358068 123760 358080
rect 122892 358040 123760 358068
rect 122892 358028 122898 358040
rect 123754 358028 123760 358040
rect 123812 358028 123818 358080
rect 123754 357416 123760 357468
rect 123812 357456 123818 357468
rect 239398 357456 239404 357468
rect 123812 357428 239404 357456
rect 123812 357416 123818 357428
rect 239398 357416 239404 357428
rect 239456 357416 239462 357468
rect 196618 356736 196624 356788
rect 196676 356776 196682 356788
rect 240134 356776 240140 356788
rect 196676 356748 240140 356776
rect 196676 356736 196682 356748
rect 240134 356736 240140 356748
rect 240192 356736 240198 356788
rect 128998 356668 129004 356720
rect 129056 356708 129062 356720
rect 168374 356708 168380 356720
rect 129056 356680 168380 356708
rect 129056 356668 129062 356680
rect 168374 356668 168380 356680
rect 168432 356708 168438 356720
rect 214650 356708 214656 356720
rect 168432 356680 214656 356708
rect 168432 356668 168438 356680
rect 214650 356668 214656 356680
rect 214708 356668 214714 356720
rect 229002 356668 229008 356720
rect 229060 356708 229066 356720
rect 256786 356708 256792 356720
rect 229060 356680 256792 356708
rect 229060 356668 229066 356680
rect 256786 356668 256792 356680
rect 256844 356668 256850 356720
rect 75178 355988 75184 356040
rect 75236 356028 75242 356040
rect 75822 356028 75828 356040
rect 75236 356000 75828 356028
rect 75236 355988 75242 356000
rect 75822 355988 75828 356000
rect 75880 356028 75886 356040
rect 191098 356028 191104 356040
rect 75880 356000 191104 356028
rect 75880 355988 75886 356000
rect 191098 355988 191104 356000
rect 191156 355988 191162 356040
rect 102226 355920 102232 355972
rect 102284 355960 102290 355972
rect 103330 355960 103336 355972
rect 102284 355932 103336 355960
rect 102284 355920 102290 355932
rect 103330 355920 103336 355932
rect 103388 355960 103394 355972
rect 214558 355960 214564 355972
rect 103388 355932 214564 355960
rect 103388 355920 103394 355932
rect 214558 355920 214564 355932
rect 214616 355920 214622 355972
rect 213178 355376 213184 355428
rect 213236 355416 213242 355428
rect 258166 355416 258172 355428
rect 213236 355388 258172 355416
rect 213236 355376 213242 355388
rect 258166 355376 258172 355388
rect 258224 355376 258230 355428
rect 214558 355308 214564 355360
rect 214616 355348 214622 355360
rect 269206 355348 269212 355360
rect 214616 355320 269212 355348
rect 214616 355308 214622 355320
rect 269206 355308 269212 355320
rect 269264 355308 269270 355360
rect 102134 354628 102140 354680
rect 102192 354668 102198 354680
rect 239490 354668 239496 354680
rect 102192 354640 239496 354668
rect 102192 354628 102198 354640
rect 239490 354628 239496 354640
rect 239548 354628 239554 354680
rect 244182 354016 244188 354068
rect 244240 354056 244246 354068
rect 262398 354056 262404 354068
rect 244240 354028 262404 354056
rect 244240 354016 244246 354028
rect 262398 354016 262404 354028
rect 262456 354016 262462 354068
rect 213822 353948 213828 354000
rect 213880 353988 213886 354000
rect 259546 353988 259552 354000
rect 213880 353960 259552 353988
rect 213880 353948 213886 353960
rect 259546 353948 259552 353960
rect 259604 353948 259610 354000
rect 153838 353268 153844 353320
rect 153896 353308 153902 353320
rect 198734 353308 198740 353320
rect 153896 353280 198740 353308
rect 153896 353268 153902 353280
rect 198734 353268 198740 353280
rect 198792 353268 198798 353320
rect 147490 353200 147496 353252
rect 147548 353240 147554 353252
rect 217318 353240 217324 353252
rect 147548 353212 217324 353240
rect 147548 353200 147554 353212
rect 217318 353200 217324 353212
rect 217376 353200 217382 353252
rect 108850 352520 108856 352572
rect 108908 352560 108914 352572
rect 280430 352560 280436 352572
rect 108908 352532 280436 352560
rect 108908 352520 108914 352532
rect 280430 352520 280436 352532
rect 280488 352520 280494 352572
rect 108390 351908 108396 351960
rect 108448 351948 108454 351960
rect 108850 351948 108856 351960
rect 108448 351920 108856 351948
rect 108448 351908 108454 351920
rect 108850 351908 108856 351920
rect 108908 351908 108914 351960
rect 162578 351160 162584 351212
rect 162636 351200 162642 351212
rect 194594 351200 194600 351212
rect 162636 351172 194600 351200
rect 162636 351160 162642 351172
rect 194594 351160 194600 351172
rect 194652 351160 194658 351212
rect 216582 351160 216588 351212
rect 216640 351200 216646 351212
rect 238110 351200 238116 351212
rect 216640 351172 238116 351200
rect 216640 351160 216646 351172
rect 238110 351160 238116 351172
rect 238168 351160 238174 351212
rect 84194 350548 84200 350600
rect 84252 350588 84258 350600
rect 270678 350588 270684 350600
rect 84252 350560 270684 350588
rect 84252 350548 84258 350560
rect 270678 350548 270684 350560
rect 270736 350588 270742 350600
rect 270954 350588 270960 350600
rect 270736 350560 270960 350588
rect 270736 350548 270742 350560
rect 270954 350548 270960 350560
rect 271012 350548 271018 350600
rect 88242 350480 88248 350532
rect 88300 350520 88306 350532
rect 220078 350520 220084 350532
rect 88300 350492 220084 350520
rect 88300 350480 88306 350492
rect 220078 350480 220084 350492
rect 220136 350480 220142 350532
rect 207658 349800 207664 349852
rect 207716 349840 207722 349852
rect 235258 349840 235264 349852
rect 207716 349812 235264 349840
rect 207716 349800 207722 349812
rect 235258 349800 235264 349812
rect 235316 349800 235322 349852
rect 146938 348440 146944 348492
rect 146996 348480 147002 348492
rect 188890 348480 188896 348492
rect 146996 348452 188896 348480
rect 146996 348440 147002 348452
rect 188890 348440 188896 348452
rect 188948 348480 188954 348492
rect 206370 348480 206376 348492
rect 188948 348452 206376 348480
rect 188948 348440 188954 348452
rect 206370 348440 206376 348452
rect 206428 348440 206434 348492
rect 209130 348440 209136 348492
rect 209188 348480 209194 348492
rect 233878 348480 233884 348492
rect 209188 348452 233884 348480
rect 209188 348440 209194 348452
rect 233878 348440 233884 348452
rect 233936 348440 233942 348492
rect 278958 348412 278964 348424
rect 113146 348384 278964 348412
rect 106918 348304 106924 348356
rect 106976 348344 106982 348356
rect 107562 348344 107568 348356
rect 106976 348316 107568 348344
rect 106976 348304 106982 348316
rect 107562 348304 107568 348316
rect 107620 348344 107626 348356
rect 113146 348344 113174 348384
rect 278958 348372 278964 348384
rect 279016 348372 279022 348424
rect 107620 348316 113174 348344
rect 107620 348304 107626 348316
rect 234430 347012 234436 347064
rect 234488 347052 234494 347064
rect 267734 347052 267740 347064
rect 234488 347024 267740 347052
rect 234488 347012 234494 347024
rect 267734 347012 267740 347024
rect 267792 347012 267798 347064
rect 134610 346468 134616 346520
rect 134668 346508 134674 346520
rect 214558 346508 214564 346520
rect 134668 346480 214564 346508
rect 134668 346468 134674 346480
rect 214558 346468 214564 346480
rect 214616 346468 214622 346520
rect 147122 346400 147128 346452
rect 147180 346440 147186 346452
rect 289998 346440 290004 346452
rect 147180 346412 290004 346440
rect 147180 346400 147186 346412
rect 289998 346400 290004 346412
rect 290056 346400 290062 346452
rect 71958 345584 71964 345636
rect 72016 345624 72022 345636
rect 73062 345624 73068 345636
rect 72016 345596 73068 345624
rect 72016 345584 72022 345596
rect 73062 345584 73068 345596
rect 73120 345584 73126 345636
rect 122098 345108 122104 345160
rect 122156 345148 122162 345160
rect 217410 345148 217416 345160
rect 122156 345120 217416 345148
rect 122156 345108 122162 345120
rect 217410 345108 217416 345120
rect 217468 345108 217474 345160
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 35158 345080 35164 345092
rect 3384 345052 35164 345080
rect 3384 345040 3390 345052
rect 35158 345040 35164 345052
rect 35216 345040 35222 345092
rect 73062 345040 73068 345092
rect 73120 345080 73126 345092
rect 292666 345080 292672 345092
rect 73120 345052 292672 345080
rect 73120 345040 73126 345052
rect 292666 345040 292672 345052
rect 292724 345040 292730 345092
rect 245010 344360 245016 344412
rect 245068 344400 245074 344412
rect 253934 344400 253940 344412
rect 245068 344372 253940 344400
rect 245068 344360 245074 344372
rect 253934 344360 253940 344372
rect 253992 344360 253998 344412
rect 15194 344292 15200 344344
rect 15252 344332 15258 344344
rect 150342 344332 150348 344344
rect 15252 344304 150348 344332
rect 15252 344292 15258 344304
rect 150342 344292 150348 344304
rect 150400 344332 150406 344344
rect 197354 344332 197360 344344
rect 150400 344304 197360 344332
rect 150400 344292 150406 344304
rect 197354 344292 197360 344304
rect 197412 344292 197418 344344
rect 197998 344292 198004 344344
rect 198056 344332 198062 344344
rect 236638 344332 236644 344344
rect 198056 344304 236644 344332
rect 198056 344292 198062 344304
rect 236638 344292 236644 344304
rect 236696 344292 236702 344344
rect 250438 344292 250444 344344
rect 250496 344332 250502 344344
rect 267734 344332 267740 344344
rect 250496 344304 267740 344332
rect 250496 344292 250502 344304
rect 267734 344292 267740 344304
rect 267792 344292 267798 344344
rect 44174 342864 44180 342916
rect 44232 342904 44238 342916
rect 189166 342904 189172 342916
rect 44232 342876 189172 342904
rect 44232 342864 44238 342876
rect 189166 342864 189172 342876
rect 189224 342864 189230 342916
rect 206462 342864 206468 342916
rect 206520 342904 206526 342916
rect 253934 342904 253940 342916
rect 206520 342876 253940 342904
rect 206520 342864 206526 342876
rect 253934 342864 253940 342876
rect 253992 342864 253998 342916
rect 124858 342524 124864 342576
rect 124916 342564 124922 342576
rect 125502 342564 125508 342576
rect 124916 342536 125508 342564
rect 124916 342524 124922 342536
rect 125502 342524 125508 342536
rect 125560 342524 125566 342576
rect 125502 342252 125508 342304
rect 125560 342292 125566 342304
rect 269390 342292 269396 342304
rect 125560 342264 269396 342292
rect 125560 342252 125566 342264
rect 269390 342252 269396 342264
rect 269448 342252 269454 342304
rect 177298 341504 177304 341556
rect 177356 341544 177362 341556
rect 185026 341544 185032 341556
rect 177356 341516 185032 341544
rect 177356 341504 177362 341516
rect 185026 341504 185032 341516
rect 185084 341504 185090 341556
rect 67450 340892 67456 340944
rect 67508 340932 67514 340944
rect 295610 340932 295616 340944
rect 67508 340904 295616 340932
rect 67508 340892 67514 340904
rect 295610 340892 295616 340904
rect 295668 340892 295674 340944
rect 215938 340144 215944 340196
rect 215996 340184 216002 340196
rect 243078 340184 243084 340196
rect 215996 340156 243084 340184
rect 215996 340144 216002 340156
rect 243078 340144 243084 340156
rect 243136 340144 243142 340196
rect 116762 339532 116768 339584
rect 116820 339572 116826 339584
rect 183554 339572 183560 339584
rect 116820 339544 183560 339572
rect 116820 339532 116826 339544
rect 183554 339532 183560 339544
rect 183612 339572 183618 339584
rect 184290 339572 184296 339584
rect 183612 339544 184296 339572
rect 183612 339532 183618 339544
rect 184290 339532 184296 339544
rect 184348 339532 184354 339584
rect 82722 339464 82728 339516
rect 82780 339504 82786 339516
rect 220078 339504 220084 339516
rect 82780 339476 220084 339504
rect 82780 339464 82786 339476
rect 220078 339464 220084 339476
rect 220136 339464 220142 339516
rect 183278 339396 183284 339448
rect 183336 339436 183342 339448
rect 186314 339436 186320 339448
rect 183336 339408 186320 339436
rect 183336 339396 183342 339408
rect 186314 339396 186320 339408
rect 186372 339396 186378 339448
rect 234338 339396 234344 339448
rect 234396 339436 234402 339448
rect 234798 339436 234804 339448
rect 234396 339408 234804 339436
rect 234396 339396 234402 339408
rect 234798 339396 234804 339408
rect 234856 339396 234862 339448
rect 187602 338784 187608 338836
rect 187660 338824 187666 338836
rect 251910 338824 251916 338836
rect 187660 338796 251916 338824
rect 187660 338784 187666 338796
rect 251910 338784 251916 338796
rect 251968 338784 251974 338836
rect 155218 338716 155224 338768
rect 155276 338756 155282 338768
rect 234798 338756 234804 338768
rect 155276 338728 234804 338756
rect 155276 338716 155282 338728
rect 234798 338716 234804 338728
rect 234856 338716 234862 338768
rect 178034 337424 178040 337476
rect 178092 337464 178098 337476
rect 237374 337464 237380 337476
rect 178092 337436 237380 337464
rect 178092 337424 178098 337436
rect 237374 337424 237380 337436
rect 237432 337424 237438 337476
rect 252002 337424 252008 337476
rect 252060 337464 252066 337476
rect 261018 337464 261024 337476
rect 252060 337436 261024 337464
rect 252060 337424 252066 337436
rect 261018 337424 261024 337436
rect 261076 337424 261082 337476
rect 217318 337356 217324 337408
rect 217376 337396 217382 337408
rect 294138 337396 294144 337408
rect 217376 337368 294144 337396
rect 217376 337356 217382 337368
rect 294138 337356 294144 337368
rect 294196 337356 294202 337408
rect 41414 336812 41420 336864
rect 41472 336852 41478 336864
rect 178034 336852 178040 336864
rect 41472 336824 178040 336852
rect 41472 336812 41478 336824
rect 178034 336812 178040 336824
rect 178092 336812 178098 336864
rect 178126 336744 178132 336796
rect 178184 336784 178190 336796
rect 212626 336784 212632 336796
rect 178184 336756 212632 336784
rect 178184 336744 178190 336756
rect 212626 336744 212632 336756
rect 212684 336744 212690 336796
rect 186130 335996 186136 336048
rect 186188 336036 186194 336048
rect 244458 336036 244464 336048
rect 186188 336008 244464 336036
rect 186188 335996 186194 336008
rect 244458 335996 244464 336008
rect 244516 335996 244522 336048
rect 137370 335316 137376 335368
rect 137428 335356 137434 335368
rect 245010 335356 245016 335368
rect 137428 335328 245016 335356
rect 137428 335316 137434 335328
rect 245010 335316 245016 335328
rect 245068 335316 245074 335368
rect 178586 334024 178592 334076
rect 178644 334064 178650 334076
rect 230566 334064 230572 334076
rect 178644 334036 230572 334064
rect 178644 334024 178650 334036
rect 230566 334024 230572 334036
rect 230624 334024 230630 334076
rect 178862 333956 178868 334008
rect 178920 333996 178926 334008
rect 242250 333996 242256 334008
rect 178920 333968 242256 333996
rect 178920 333956 178926 333968
rect 242250 333956 242256 333968
rect 242308 333956 242314 334008
rect 210418 333208 210424 333260
rect 210476 333248 210482 333260
rect 274634 333248 274640 333260
rect 210476 333220 274640 333248
rect 210476 333208 210482 333220
rect 274634 333208 274640 333220
rect 274692 333208 274698 333260
rect 169018 332664 169024 332716
rect 169076 332704 169082 332716
rect 200206 332704 200212 332716
rect 169076 332676 200212 332704
rect 169076 332664 169082 332676
rect 200206 332664 200212 332676
rect 200264 332664 200270 332716
rect 141602 332596 141608 332648
rect 141660 332636 141666 332648
rect 247126 332636 247132 332648
rect 141660 332608 247132 332636
rect 141660 332596 141666 332608
rect 247126 332596 247132 332608
rect 247184 332636 247190 332648
rect 247678 332636 247684 332648
rect 247184 332608 247684 332636
rect 247184 332596 247190 332608
rect 247678 332596 247684 332608
rect 247736 332596 247742 332648
rect 219342 331916 219348 331968
rect 219400 331956 219406 331968
rect 260098 331956 260104 331968
rect 219400 331928 260104 331956
rect 219400 331916 219406 331928
rect 260098 331916 260104 331928
rect 260156 331916 260162 331968
rect 141694 331848 141700 331900
rect 141752 331888 141758 331900
rect 183370 331888 183376 331900
rect 141752 331860 183376 331888
rect 141752 331848 141758 331860
rect 183370 331848 183376 331860
rect 183428 331888 183434 331900
rect 235994 331888 236000 331900
rect 183428 331860 236000 331888
rect 183428 331848 183434 331860
rect 235994 331848 236000 331860
rect 236052 331848 236058 331900
rect 163498 331236 163504 331288
rect 163556 331276 163562 331288
rect 191834 331276 191840 331288
rect 163556 331248 191840 331276
rect 163556 331236 163562 331248
rect 191834 331236 191840 331248
rect 191892 331276 191898 331288
rect 193030 331276 193036 331288
rect 191892 331248 193036 331276
rect 191892 331236 191898 331248
rect 193030 331236 193036 331248
rect 193088 331236 193094 331288
rect 127618 330488 127624 330540
rect 127676 330528 127682 330540
rect 204162 330528 204168 330540
rect 127676 330500 204168 330528
rect 127676 330488 127682 330500
rect 204162 330488 204168 330500
rect 204220 330488 204226 330540
rect 246298 330488 246304 330540
rect 246356 330528 246362 330540
rect 259454 330528 259460 330540
rect 246356 330500 259460 330528
rect 246356 330488 246362 330500
rect 259454 330488 259460 330500
rect 259512 330488 259518 330540
rect 264882 330488 264888 330540
rect 264940 330528 264946 330540
rect 272150 330528 272156 330540
rect 264940 330500 272156 330528
rect 264940 330488 264946 330500
rect 272150 330488 272156 330500
rect 272208 330488 272214 330540
rect 205726 329876 205732 329928
rect 205784 329916 205790 329928
rect 245654 329916 245660 329928
rect 205784 329888 245660 329916
rect 205784 329876 205790 329888
rect 245654 329876 245660 329888
rect 245712 329876 245718 329928
rect 166350 329808 166356 329860
rect 166408 329848 166414 329860
rect 166718 329848 166724 329860
rect 166408 329820 166724 329848
rect 166408 329808 166414 329820
rect 166718 329808 166724 329820
rect 166776 329848 166782 329860
rect 258166 329848 258172 329860
rect 166776 329820 258172 329848
rect 166776 329808 166782 329820
rect 258166 329808 258172 329820
rect 258224 329808 258230 329860
rect 153010 329740 153016 329792
rect 153068 329780 153074 329792
rect 157334 329780 157340 329792
rect 153068 329752 157340 329780
rect 153068 329740 153074 329752
rect 157334 329740 157340 329752
rect 157392 329740 157398 329792
rect 8294 329060 8300 329112
rect 8352 329100 8358 329112
rect 153194 329100 153200 329112
rect 8352 329072 153200 329100
rect 8352 329060 8358 329072
rect 153194 329060 153200 329072
rect 153252 329060 153258 329112
rect 186222 329060 186228 329112
rect 186280 329100 186286 329112
rect 187510 329100 187516 329112
rect 186280 329072 187516 329100
rect 186280 329060 186286 329072
rect 187510 329060 187516 329072
rect 187568 329100 187574 329112
rect 205726 329100 205732 329112
rect 187568 329072 205732 329100
rect 187568 329060 187574 329072
rect 205726 329060 205732 329072
rect 205784 329060 205790 329112
rect 233878 329060 233884 329112
rect 233936 329100 233942 329112
rect 253198 329100 253204 329112
rect 233936 329072 253204 329100
rect 233936 329060 233942 329072
rect 253198 329060 253204 329072
rect 253256 329060 253262 329112
rect 157334 328448 157340 328500
rect 157392 328488 157398 328500
rect 243170 328488 243176 328500
rect 157392 328460 243176 328488
rect 157392 328448 157398 328460
rect 243170 328448 243176 328460
rect 243228 328448 243234 328500
rect 193030 328176 193036 328228
rect 193088 328216 193094 328228
rect 195974 328216 195980 328228
rect 193088 328188 195980 328216
rect 193088 328176 193094 328188
rect 195974 328176 195980 328188
rect 196032 328176 196038 328228
rect 96706 327700 96712 327752
rect 96764 327740 96770 327752
rect 249886 327740 249892 327752
rect 96764 327712 249892 327740
rect 96764 327700 96770 327712
rect 249886 327700 249892 327712
rect 249944 327700 249950 327752
rect 241514 326408 241520 326460
rect 241572 326448 241578 326460
rect 242342 326448 242348 326460
rect 241572 326420 242348 326448
rect 241572 326408 241578 326420
rect 242342 326408 242348 326420
rect 242400 326408 242406 326460
rect 251818 326408 251824 326460
rect 251876 326448 251882 326460
rect 260834 326448 260840 326460
rect 251876 326420 260840 326448
rect 251876 326408 251882 326420
rect 260834 326408 260840 326420
rect 260892 326408 260898 326460
rect 33134 326340 33140 326392
rect 33192 326380 33198 326392
rect 154022 326380 154028 326392
rect 33192 326352 154028 326380
rect 33192 326340 33198 326352
rect 154022 326340 154028 326352
rect 154080 326340 154086 326392
rect 184290 326340 184296 326392
rect 184348 326380 184354 326392
rect 251910 326380 251916 326392
rect 184348 326352 251916 326380
rect 184348 326340 184354 326352
rect 251910 326340 251916 326352
rect 251968 326340 251974 326392
rect 155310 325660 155316 325712
rect 155368 325700 155374 325712
rect 241514 325700 241520 325712
rect 155368 325672 241520 325700
rect 155368 325660 155374 325672
rect 241514 325660 241520 325672
rect 241572 325660 241578 325712
rect 280522 325660 280528 325712
rect 280580 325700 280586 325712
rect 580902 325700 580908 325712
rect 280580 325672 580908 325700
rect 280580 325660 280586 325672
rect 580902 325660 580908 325672
rect 580960 325660 580966 325712
rect 153930 324980 153936 325032
rect 153988 325020 153994 325032
rect 215294 325020 215300 325032
rect 153988 324992 215300 325020
rect 153988 324980 153994 324992
rect 215294 324980 215300 324992
rect 215352 325020 215358 325032
rect 256878 325020 256884 325032
rect 215352 324992 256884 325020
rect 215352 324980 215358 324992
rect 256878 324980 256884 324992
rect 256936 324980 256942 325032
rect 88978 324912 88984 324964
rect 89036 324952 89042 324964
rect 166350 324952 166356 324964
rect 89036 324924 166356 324952
rect 89036 324912 89042 324924
rect 166350 324912 166356 324924
rect 166408 324912 166414 324964
rect 193122 324912 193128 324964
rect 193180 324952 193186 324964
rect 255498 324952 255504 324964
rect 193180 324924 255504 324952
rect 193180 324912 193186 324924
rect 255498 324912 255504 324924
rect 255556 324912 255562 324964
rect 151078 323620 151084 323672
rect 151136 323660 151142 323672
rect 162118 323660 162124 323672
rect 151136 323632 162124 323660
rect 151136 323620 151142 323632
rect 162118 323620 162124 323632
rect 162176 323620 162182 323672
rect 176010 323620 176016 323672
rect 176068 323660 176074 323672
rect 204254 323660 204260 323672
rect 176068 323632 204260 323660
rect 176068 323620 176074 323632
rect 204254 323620 204260 323632
rect 204312 323620 204318 323672
rect 211798 323620 211804 323672
rect 211856 323660 211862 323672
rect 246390 323660 246396 323672
rect 211856 323632 246396 323660
rect 211856 323620 211862 323632
rect 246390 323620 246396 323632
rect 246448 323620 246454 323672
rect 152550 323552 152556 323604
rect 152608 323592 152614 323604
rect 183462 323592 183468 323604
rect 152608 323564 183468 323592
rect 152608 323552 152614 323564
rect 183462 323552 183468 323564
rect 183520 323592 183526 323604
rect 209774 323592 209780 323604
rect 183520 323564 209780 323592
rect 183520 323552 183526 323564
rect 209774 323552 209780 323564
rect 209832 323552 209838 323604
rect 220078 323552 220084 323604
rect 220136 323592 220142 323604
rect 262214 323592 262220 323604
rect 220136 323564 262220 323592
rect 220136 323552 220142 323564
rect 262214 323552 262220 323564
rect 262272 323552 262278 323604
rect 115198 321648 115204 321700
rect 115256 321688 115262 321700
rect 185670 321688 185676 321700
rect 115256 321660 185676 321688
rect 115256 321648 115262 321660
rect 185670 321648 185676 321660
rect 185728 321648 185734 321700
rect 155862 321580 155868 321632
rect 155920 321620 155926 321632
rect 158806 321620 158812 321632
rect 155920 321592 158812 321620
rect 155920 321580 155926 321592
rect 158806 321580 158812 321592
rect 158864 321620 158870 321632
rect 263778 321620 263784 321632
rect 158864 321592 263784 321620
rect 158864 321580 158870 321592
rect 263778 321580 263784 321592
rect 263836 321580 263842 321632
rect 126882 321512 126888 321564
rect 126940 321552 126946 321564
rect 281534 321552 281540 321564
rect 126940 321524 281540 321552
rect 126940 321512 126946 321524
rect 281534 321512 281540 321524
rect 281592 321512 281598 321564
rect 281534 321308 281540 321360
rect 281592 321348 281598 321360
rect 281810 321348 281816 321360
rect 281592 321320 281816 321348
rect 281592 321308 281598 321320
rect 281810 321308 281816 321320
rect 281868 321308 281874 321360
rect 104250 320832 104256 320884
rect 104308 320872 104314 320884
rect 125686 320872 125692 320884
rect 104308 320844 125692 320872
rect 104308 320832 104314 320844
rect 125686 320832 125692 320844
rect 125744 320872 125750 320884
rect 126882 320872 126888 320884
rect 125744 320844 126888 320872
rect 125744 320832 125750 320844
rect 126882 320832 126888 320844
rect 126940 320832 126946 320884
rect 106182 320152 106188 320204
rect 106240 320192 106246 320204
rect 261018 320192 261024 320204
rect 106240 320164 261024 320192
rect 106240 320152 106246 320164
rect 261018 320152 261024 320164
rect 261076 320152 261082 320204
rect 251818 320084 251824 320136
rect 251876 320124 251882 320136
rect 252002 320124 252008 320136
rect 251876 320096 252008 320124
rect 251876 320084 251882 320096
rect 252002 320084 252008 320096
rect 252060 320084 252066 320136
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 15838 319444 15844 319456
rect 4120 319416 15844 319444
rect 4120 319404 4126 319416
rect 15838 319404 15844 319416
rect 15896 319404 15902 319456
rect 188338 319404 188344 319456
rect 188396 319444 188402 319456
rect 267918 319444 267924 319456
rect 188396 319416 267924 319444
rect 188396 319404 188402 319416
rect 267918 319404 267924 319416
rect 267976 319404 267982 319456
rect 181898 319064 181904 319116
rect 181956 319104 181962 319116
rect 187050 319104 187056 319116
rect 181956 319076 187056 319104
rect 181956 319064 181962 319076
rect 187050 319064 187056 319076
rect 187108 319064 187114 319116
rect 162118 318792 162124 318844
rect 162176 318832 162182 318844
rect 251818 318832 251824 318844
rect 162176 318804 251824 318832
rect 162176 318792 162182 318804
rect 251818 318792 251824 318804
rect 251876 318792 251882 318844
rect 182818 318044 182824 318096
rect 182876 318084 182882 318096
rect 185026 318084 185032 318096
rect 182876 318056 185032 318084
rect 182876 318044 182882 318056
rect 185026 318044 185032 318056
rect 185084 318084 185090 318096
rect 233878 318084 233884 318096
rect 185084 318056 233884 318084
rect 185084 318044 185090 318056
rect 233878 318044 233884 318056
rect 233936 318044 233942 318096
rect 240870 318044 240876 318096
rect 240928 318084 240934 318096
rect 256786 318084 256792 318096
rect 240928 318056 256792 318084
rect 240928 318044 240934 318056
rect 256786 318044 256792 318056
rect 256844 318044 256850 318096
rect 149974 317500 149980 317552
rect 150032 317540 150038 317552
rect 182174 317540 182180 317552
rect 150032 317512 182180 317540
rect 150032 317500 150038 317512
rect 182174 317500 182180 317512
rect 182232 317500 182238 317552
rect 178678 317432 178684 317484
rect 178736 317472 178742 317484
rect 236638 317472 236644 317484
rect 178736 317444 236644 317472
rect 178736 317432 178742 317444
rect 236638 317432 236644 317444
rect 236696 317432 236702 317484
rect 246298 317432 246304 317484
rect 246356 317472 246362 317484
rect 250990 317472 250996 317484
rect 246356 317444 250996 317472
rect 246356 317432 246362 317444
rect 250990 317432 250996 317444
rect 251048 317432 251054 317484
rect 75270 317364 75276 317416
rect 75328 317404 75334 317416
rect 81434 317404 81440 317416
rect 75328 317376 81440 317404
rect 75328 317364 75334 317376
rect 81434 317364 81440 317376
rect 81492 317364 81498 317416
rect 151630 316752 151636 316804
rect 151688 316792 151694 316804
rect 169662 316792 169668 316804
rect 151688 316764 169668 316792
rect 151688 316752 151694 316764
rect 169662 316752 169668 316764
rect 169720 316752 169726 316804
rect 32398 316684 32404 316736
rect 32456 316724 32462 316736
rect 159358 316724 159364 316736
rect 32456 316696 159364 316724
rect 32456 316684 32462 316696
rect 159358 316684 159364 316696
rect 159416 316724 159422 316736
rect 263594 316724 263600 316736
rect 159416 316696 263600 316724
rect 159416 316684 159422 316696
rect 263594 316684 263600 316696
rect 263652 316684 263658 316736
rect 169662 316004 169668 316056
rect 169720 316044 169726 316056
rect 264974 316044 264980 316056
rect 169720 316016 264980 316044
rect 169720 316004 169726 316016
rect 264974 316004 264980 316016
rect 265032 316004 265038 316056
rect 89530 315256 89536 315308
rect 89588 315296 89594 315308
rect 99466 315296 99472 315308
rect 89588 315268 99472 315296
rect 89588 315256 89594 315268
rect 99466 315256 99472 315268
rect 99524 315256 99530 315308
rect 256694 315256 256700 315308
rect 256752 315296 256758 315308
rect 257430 315296 257436 315308
rect 256752 315268 257436 315296
rect 256752 315256 256758 315268
rect 257430 315256 257436 315268
rect 257488 315296 257494 315308
rect 295518 315296 295524 315308
rect 257488 315268 295524 315296
rect 257488 315256 257494 315268
rect 295518 315256 295524 315268
rect 295576 315256 295582 315308
rect 160738 314712 160744 314764
rect 160796 314752 160802 314764
rect 256694 314752 256700 314764
rect 160796 314724 256700 314752
rect 160796 314712 160802 314724
rect 256694 314712 256700 314724
rect 256752 314712 256758 314764
rect 60642 314644 60648 314696
rect 60700 314684 60706 314696
rect 263686 314684 263692 314696
rect 60700 314656 263692 314684
rect 60700 314644 60706 314656
rect 263686 314644 263692 314656
rect 263744 314644 263750 314696
rect 182174 313964 182180 314016
rect 182232 314004 182238 314016
rect 247770 314004 247776 314016
rect 182232 313976 247776 314004
rect 182232 313964 182238 313976
rect 247770 313964 247776 313976
rect 247828 313964 247834 314016
rect 129090 313896 129096 313948
rect 129148 313936 129154 313948
rect 260926 313936 260932 313948
rect 129148 313908 260932 313936
rect 129148 313896 129154 313908
rect 260926 313896 260932 313908
rect 260984 313896 260990 313948
rect 104434 313284 104440 313336
rect 104492 313324 104498 313336
rect 124858 313324 124864 313336
rect 104492 313296 124864 313324
rect 104492 313284 104498 313296
rect 124858 313284 124864 313296
rect 124916 313324 124922 313336
rect 129090 313324 129096 313336
rect 124916 313296 129096 313324
rect 124916 313284 124922 313296
rect 129090 313284 129096 313296
rect 129148 313284 129154 313336
rect 249610 313284 249616 313336
rect 249668 313324 249674 313336
rect 296714 313324 296720 313336
rect 249668 313296 296720 313324
rect 249668 313284 249674 313296
rect 296714 313284 296720 313296
rect 296772 313284 296778 313336
rect 104342 312604 104348 312656
rect 104400 312644 104406 312656
rect 115198 312644 115204 312656
rect 104400 312616 115204 312644
rect 104400 312604 104406 312616
rect 115198 312604 115204 312616
rect 115256 312604 115262 312656
rect 242158 312604 242164 312656
rect 242216 312644 242222 312656
rect 252738 312644 252744 312656
rect 242216 312616 252744 312644
rect 242216 312604 242222 312616
rect 252738 312604 252744 312616
rect 252796 312604 252802 312656
rect 73798 312536 73804 312588
rect 73856 312576 73862 312588
rect 80238 312576 80244 312588
rect 73856 312548 80244 312576
rect 73856 312536 73862 312548
rect 80238 312536 80244 312548
rect 80296 312536 80302 312588
rect 108206 312536 108212 312588
rect 108264 312576 108270 312588
rect 142154 312576 142160 312588
rect 108264 312548 142160 312576
rect 108264 312536 108270 312548
rect 142154 312536 142160 312548
rect 142212 312576 142218 312588
rect 262490 312576 262496 312588
rect 142212 312548 262496 312576
rect 142212 312536 142218 312548
rect 262490 312536 262496 312548
rect 262548 312536 262554 312588
rect 148410 311856 148416 311908
rect 148468 311896 148474 311908
rect 217410 311896 217416 311908
rect 148468 311868 217416 311896
rect 148468 311856 148474 311868
rect 217410 311856 217416 311868
rect 217468 311856 217474 311908
rect 149790 311352 149796 311364
rect 142126 311324 149796 311352
rect 126330 311176 126336 311228
rect 126388 311216 126394 311228
rect 142126 311216 142154 311324
rect 149790 311312 149796 311324
rect 149848 311312 149854 311364
rect 126388 311188 142154 311216
rect 126388 311176 126394 311188
rect 82906 311108 82912 311160
rect 82964 311148 82970 311160
rect 147122 311148 147128 311160
rect 82964 311120 147128 311148
rect 82964 311108 82970 311120
rect 147122 311108 147128 311120
rect 147180 311108 147186 311160
rect 164970 311108 164976 311160
rect 165028 311148 165034 311160
rect 173158 311148 173164 311160
rect 165028 311120 173164 311148
rect 165028 311108 165034 311120
rect 173158 311108 173164 311120
rect 173216 311148 173222 311160
rect 218054 311148 218060 311160
rect 173216 311120 218060 311148
rect 173216 311108 173222 311120
rect 218054 311108 218060 311120
rect 218112 311108 218118 311160
rect 239398 311108 239404 311160
rect 239456 311148 239462 311160
rect 255406 311148 255412 311160
rect 239456 311120 255412 311148
rect 239456 311108 239462 311120
rect 255406 311108 255412 311120
rect 255464 311108 255470 311160
rect 155402 310496 155408 310548
rect 155460 310536 155466 310548
rect 276290 310536 276296 310548
rect 155460 310508 276296 310536
rect 155460 310496 155466 310508
rect 276290 310496 276296 310508
rect 276348 310496 276354 310548
rect 97258 309816 97264 309868
rect 97316 309856 97322 309868
rect 108206 309856 108212 309868
rect 97316 309828 108212 309856
rect 97316 309816 97322 309828
rect 108206 309816 108212 309828
rect 108264 309816 108270 309868
rect 163774 309816 163780 309868
rect 163832 309856 163838 309868
rect 257338 309856 257344 309868
rect 163832 309828 257344 309856
rect 163832 309816 163838 309828
rect 257338 309816 257344 309828
rect 257396 309856 257402 309868
rect 259546 309856 259552 309868
rect 257396 309828 259552 309856
rect 257396 309816 257402 309828
rect 259546 309816 259552 309828
rect 259604 309816 259610 309868
rect 61746 309748 61752 309800
rect 61804 309788 61810 309800
rect 166442 309788 166448 309800
rect 61804 309760 166448 309788
rect 61804 309748 61810 309760
rect 166442 309748 166448 309760
rect 166500 309748 166506 309800
rect 230474 309748 230480 309800
rect 230532 309788 230538 309800
rect 252646 309788 252652 309800
rect 230532 309760 252652 309788
rect 230532 309748 230538 309760
rect 252646 309748 252652 309760
rect 252704 309748 252710 309800
rect 189074 309136 189080 309188
rect 189132 309176 189138 309188
rect 190362 309176 190368 309188
rect 189132 309148 190368 309176
rect 189132 309136 189138 309148
rect 190362 309136 190368 309148
rect 190420 309176 190426 309188
rect 218698 309176 218704 309188
rect 190420 309148 218704 309176
rect 190420 309136 190426 309148
rect 218698 309136 218704 309148
rect 218756 309136 218762 309188
rect 178586 308456 178592 308508
rect 178644 308496 178650 308508
rect 189074 308496 189080 308508
rect 178644 308468 189080 308496
rect 178644 308456 178650 308468
rect 189074 308456 189080 308468
rect 189132 308456 189138 308508
rect 99190 308388 99196 308440
rect 99248 308428 99254 308440
rect 125502 308428 125508 308440
rect 99248 308400 125508 308428
rect 99248 308388 99254 308400
rect 125502 308388 125508 308400
rect 125560 308428 125566 308440
rect 131114 308428 131120 308440
rect 125560 308400 131120 308428
rect 125560 308388 125566 308400
rect 131114 308388 131120 308400
rect 131172 308388 131178 308440
rect 151170 308388 151176 308440
rect 151228 308428 151234 308440
rect 157242 308428 157248 308440
rect 151228 308400 157248 308428
rect 151228 308388 151234 308400
rect 157242 308388 157248 308400
rect 157300 308428 157306 308440
rect 207566 308428 207572 308440
rect 157300 308400 207572 308428
rect 157300 308388 157306 308400
rect 207566 308388 207572 308400
rect 207624 308388 207630 308440
rect 224862 308388 224868 308440
rect 224920 308428 224926 308440
rect 255590 308428 255596 308440
rect 224920 308400 255596 308428
rect 224920 308388 224926 308400
rect 255590 308388 255596 308400
rect 255648 308388 255654 308440
rect 189718 307776 189724 307828
rect 189776 307816 189782 307828
rect 225966 307816 225972 307828
rect 189776 307788 225972 307816
rect 189776 307776 189782 307788
rect 225966 307776 225972 307788
rect 226024 307776 226030 307828
rect 239490 307776 239496 307828
rect 239548 307816 239554 307828
rect 241422 307816 241428 307828
rect 239548 307788 241428 307816
rect 239548 307776 239554 307788
rect 241422 307776 241428 307788
rect 241480 307776 241486 307828
rect 138014 307708 138020 307760
rect 138072 307748 138078 307760
rect 149974 307748 149980 307760
rect 138072 307720 149980 307748
rect 138072 307708 138078 307720
rect 149974 307708 149980 307720
rect 150032 307708 150038 307760
rect 173710 307708 173716 307760
rect 173768 307748 173774 307760
rect 175274 307748 175280 307760
rect 173768 307720 175280 307748
rect 173768 307708 173774 307720
rect 175274 307708 175280 307720
rect 175332 307708 175338 307760
rect 196250 307708 196256 307760
rect 196308 307748 196314 307760
rect 196710 307748 196716 307760
rect 196308 307720 196716 307748
rect 196308 307708 196314 307720
rect 196710 307708 196716 307720
rect 196768 307708 196774 307760
rect 176746 307204 176752 307216
rect 161446 307176 176752 307204
rect 71130 307096 71136 307148
rect 71188 307136 71194 307148
rect 77386 307136 77392 307148
rect 71188 307108 77392 307136
rect 71188 307096 71194 307108
rect 77386 307096 77392 307108
rect 77444 307096 77450 307148
rect 122190 307096 122196 307148
rect 122248 307136 122254 307148
rect 122248 307108 142154 307136
rect 122248 307096 122254 307108
rect 74626 307028 74632 307080
rect 74684 307068 74690 307080
rect 138014 307068 138020 307080
rect 74684 307040 138020 307068
rect 74684 307028 74690 307040
rect 138014 307028 138020 307040
rect 138072 307028 138078 307080
rect 142126 307068 142154 307108
rect 145558 307068 145564 307080
rect 142126 307040 145564 307068
rect 145558 307028 145564 307040
rect 145616 307068 145622 307080
rect 161446 307068 161474 307176
rect 176746 307164 176752 307176
rect 176804 307164 176810 307216
rect 176010 307096 176016 307148
rect 176068 307136 176074 307148
rect 176470 307136 176476 307148
rect 176068 307108 176476 307136
rect 176068 307096 176074 307108
rect 176470 307096 176476 307108
rect 176528 307096 176534 307148
rect 145616 307040 161474 307068
rect 145616 307028 145622 307040
rect 176746 307028 176752 307080
rect 176804 307068 176810 307080
rect 196250 307068 196256 307080
rect 176804 307040 196256 307068
rect 176804 307028 176810 307040
rect 196250 307028 196256 307040
rect 196308 307028 196314 307080
rect 236638 307028 236644 307080
rect 236696 307068 236702 307080
rect 267826 307068 267832 307080
rect 236696 307040 267832 307068
rect 236696 307028 236702 307040
rect 267826 307028 267832 307040
rect 267884 307028 267890 307080
rect 169478 306552 169484 306604
rect 169536 306592 169542 306604
rect 172514 306592 172520 306604
rect 169536 306564 172520 306592
rect 169536 306552 169542 306564
rect 172514 306552 172520 306564
rect 172572 306552 172578 306604
rect 176010 306348 176016 306400
rect 176068 306388 176074 306400
rect 259730 306388 259736 306400
rect 176068 306360 259736 306388
rect 176068 306348 176074 306360
rect 259730 306348 259736 306360
rect 259788 306348 259794 306400
rect 67358 305600 67364 305652
rect 67416 305640 67422 305652
rect 88978 305640 88984 305652
rect 67416 305612 88984 305640
rect 67416 305600 67422 305612
rect 88978 305600 88984 305612
rect 89036 305600 89042 305652
rect 91186 305600 91192 305652
rect 91244 305640 91250 305652
rect 104434 305640 104440 305652
rect 91244 305612 104440 305640
rect 91244 305600 91250 305612
rect 104434 305600 104440 305612
rect 104492 305600 104498 305652
rect 109034 305600 109040 305652
rect 109092 305640 109098 305652
rect 118786 305640 118792 305652
rect 109092 305612 118792 305640
rect 109092 305600 109098 305612
rect 118786 305600 118792 305612
rect 118844 305600 118850 305652
rect 119338 305600 119344 305652
rect 119396 305640 119402 305652
rect 144270 305640 144276 305652
rect 119396 305612 144276 305640
rect 119396 305600 119402 305612
rect 144270 305600 144276 305612
rect 144328 305600 144334 305652
rect 185670 305600 185676 305652
rect 185728 305640 185734 305652
rect 193858 305640 193864 305652
rect 185728 305612 193864 305640
rect 185728 305600 185734 305612
rect 193858 305600 193864 305612
rect 193916 305600 193922 305652
rect 206370 305600 206376 305652
rect 206428 305640 206434 305652
rect 215386 305640 215392 305652
rect 206428 305612 215392 305640
rect 206428 305600 206434 305612
rect 215386 305600 215392 305612
rect 215444 305600 215450 305652
rect 4062 305124 4068 305176
rect 4120 305164 4126 305176
rect 7558 305164 7564 305176
rect 4120 305136 7564 305164
rect 4120 305124 4126 305136
rect 7558 305124 7564 305136
rect 7616 305124 7622 305176
rect 193582 305056 193588 305108
rect 193640 305096 193646 305108
rect 228358 305096 228364 305108
rect 193640 305068 228364 305096
rect 193640 305056 193646 305068
rect 228358 305056 228364 305068
rect 228416 305056 228422 305108
rect 252462 305056 252468 305108
rect 252520 305096 252526 305108
rect 258074 305096 258080 305108
rect 252520 305068 258080 305096
rect 252520 305056 252526 305068
rect 258074 305056 258080 305068
rect 258132 305096 258138 305108
rect 258718 305096 258724 305108
rect 258132 305068 258724 305096
rect 258132 305056 258138 305068
rect 258718 305056 258724 305068
rect 258776 305056 258782 305108
rect 80054 304988 80060 305040
rect 80112 305028 80118 305040
rect 109034 305028 109040 305040
rect 80112 305000 109040 305028
rect 80112 304988 80118 305000
rect 109034 304988 109040 305000
rect 109092 304988 109098 305040
rect 144822 304988 144828 305040
rect 144880 305028 144886 305040
rect 197446 305028 197452 305040
rect 144880 305000 197452 305028
rect 144880 304988 144886 305000
rect 197446 304988 197452 305000
rect 197504 304988 197510 305040
rect 253382 304988 253388 305040
rect 253440 305028 253446 305040
rect 284478 305028 284484 305040
rect 253440 305000 284484 305028
rect 253440 304988 253446 305000
rect 284478 304988 284484 305000
rect 284536 304988 284542 305040
rect 223390 304920 223396 304972
rect 223448 304960 223454 304972
rect 227622 304960 227628 304972
rect 223448 304932 227628 304960
rect 223448 304920 223454 304932
rect 227622 304920 227628 304932
rect 227680 304960 227686 304972
rect 229830 304960 229836 304972
rect 227680 304932 229836 304960
rect 227680 304920 227686 304932
rect 229830 304920 229836 304932
rect 229888 304920 229894 304972
rect 251910 304784 251916 304836
rect 251968 304824 251974 304836
rect 258258 304824 258264 304836
rect 251968 304796 258264 304824
rect 251968 304784 251974 304796
rect 258258 304784 258264 304796
rect 258316 304784 258322 304836
rect 232222 304580 232228 304632
rect 232280 304620 232286 304632
rect 240778 304620 240784 304632
rect 232280 304592 240784 304620
rect 232280 304580 232286 304592
rect 240778 304580 240784 304592
rect 240836 304580 240842 304632
rect 123570 304308 123576 304360
rect 123628 304348 123634 304360
rect 144178 304348 144184 304360
rect 123628 304320 144184 304348
rect 123628 304308 123634 304320
rect 144178 304308 144184 304320
rect 144236 304308 144242 304360
rect 218422 304308 218428 304360
rect 218480 304348 218486 304360
rect 219342 304348 219348 304360
rect 218480 304320 219348 304348
rect 218480 304308 218486 304320
rect 219342 304308 219348 304320
rect 219400 304308 219406 304360
rect 242434 304308 242440 304360
rect 242492 304348 242498 304360
rect 252462 304348 252468 304360
rect 242492 304320 252468 304348
rect 242492 304308 242498 304320
rect 252462 304308 252468 304320
rect 252520 304308 252526 304360
rect 96614 304240 96620 304292
rect 96672 304280 96678 304292
rect 147214 304280 147220 304292
rect 96672 304252 147220 304280
rect 96672 304240 96678 304252
rect 147214 304240 147220 304252
rect 147272 304240 147278 304292
rect 181438 304240 181444 304292
rect 181496 304280 181502 304292
rect 229002 304280 229008 304292
rect 181496 304252 229008 304280
rect 181496 304240 181502 304252
rect 229002 304240 229008 304252
rect 229060 304240 229066 304292
rect 247770 304240 247776 304292
rect 247828 304280 247834 304292
rect 258350 304280 258356 304292
rect 247828 304252 258356 304280
rect 247828 304240 247834 304252
rect 258350 304240 258356 304252
rect 258408 304240 258414 304292
rect 262674 304240 262680 304292
rect 262732 304280 262738 304292
rect 298186 304280 298192 304292
rect 262732 304252 298192 304280
rect 262732 304240 262738 304252
rect 298186 304240 298192 304252
rect 298244 304240 298250 304292
rect 232498 303696 232504 303748
rect 232556 303736 232562 303748
rect 233970 303736 233976 303748
rect 232556 303708 233976 303736
rect 232556 303696 232562 303708
rect 233970 303696 233976 303708
rect 234028 303696 234034 303748
rect 148318 303628 148324 303680
rect 148376 303668 148382 303680
rect 213178 303668 213184 303680
rect 148376 303640 213184 303668
rect 148376 303628 148382 303640
rect 213178 303628 213184 303640
rect 213236 303628 213242 303680
rect 214558 303628 214564 303680
rect 214616 303668 214622 303680
rect 217226 303668 217232 303680
rect 214616 303640 217232 303668
rect 214616 303628 214622 303640
rect 217226 303628 217232 303640
rect 217284 303628 217290 303680
rect 220906 303628 220912 303680
rect 220964 303668 220970 303680
rect 221734 303668 221740 303680
rect 220964 303640 221740 303668
rect 220964 303628 220970 303640
rect 221734 303628 221740 303640
rect 221792 303628 221798 303680
rect 223574 303628 223580 303680
rect 223632 303668 223638 303680
rect 224126 303668 224132 303680
rect 223632 303640 224132 303668
rect 223632 303628 223638 303640
rect 224126 303628 224132 303640
rect 224184 303628 224190 303680
rect 225046 303628 225052 303680
rect 225104 303668 225110 303680
rect 226242 303668 226248 303680
rect 225104 303640 226248 303668
rect 225104 303628 225110 303640
rect 226242 303628 226248 303640
rect 226300 303628 226306 303680
rect 230566 303628 230572 303680
rect 230624 303668 230630 303680
rect 231302 303668 231308 303680
rect 230624 303640 231308 303668
rect 230624 303628 230630 303640
rect 231302 303628 231308 303640
rect 231360 303628 231366 303680
rect 233878 303628 233884 303680
rect 233936 303668 233942 303680
rect 234614 303668 234620 303680
rect 233936 303640 234620 303668
rect 233936 303628 233942 303640
rect 234614 303628 234620 303640
rect 234672 303628 234678 303680
rect 237374 303628 237380 303680
rect 237432 303668 237438 303680
rect 237926 303668 237932 303680
rect 237432 303640 237932 303668
rect 237432 303628 237438 303640
rect 237926 303628 237932 303640
rect 237984 303628 237990 303680
rect 242250 303628 242256 303680
rect 242308 303668 242314 303680
rect 244182 303668 244188 303680
rect 242308 303640 244188 303668
rect 242308 303628 242314 303640
rect 244182 303628 244188 303640
rect 244240 303628 244246 303680
rect 248690 303628 248696 303680
rect 248748 303668 248754 303680
rect 249334 303668 249340 303680
rect 248748 303640 249340 303668
rect 248748 303628 248754 303640
rect 249334 303628 249340 303640
rect 249392 303628 249398 303680
rect 201586 303560 201592 303612
rect 201644 303560 201650 303612
rect 202874 303560 202880 303612
rect 202932 303600 202938 303612
rect 203702 303600 203708 303612
rect 202932 303572 203708 303600
rect 202932 303560 202938 303572
rect 203702 303560 203708 303572
rect 203760 303560 203766 303612
rect 204254 303560 204260 303612
rect 204312 303600 204318 303612
rect 204806 303600 204812 303612
rect 204312 303572 204812 303600
rect 204312 303560 204318 303572
rect 204806 303560 204812 303572
rect 204864 303560 204870 303612
rect 201604 303408 201632 303560
rect 201586 303356 201592 303408
rect 201644 303356 201650 303408
rect 216582 303356 216588 303408
rect 216640 303396 216646 303408
rect 218974 303396 218980 303408
rect 216640 303368 218980 303396
rect 216640 303356 216646 303368
rect 218974 303356 218980 303368
rect 219032 303356 219038 303408
rect 233418 303152 233424 303204
rect 233476 303192 233482 303204
rect 234430 303192 234436 303204
rect 233476 303164 234436 303192
rect 233476 303152 233482 303164
rect 234430 303152 234436 303164
rect 234488 303152 234494 303204
rect 121454 302880 121460 302932
rect 121512 302920 121518 302932
rect 216582 302920 216588 302932
rect 121512 302892 216588 302920
rect 121512 302880 121518 302892
rect 216582 302880 216588 302892
rect 216640 302880 216646 302932
rect 240594 302268 240600 302320
rect 240652 302308 240658 302320
rect 262306 302308 262312 302320
rect 240652 302280 262312 302308
rect 240652 302268 240658 302280
rect 262306 302268 262312 302280
rect 262364 302308 262370 302320
rect 262674 302308 262680 302320
rect 262364 302280 262680 302308
rect 262364 302268 262370 302280
rect 262674 302268 262680 302280
rect 262732 302268 262738 302320
rect 73062 302200 73068 302252
rect 73120 302240 73126 302252
rect 164970 302240 164976 302252
rect 73120 302212 164976 302240
rect 73120 302200 73126 302212
rect 164970 302200 164976 302212
rect 165028 302200 165034 302252
rect 187050 302200 187056 302252
rect 187108 302240 187114 302252
rect 233418 302240 233424 302252
rect 187108 302212 233424 302240
rect 187108 302200 187114 302212
rect 233418 302200 233424 302212
rect 233476 302200 233482 302252
rect 268102 302240 268108 302252
rect 243556 302212 268108 302240
rect 231118 302132 231124 302184
rect 231176 302172 231182 302184
rect 243556 302172 243584 302212
rect 268102 302200 268108 302212
rect 268160 302200 268166 302252
rect 231176 302144 243584 302172
rect 231176 302132 231182 302144
rect 258718 302132 258724 302184
rect 258776 302172 258782 302184
rect 266354 302172 266360 302184
rect 258776 302144 266360 302172
rect 258776 302132 258782 302144
rect 266354 302132 266360 302144
rect 266412 302132 266418 302184
rect 86218 301520 86224 301572
rect 86276 301560 86282 301572
rect 129182 301560 129188 301572
rect 86276 301532 129188 301560
rect 86276 301520 86282 301532
rect 129182 301520 129188 301532
rect 129240 301520 129246 301572
rect 242342 301520 242348 301572
rect 242400 301560 242406 301572
rect 242400 301532 244274 301560
rect 242400 301520 242406 301532
rect 34514 301452 34520 301504
rect 34572 301492 34578 301504
rect 179322 301492 179328 301504
rect 34572 301464 179328 301492
rect 34572 301452 34578 301464
rect 179322 301452 179328 301464
rect 179380 301452 179386 301504
rect 244246 301492 244274 301532
rect 254118 301492 254124 301504
rect 244246 301464 254124 301492
rect 254118 301452 254124 301464
rect 254176 301452 254182 301504
rect 244366 301384 244372 301436
rect 244424 301424 244430 301436
rect 245102 301424 245108 301436
rect 244424 301396 245108 301424
rect 244424 301384 244430 301396
rect 245102 301384 245108 301396
rect 245160 301384 245166 301436
rect 215662 301084 215668 301096
rect 200086 301056 215668 301084
rect 193674 300908 193680 300960
rect 193732 300948 193738 300960
rect 197630 300948 197636 300960
rect 193732 300920 197636 300948
rect 193732 300908 193738 300920
rect 197630 300908 197636 300920
rect 197688 300908 197694 300960
rect 166258 300840 166264 300892
rect 166316 300880 166322 300892
rect 200086 300880 200114 301056
rect 215662 301044 215668 301056
rect 215720 301044 215726 301096
rect 211062 300976 211068 301028
rect 211120 300976 211126 301028
rect 166316 300852 200114 300880
rect 166316 300840 166322 300852
rect 156598 300772 156604 300824
rect 156656 300812 156662 300824
rect 160830 300812 160836 300824
rect 156656 300784 160836 300812
rect 156656 300772 156662 300784
rect 160830 300772 160836 300784
rect 160888 300812 160894 300824
rect 191098 300812 191104 300824
rect 160888 300784 191104 300812
rect 160888 300772 160894 300784
rect 191098 300772 191104 300784
rect 191156 300772 191162 300824
rect 129182 300160 129188 300212
rect 129240 300200 129246 300212
rect 141694 300200 141700 300212
rect 129240 300172 141700 300200
rect 129240 300160 129246 300172
rect 141694 300160 141700 300172
rect 141752 300160 141758 300212
rect 190914 300160 190920 300212
rect 190972 300200 190978 300212
rect 211080 300200 211108 300976
rect 216858 300908 216864 300960
rect 216916 300948 216922 300960
rect 227714 300948 227720 300960
rect 216916 300920 227720 300948
rect 216916 300908 216922 300920
rect 227714 300908 227720 300920
rect 227772 300908 227778 300960
rect 249242 300908 249248 300960
rect 249300 300948 249306 300960
rect 258718 300948 258724 300960
rect 249300 300920 258724 300948
rect 249300 300908 249306 300920
rect 258718 300908 258724 300920
rect 258776 300908 258782 300960
rect 190972 300172 211108 300200
rect 190972 300160 190978 300172
rect 255314 300160 255320 300212
rect 255372 300200 255378 300212
rect 274634 300200 274640 300212
rect 255372 300172 274640 300200
rect 255372 300160 255378 300172
rect 274634 300160 274640 300172
rect 274692 300160 274698 300212
rect 140222 300092 140228 300144
rect 140280 300132 140286 300144
rect 193582 300132 193588 300144
rect 140280 300104 193588 300132
rect 140280 300092 140286 300104
rect 193582 300092 193588 300104
rect 193640 300092 193646 300144
rect 252462 300092 252468 300144
rect 252520 300132 252526 300144
rect 254026 300132 254032 300144
rect 252520 300104 254032 300132
rect 252520 300092 252526 300104
rect 254026 300092 254032 300104
rect 254084 300092 254090 300144
rect 258718 300092 258724 300144
rect 258776 300132 258782 300144
rect 282914 300132 282920 300144
rect 258776 300104 282920 300132
rect 258776 300092 258782 300104
rect 282914 300092 282920 300104
rect 282972 300092 282978 300144
rect 253014 299412 253020 299464
rect 253072 299452 253078 299464
rect 272058 299452 272064 299464
rect 253072 299424 272064 299452
rect 253072 299412 253078 299424
rect 272058 299412 272064 299424
rect 272116 299412 272122 299464
rect 159542 298800 159548 298852
rect 159600 298840 159606 298852
rect 188982 298840 188988 298852
rect 159600 298812 188988 298840
rect 159600 298800 159606 298812
rect 188982 298800 188988 298812
rect 189040 298840 189046 298852
rect 191742 298840 191748 298852
rect 189040 298812 191748 298840
rect 189040 298800 189046 298812
rect 191742 298800 191748 298812
rect 191800 298800 191806 298852
rect 138750 298732 138756 298784
rect 138808 298772 138814 298784
rect 187694 298772 187700 298784
rect 138808 298744 187700 298772
rect 138808 298732 138814 298744
rect 187694 298732 187700 298744
rect 187752 298732 187758 298784
rect 256602 298120 256608 298172
rect 256660 298160 256666 298172
rect 261478 298160 261484 298172
rect 256660 298132 261484 298160
rect 256660 298120 256666 298132
rect 261478 298120 261484 298132
rect 261536 298120 261542 298172
rect 304258 298120 304264 298172
rect 304316 298160 304322 298172
rect 580166 298160 580172 298172
rect 304316 298132 580172 298160
rect 304316 298120 304322 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 168466 298052 168472 298104
rect 168524 298092 168530 298104
rect 189718 298092 189724 298104
rect 168524 298064 189724 298092
rect 168524 298052 168530 298064
rect 189718 298052 189724 298064
rect 189776 298052 189782 298104
rect 122926 297372 122932 297424
rect 122984 297412 122990 297424
rect 132402 297412 132408 297424
rect 122984 297384 132408 297412
rect 122984 297372 122990 297384
rect 132402 297372 132408 297384
rect 132460 297412 132466 297424
rect 184842 297412 184848 297424
rect 132460 297384 184848 297412
rect 132460 297372 132466 297384
rect 184842 297372 184848 297384
rect 184900 297412 184906 297424
rect 191742 297412 191748 297424
rect 184900 297384 191748 297412
rect 184900 297372 184906 297384
rect 191742 297372 191748 297384
rect 191800 297372 191806 297424
rect 88426 297168 88432 297220
rect 88484 297208 88490 297220
rect 89530 297208 89536 297220
rect 88484 297180 89536 297208
rect 88484 297168 88490 297180
rect 89530 297168 89536 297180
rect 89588 297168 89594 297220
rect 89530 296692 89536 296744
rect 89588 296732 89594 296744
rect 115382 296732 115388 296744
rect 89588 296704 115388 296732
rect 89588 296692 89594 296704
rect 115382 296692 115388 296704
rect 115440 296692 115446 296744
rect 255314 296692 255320 296744
rect 255372 296732 255378 296744
rect 267918 296732 267924 296744
rect 255372 296704 267924 296732
rect 255372 296692 255378 296704
rect 267918 296692 267924 296704
rect 267976 296692 267982 296744
rect 256602 296012 256608 296064
rect 256660 296052 256666 296064
rect 272058 296052 272064 296064
rect 256660 296024 272064 296052
rect 256660 296012 256666 296024
rect 272058 296012 272064 296024
rect 272116 296012 272122 296064
rect 161934 295944 161940 295996
rect 161992 295984 161998 295996
rect 175182 295984 175188 295996
rect 161992 295956 175188 295984
rect 161992 295944 161998 295956
rect 175182 295944 175188 295956
rect 175240 295984 175246 295996
rect 185670 295984 185676 295996
rect 175240 295956 185676 295984
rect 175240 295944 175246 295956
rect 185670 295944 185676 295956
rect 185728 295944 185734 295996
rect 258534 295944 258540 295996
rect 258592 295984 258598 295996
rect 288710 295984 288716 295996
rect 258592 295956 288716 295984
rect 258592 295944 258598 295956
rect 288710 295944 288716 295956
rect 288768 295944 288774 295996
rect 165522 295332 165528 295384
rect 165580 295372 165586 295384
rect 168374 295372 168380 295384
rect 165580 295344 168380 295372
rect 165580 295332 165586 295344
rect 168374 295332 168380 295344
rect 168432 295332 168438 295384
rect 256602 295264 256608 295316
rect 256660 295304 256666 295316
rect 267734 295304 267740 295316
rect 256660 295276 267740 295304
rect 256660 295264 256666 295276
rect 267734 295264 267740 295276
rect 267792 295304 267798 295316
rect 274818 295304 274824 295316
rect 267792 295276 274824 295304
rect 267792 295264 267798 295276
rect 274818 295264 274824 295276
rect 274876 295264 274882 295316
rect 155954 294652 155960 294704
rect 156012 294692 156018 294704
rect 156598 294692 156604 294704
rect 156012 294664 156604 294692
rect 156012 294652 156018 294664
rect 156598 294652 156604 294664
rect 156656 294652 156662 294704
rect 137462 294584 137468 294636
rect 137520 294624 137526 294636
rect 144730 294624 144736 294636
rect 137520 294596 144736 294624
rect 137520 294584 137526 294596
rect 144730 294584 144736 294596
rect 144788 294624 144794 294636
rect 175182 294624 175188 294636
rect 144788 294596 175188 294624
rect 144788 294584 144794 294596
rect 175182 294584 175188 294596
rect 175240 294584 175246 294636
rect 69658 293972 69664 294024
rect 69716 294012 69722 294024
rect 155954 294012 155960 294024
rect 69716 293984 155960 294012
rect 69716 293972 69722 293984
rect 155954 293972 155960 293984
rect 156012 293972 156018 294024
rect 175182 293972 175188 294024
rect 175240 294012 175246 294024
rect 191742 294012 191748 294024
rect 175240 293984 191748 294012
rect 175240 293972 175246 293984
rect 191742 293972 191748 293984
rect 191800 293972 191806 294024
rect 256326 293972 256332 294024
rect 256384 294012 256390 294024
rect 289998 294012 290004 294024
rect 256384 293984 290004 294012
rect 256384 293972 256390 293984
rect 289998 293972 290004 293984
rect 290056 293972 290062 294024
rect 92566 293904 92572 293956
rect 92624 293944 92630 293956
rect 93762 293944 93768 293956
rect 92624 293916 93768 293944
rect 92624 293904 92630 293916
rect 93762 293904 93768 293916
rect 93820 293944 93826 293956
rect 122926 293944 122932 293956
rect 93820 293916 122932 293944
rect 93820 293904 93826 293916
rect 122926 293904 122932 293916
rect 122984 293904 122990 293956
rect 261570 293904 261576 293956
rect 261628 293944 261634 293956
rect 262214 293944 262220 293956
rect 261628 293916 262220 293944
rect 261628 293904 261634 293916
rect 262214 293904 262220 293916
rect 262272 293904 262278 293956
rect 302326 293944 302332 293956
rect 263566 293916 302332 293944
rect 261478 293836 261484 293888
rect 261536 293876 261542 293888
rect 263566 293876 263594 293916
rect 302326 293904 302332 293916
rect 302384 293904 302390 293956
rect 261536 293848 263594 293876
rect 261536 293836 261542 293848
rect 255958 293224 255964 293276
rect 256016 293264 256022 293276
rect 258810 293264 258816 293276
rect 256016 293236 258816 293264
rect 256016 293224 256022 293236
rect 258810 293224 258816 293236
rect 258868 293224 258874 293276
rect 256142 293088 256148 293140
rect 256200 293128 256206 293140
rect 260742 293128 260748 293140
rect 256200 293100 260748 293128
rect 256200 293088 256206 293100
rect 260742 293088 260748 293100
rect 260800 293088 260806 293140
rect 168374 292612 168380 292664
rect 168432 292652 168438 292664
rect 169110 292652 169116 292664
rect 168432 292624 169116 292652
rect 168432 292612 168438 292624
rect 169110 292612 169116 292624
rect 169168 292652 169174 292664
rect 191558 292652 191564 292664
rect 169168 292624 191564 292652
rect 169168 292612 169174 292624
rect 191558 292612 191564 292624
rect 191616 292612 191622 292664
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 22830 292584 22836 292596
rect 3568 292556 22836 292584
rect 3568 292544 3574 292556
rect 22830 292544 22836 292556
rect 22888 292544 22894 292596
rect 84562 292544 84568 292596
rect 84620 292584 84626 292596
rect 177850 292584 177856 292596
rect 84620 292556 177856 292584
rect 84620 292544 84626 292556
rect 177850 292544 177856 292556
rect 177908 292544 177914 292596
rect 184750 292544 184756 292596
rect 184808 292584 184814 292596
rect 188706 292584 188712 292596
rect 184808 292556 188712 292584
rect 184808 292544 184814 292556
rect 188706 292544 188712 292556
rect 188764 292544 188770 292596
rect 99282 292476 99288 292528
rect 99340 292516 99346 292528
rect 157150 292516 157156 292528
rect 99340 292488 157156 292516
rect 99340 292476 99346 292488
rect 157150 292476 157156 292488
rect 157208 292516 157214 292528
rect 168374 292516 168380 292528
rect 157208 292488 168380 292516
rect 157208 292476 157214 292488
rect 168374 292476 168380 292488
rect 168432 292476 168438 292528
rect 255958 292136 255964 292188
rect 256016 292176 256022 292188
rect 256878 292176 256884 292188
rect 256016 292148 256884 292176
rect 256016 292136 256022 292148
rect 256878 292136 256884 292148
rect 256936 292176 256942 292188
rect 258626 292176 258632 292188
rect 256936 292148 258632 292176
rect 256936 292136 256942 292148
rect 258626 292136 258632 292148
rect 258684 292136 258690 292188
rect 177850 292068 177856 292120
rect 177908 292108 177914 292120
rect 178862 292108 178868 292120
rect 177908 292080 178868 292108
rect 177908 292068 177914 292080
rect 178862 292068 178868 292080
rect 178920 292068 178926 292120
rect 178954 291864 178960 291916
rect 179012 291904 179018 291916
rect 188338 291904 188344 291916
rect 179012 291876 188344 291904
rect 179012 291864 179018 291876
rect 188338 291864 188344 291876
rect 188396 291864 188402 291916
rect 60458 291796 60464 291848
rect 60516 291836 60522 291848
rect 75178 291836 75184 291848
rect 60516 291808 75184 291836
rect 60516 291796 60522 291808
rect 75178 291796 75184 291808
rect 75236 291796 75242 291848
rect 151354 291796 151360 291848
rect 151412 291836 151418 291848
rect 189810 291836 189816 291848
rect 151412 291808 189816 291836
rect 151412 291796 151418 291808
rect 189810 291796 189816 291808
rect 189868 291796 189874 291848
rect 257338 291796 257344 291848
rect 257396 291836 257402 291848
rect 261018 291836 261024 291848
rect 257396 291808 261024 291836
rect 257396 291796 257402 291808
rect 261018 291796 261024 291808
rect 261076 291796 261082 291848
rect 98362 291252 98368 291304
rect 98420 291292 98426 291304
rect 99282 291292 99288 291304
rect 98420 291264 99288 291292
rect 98420 291252 98426 291264
rect 99282 291252 99288 291264
rect 99340 291252 99346 291304
rect 89530 291184 89536 291236
rect 89588 291224 89594 291236
rect 121546 291224 121552 291236
rect 89588 291196 121552 291224
rect 89588 291184 89594 291196
rect 121546 291184 121552 291196
rect 121604 291184 121610 291236
rect 255498 290980 255504 291032
rect 255556 291020 255562 291032
rect 258166 291020 258172 291032
rect 255556 290992 258172 291020
rect 255556 290980 255562 290992
rect 258166 290980 258172 290992
rect 258224 290980 258230 291032
rect 71866 290436 71872 290488
rect 71924 290476 71930 290488
rect 161934 290476 161940 290488
rect 71924 290448 161940 290476
rect 71924 290436 71930 290448
rect 161934 290436 161940 290448
rect 161992 290436 161998 290488
rect 188706 290028 188712 290080
rect 188764 290068 188770 290080
rect 188982 290068 188988 290080
rect 188764 290040 188988 290068
rect 188764 290028 188770 290040
rect 188982 290028 188988 290040
rect 189040 290068 189046 290080
rect 191190 290068 191196 290080
rect 189040 290040 191196 290068
rect 189040 290028 189046 290040
rect 191190 290028 191196 290040
rect 191248 290028 191254 290080
rect 162210 289824 162216 289876
rect 162268 289864 162274 289876
rect 191650 289864 191656 289876
rect 162268 289836 191656 289864
rect 162268 289824 162274 289836
rect 191650 289824 191656 289836
rect 191708 289824 191714 289876
rect 162762 289756 162768 289808
rect 162820 289796 162826 289808
rect 191742 289796 191748 289808
rect 162820 289768 191748 289796
rect 162820 289756 162826 289768
rect 191742 289756 191748 289768
rect 191800 289756 191806 289808
rect 260742 289756 260748 289808
rect 260800 289796 260806 289808
rect 269206 289796 269212 289808
rect 260800 289768 269212 289796
rect 260800 289756 260806 289768
rect 269206 289756 269212 289768
rect 269264 289756 269270 289808
rect 255498 289688 255504 289740
rect 255556 289728 255562 289740
rect 262490 289728 262496 289740
rect 255556 289700 262496 289728
rect 255556 289688 255562 289700
rect 262490 289688 262496 289700
rect 262548 289688 262554 289740
rect 76190 289416 76196 289468
rect 76248 289456 76254 289468
rect 76558 289456 76564 289468
rect 76248 289428 76564 289456
rect 76248 289416 76254 289428
rect 76558 289416 76564 289428
rect 76616 289416 76622 289468
rect 64782 289076 64788 289128
rect 64840 289116 64846 289128
rect 151078 289116 151084 289128
rect 64840 289088 151084 289116
rect 64840 289076 64846 289088
rect 151078 289076 151084 289088
rect 151136 289076 151142 289128
rect 159450 289076 159456 289128
rect 159508 289116 159514 289128
rect 162762 289116 162768 289128
rect 159508 289088 162768 289116
rect 159508 289076 159514 289088
rect 162762 289076 162768 289088
rect 162820 289076 162826 289128
rect 45462 288396 45468 288448
rect 45520 288436 45526 288448
rect 76190 288436 76196 288448
rect 45520 288408 76196 288436
rect 45520 288396 45526 288408
rect 76190 288396 76196 288408
rect 76248 288396 76254 288448
rect 79226 288396 79232 288448
rect 79284 288436 79290 288448
rect 79962 288436 79968 288448
rect 79284 288408 79968 288436
rect 79284 288396 79290 288408
rect 79962 288396 79968 288408
rect 80020 288436 80026 288448
rect 159450 288436 159456 288448
rect 80020 288408 159456 288436
rect 80020 288396 80026 288408
rect 159450 288396 159456 288408
rect 159508 288396 159514 288448
rect 35158 288328 35164 288380
rect 35216 288368 35222 288380
rect 70578 288368 70584 288380
rect 35216 288340 70584 288368
rect 35216 288328 35222 288340
rect 70578 288328 70584 288340
rect 70636 288368 70642 288380
rect 71038 288368 71044 288380
rect 70636 288340 71044 288368
rect 70636 288328 70642 288340
rect 71038 288328 71044 288340
rect 71096 288328 71102 288380
rect 255498 288328 255504 288380
rect 255556 288368 255562 288380
rect 281534 288368 281540 288380
rect 255556 288340 281540 288368
rect 255556 288328 255562 288340
rect 281534 288328 281540 288340
rect 281592 288328 281598 288380
rect 255314 288260 255320 288312
rect 255372 288300 255378 288312
rect 263778 288300 263784 288312
rect 255372 288272 263784 288300
rect 255372 288260 255378 288272
rect 263778 288260 263784 288272
rect 263836 288260 263842 288312
rect 74626 287784 74632 287836
rect 74684 287824 74690 287836
rect 75362 287824 75368 287836
rect 74684 287796 75368 287824
rect 74684 287784 74690 287796
rect 75362 287784 75368 287796
rect 75420 287784 75426 287836
rect 92474 287784 92480 287836
rect 92532 287824 92538 287836
rect 92934 287824 92940 287836
rect 92532 287796 92940 287824
rect 92532 287784 92538 287796
rect 92934 287784 92940 287796
rect 92992 287784 92998 287836
rect 68278 287716 68284 287768
rect 68336 287756 68342 287768
rect 158806 287756 158812 287768
rect 68336 287728 158812 287756
rect 68336 287716 68342 287728
rect 158806 287716 158812 287728
rect 158864 287716 158870 287768
rect 78582 287648 78588 287700
rect 78640 287688 78646 287700
rect 184198 287688 184204 287700
rect 78640 287660 184204 287688
rect 78640 287648 78646 287660
rect 184198 287648 184204 287660
rect 184256 287648 184262 287700
rect 182910 287512 182916 287564
rect 182968 287552 182974 287564
rect 190178 287552 190184 287564
rect 182968 287524 190184 287552
rect 182968 287512 182974 287524
rect 190178 287512 190184 287524
rect 190236 287512 190242 287564
rect 170490 286968 170496 287020
rect 170548 287008 170554 287020
rect 191742 287008 191748 287020
rect 170548 286980 191748 287008
rect 170548 286968 170554 286980
rect 191742 286968 191748 286980
rect 191800 286968 191806 287020
rect 255406 286628 255412 286680
rect 255464 286668 255470 286680
rect 257338 286668 257344 286680
rect 255464 286640 257344 286668
rect 255464 286628 255470 286640
rect 257338 286628 257344 286640
rect 257396 286628 257402 286680
rect 80422 286424 80428 286476
rect 80480 286464 80486 286476
rect 81250 286464 81256 286476
rect 80480 286436 81256 286464
rect 80480 286424 80486 286436
rect 81250 286424 81256 286436
rect 81308 286464 81314 286476
rect 83458 286464 83464 286476
rect 81308 286436 83464 286464
rect 81308 286424 81314 286436
rect 83458 286424 83464 286436
rect 83516 286424 83522 286476
rect 144178 286288 144184 286340
rect 144236 286328 144242 286340
rect 187050 286328 187056 286340
rect 144236 286300 187056 286328
rect 144236 286288 144242 286300
rect 187050 286288 187056 286300
rect 187108 286288 187114 286340
rect 255498 286288 255504 286340
rect 255556 286328 255562 286340
rect 258350 286328 258356 286340
rect 255556 286300 258356 286328
rect 255556 286288 255562 286300
rect 258350 286288 258356 286300
rect 258408 286328 258414 286340
rect 260834 286328 260840 286340
rect 258408 286300 260840 286328
rect 258408 286288 258414 286300
rect 260834 286288 260840 286300
rect 260892 286288 260898 286340
rect 81986 286084 81992 286136
rect 82044 286124 82050 286136
rect 82722 286124 82728 286136
rect 82044 286096 82728 286124
rect 82044 286084 82050 286096
rect 82722 286084 82728 286096
rect 82780 286124 82786 286136
rect 84654 286124 84660 286136
rect 82780 286096 84660 286124
rect 82780 286084 82786 286096
rect 84654 286084 84660 286096
rect 84712 286084 84718 286136
rect 95326 286084 95332 286136
rect 95384 286124 95390 286136
rect 97258 286124 97264 286136
rect 95384 286096 97264 286124
rect 95384 286084 95390 286096
rect 97258 286084 97264 286096
rect 97316 286084 97322 286136
rect 69014 285852 69020 285864
rect 60706 285824 69020 285852
rect 52178 285744 52184 285796
rect 52236 285784 52242 285796
rect 60706 285784 60734 285824
rect 69014 285812 69020 285824
rect 69072 285812 69078 285864
rect 73798 285852 73804 285864
rect 70366 285824 73804 285852
rect 70366 285784 70394 285824
rect 73798 285812 73804 285824
rect 73856 285812 73862 285864
rect 52236 285756 60734 285784
rect 65536 285756 70394 285784
rect 52236 285744 52242 285756
rect 53558 285676 53564 285728
rect 53616 285716 53622 285728
rect 65536 285716 65564 285756
rect 53616 285688 65564 285716
rect 53616 285676 53622 285688
rect 69014 285676 69020 285728
rect 69072 285716 69078 285728
rect 72418 285716 72424 285728
rect 69072 285688 72424 285716
rect 69072 285676 69078 285688
rect 72418 285676 72424 285688
rect 72476 285676 72482 285728
rect 87506 285676 87512 285728
rect 87564 285716 87570 285728
rect 90358 285716 90364 285728
rect 87564 285688 90364 285716
rect 87564 285676 87570 285688
rect 90358 285676 90364 285688
rect 90416 285676 90422 285728
rect 90818 285676 90824 285728
rect 90876 285716 90882 285728
rect 118050 285716 118056 285728
rect 90876 285688 118056 285716
rect 90876 285676 90882 285688
rect 118050 285676 118056 285688
rect 118108 285676 118114 285728
rect 167638 285676 167644 285728
rect 167696 285716 167702 285728
rect 170490 285716 170496 285728
rect 167696 285688 170496 285716
rect 167696 285676 167702 285688
rect 170490 285676 170496 285688
rect 170548 285676 170554 285728
rect 255406 285608 255412 285660
rect 255464 285648 255470 285660
rect 260926 285648 260932 285660
rect 255464 285620 260932 285648
rect 255464 285608 255470 285620
rect 260926 285608 260932 285620
rect 260984 285608 260990 285660
rect 54294 284928 54300 284980
rect 54352 284968 54358 284980
rect 87598 284968 87604 284980
rect 54352 284940 87604 284968
rect 54352 284928 54358 284940
rect 87598 284928 87604 284940
rect 87656 284928 87662 284980
rect 176562 284928 176568 284980
rect 176620 284968 176626 284980
rect 185578 284968 185584 284980
rect 176620 284940 185584 284968
rect 176620 284928 176626 284940
rect 185578 284928 185584 284940
rect 185636 284928 185642 284980
rect 91094 284384 91100 284436
rect 91152 284424 91158 284436
rect 98454 284424 98460 284436
rect 91152 284396 98460 284424
rect 91152 284384 91158 284396
rect 98454 284384 98460 284396
rect 98512 284384 98518 284436
rect 37918 284316 37924 284368
rect 37976 284356 37982 284368
rect 54294 284356 54300 284368
rect 37976 284328 54300 284356
rect 37976 284316 37982 284328
rect 54294 284316 54300 284328
rect 54352 284356 54358 284368
rect 54846 284356 54852 284368
rect 54352 284328 54852 284356
rect 54352 284316 54358 284328
rect 54846 284316 54852 284328
rect 54904 284316 54910 284368
rect 58894 284316 58900 284368
rect 58952 284356 58958 284368
rect 71866 284356 71872 284368
rect 58952 284328 71872 284356
rect 58952 284316 58958 284328
rect 71866 284316 71872 284328
rect 71924 284316 71930 284368
rect 88150 284316 88156 284368
rect 88208 284356 88214 284368
rect 99374 284356 99380 284368
rect 88208 284328 99380 284356
rect 88208 284316 88214 284328
rect 99374 284316 99380 284328
rect 99432 284316 99438 284368
rect 128262 284316 128268 284368
rect 128320 284356 128326 284368
rect 191742 284356 191748 284368
rect 128320 284328 191748 284356
rect 128320 284316 128326 284328
rect 191742 284316 191748 284328
rect 191800 284316 191806 284368
rect 266538 284316 266544 284368
rect 266596 284356 266602 284368
rect 266722 284356 266728 284368
rect 266596 284328 266728 284356
rect 266596 284316 266602 284328
rect 266722 284316 266728 284328
rect 266780 284316 266786 284368
rect 255406 284248 255412 284300
rect 255464 284288 255470 284300
rect 295610 284288 295616 284300
rect 255464 284260 295616 284288
rect 255464 284248 255470 284260
rect 295610 284248 295616 284260
rect 295668 284248 295674 284300
rect 169662 284112 169668 284164
rect 169720 284152 169726 284164
rect 169938 284152 169944 284164
rect 169720 284124 169944 284152
rect 169720 284112 169726 284124
rect 169938 284112 169944 284124
rect 169996 284112 170002 284164
rect 86080 283704 86086 283756
rect 86138 283744 86144 283756
rect 86862 283744 86868 283756
rect 86138 283716 86868 283744
rect 86138 283704 86144 283716
rect 86862 283704 86868 283716
rect 86920 283704 86926 283756
rect 52362 283568 52368 283620
rect 52420 283608 52426 283620
rect 56410 283608 56416 283620
rect 52420 283580 56416 283608
rect 52420 283568 52426 283580
rect 56410 283568 56416 283580
rect 56468 283608 56474 283620
rect 66254 283608 66260 283620
rect 56468 283580 66260 283608
rect 56468 283568 56474 283580
rect 66254 283568 66260 283580
rect 66312 283568 66318 283620
rect 162762 283568 162768 283620
rect 162820 283608 162826 283620
rect 176010 283608 176016 283620
rect 162820 283580 176016 283608
rect 162820 283568 162826 283580
rect 176010 283568 176016 283580
rect 176068 283568 176074 283620
rect 88610 283364 88616 283416
rect 88668 283404 88674 283416
rect 88978 283404 88984 283416
rect 88668 283376 88984 283404
rect 88668 283364 88674 283376
rect 88978 283364 88984 283376
rect 89036 283364 89042 283416
rect 98086 283364 98092 283416
rect 98144 283404 98150 283416
rect 98362 283404 98368 283416
rect 98144 283376 98368 283404
rect 98144 283364 98150 283376
rect 98362 283364 98368 283376
rect 98420 283364 98426 283416
rect 255498 283364 255504 283416
rect 255556 283404 255562 283416
rect 259730 283404 259736 283416
rect 255556 283376 259736 283404
rect 255556 283364 255562 283376
rect 259730 283364 259736 283376
rect 259788 283364 259794 283416
rect 68646 283228 68652 283280
rect 68704 283268 68710 283280
rect 69382 283268 69388 283280
rect 68704 283240 69388 283268
rect 68704 283228 68710 283240
rect 69382 283228 69388 283240
rect 69440 283268 69446 283280
rect 70302 283268 70308 283280
rect 69440 283240 70308 283268
rect 69440 283228 69446 283240
rect 70302 283228 70308 283240
rect 70360 283228 70366 283280
rect 83550 283228 83556 283280
rect 83608 283268 83614 283280
rect 84010 283268 84016 283280
rect 83608 283240 84016 283268
rect 83608 283228 83614 283240
rect 84010 283228 84016 283240
rect 84068 283228 84074 283280
rect 67542 283024 67548 283076
rect 67600 283064 67606 283076
rect 67600 283036 70394 283064
rect 67600 283024 67606 283036
rect 69658 282996 69664 283008
rect 69492 282968 69664 282996
rect 69014 282684 69020 282736
rect 69072 282724 69078 282736
rect 69492 282724 69520 282968
rect 69658 282956 69664 282968
rect 69716 282956 69722 283008
rect 70366 282996 70394 283036
rect 158714 282996 158720 283008
rect 70366 282968 158720 282996
rect 158714 282956 158720 282968
rect 158772 282956 158778 283008
rect 162762 282928 162768 282940
rect 69072 282696 69520 282724
rect 69768 282900 162768 282928
rect 69072 282684 69078 282696
rect 68922 282616 68928 282668
rect 68980 282656 68986 282668
rect 69768 282656 69796 282900
rect 162762 282888 162768 282900
rect 162820 282888 162826 282940
rect 175918 282888 175924 282940
rect 175976 282928 175982 282940
rect 180150 282928 180156 282940
rect 175976 282900 180156 282928
rect 175976 282888 175982 282900
rect 180150 282888 180156 282900
rect 180208 282928 180214 282940
rect 191742 282928 191748 282940
rect 180208 282900 191748 282928
rect 180208 282888 180214 282900
rect 191742 282888 191748 282900
rect 191800 282888 191806 282940
rect 98454 282820 98460 282872
rect 98512 282860 98518 282872
rect 163774 282860 163780 282872
rect 98512 282832 163780 282860
rect 98512 282820 98518 282832
rect 163774 282820 163780 282832
rect 163832 282820 163838 282872
rect 255498 282820 255504 282872
rect 255556 282860 255562 282872
rect 263594 282860 263600 282872
rect 255556 282832 263600 282860
rect 255556 282820 255562 282832
rect 263594 282820 263600 282832
rect 263652 282820 263658 282872
rect 68980 282628 69796 282656
rect 68980 282616 68986 282628
rect 68554 282140 68560 282192
rect 68612 282180 68618 282192
rect 98914 282180 98920 282192
rect 68612 282152 98920 282180
rect 68612 282140 68618 282152
rect 98914 282140 98920 282152
rect 98972 282140 98978 282192
rect 169018 282140 169024 282192
rect 169076 282180 169082 282192
rect 182818 282180 182824 282192
rect 169076 282152 182824 282180
rect 169076 282140 169082 282152
rect 182818 282140 182824 282152
rect 182876 282140 182882 282192
rect 259270 282140 259276 282192
rect 259328 282180 259334 282192
rect 267826 282180 267832 282192
rect 259328 282152 267832 282180
rect 259328 282140 259334 282152
rect 267826 282140 267832 282152
rect 267884 282140 267890 282192
rect 273438 282140 273444 282192
rect 273496 282180 273502 282192
rect 291378 282180 291384 282192
rect 273496 282152 291384 282180
rect 273496 282140 273502 282152
rect 291378 282140 291384 282152
rect 291436 282140 291442 282192
rect 255406 281936 255412 281988
rect 255464 281976 255470 281988
rect 259362 281976 259368 281988
rect 255464 281948 259368 281976
rect 255464 281936 255470 281948
rect 259362 281936 259368 281948
rect 259420 281936 259426 281988
rect 184290 281596 184296 281648
rect 184348 281636 184354 281648
rect 192018 281636 192024 281648
rect 184348 281608 192024 281636
rect 184348 281596 184354 281608
rect 192018 281596 192024 281608
rect 192076 281596 192082 281648
rect 100754 281528 100760 281580
rect 100812 281568 100818 281580
rect 108482 281568 108488 281580
rect 100812 281540 108488 281568
rect 100812 281528 100818 281540
rect 108482 281528 108488 281540
rect 108540 281528 108546 281580
rect 155494 281528 155500 281580
rect 155552 281568 155558 281580
rect 191742 281568 191748 281580
rect 155552 281540 191748 281568
rect 155552 281528 155558 281540
rect 191742 281528 191748 281540
rect 191800 281528 191806 281580
rect 100846 281460 100852 281512
rect 100904 281500 100910 281512
rect 103422 281500 103428 281512
rect 100904 281472 103428 281500
rect 100904 281460 100910 281472
rect 103422 281460 103428 281472
rect 103480 281500 103486 281512
rect 107562 281500 107568 281512
rect 103480 281472 107568 281500
rect 103480 281460 103486 281472
rect 107562 281460 107568 281472
rect 107620 281460 107626 281512
rect 255498 281460 255504 281512
rect 255556 281500 255562 281512
rect 276106 281500 276112 281512
rect 255556 281472 276112 281500
rect 255556 281460 255562 281472
rect 276106 281460 276112 281472
rect 276164 281460 276170 281512
rect 255406 281392 255412 281444
rect 255464 281432 255470 281444
rect 263686 281432 263692 281444
rect 255464 281404 263692 281432
rect 255464 281392 255470 281404
rect 263686 281392 263692 281404
rect 263744 281392 263750 281444
rect 160830 280780 160836 280832
rect 160888 280820 160894 280832
rect 161382 280820 161388 280832
rect 160888 280792 161388 280820
rect 160888 280780 160894 280792
rect 161382 280780 161388 280792
rect 161440 280820 161446 280832
rect 191742 280820 191748 280832
rect 161440 280792 191748 280820
rect 161440 280780 161446 280792
rect 191742 280780 191748 280792
rect 191800 280780 191806 280832
rect 175918 280644 175924 280696
rect 175976 280684 175982 280696
rect 178770 280684 178776 280696
rect 175976 280656 178776 280684
rect 175976 280644 175982 280656
rect 178770 280644 178776 280656
rect 178828 280644 178834 280696
rect 43438 280168 43444 280220
rect 43496 280208 43502 280220
rect 66714 280208 66720 280220
rect 43496 280180 66720 280208
rect 43496 280168 43502 280180
rect 66714 280168 66720 280180
rect 66772 280208 66778 280220
rect 68922 280208 68928 280220
rect 66772 280180 68928 280208
rect 66772 280168 66778 280180
rect 68922 280168 68928 280180
rect 68980 280168 68986 280220
rect 107010 280168 107016 280220
rect 107068 280208 107074 280220
rect 114462 280208 114468 280220
rect 107068 280180 114468 280208
rect 107068 280168 107074 280180
rect 114462 280168 114468 280180
rect 114520 280208 114526 280220
rect 114646 280208 114652 280220
rect 114520 280180 114652 280208
rect 114520 280168 114526 280180
rect 114646 280168 114652 280180
rect 114704 280168 114710 280220
rect 263594 280168 263600 280220
rect 263652 280208 263658 280220
rect 264238 280208 264244 280220
rect 263652 280180 264244 280208
rect 263652 280168 263658 280180
rect 264238 280168 264244 280180
rect 264296 280208 264302 280220
rect 292574 280208 292580 280220
rect 264296 280180 292580 280208
rect 264296 280168 264302 280180
rect 292574 280168 292580 280180
rect 292632 280168 292638 280220
rect 100754 280100 100760 280152
rect 100812 280140 100818 280152
rect 130470 280140 130476 280152
rect 100812 280112 103514 280140
rect 100812 280100 100818 280112
rect 103486 280004 103514 280112
rect 109006 280112 130476 280140
rect 109006 280004 109034 280112
rect 130470 280100 130476 280112
rect 130528 280100 130534 280152
rect 255498 280100 255504 280152
rect 255556 280140 255562 280152
rect 269390 280140 269396 280152
rect 255556 280112 269396 280140
rect 255556 280100 255562 280112
rect 269390 280100 269396 280112
rect 269448 280100 269454 280152
rect 103486 279976 109034 280004
rect 7558 279420 7564 279472
rect 7616 279460 7622 279472
rect 35802 279460 35808 279472
rect 7616 279432 35808 279460
rect 7616 279420 7622 279432
rect 35802 279420 35808 279432
rect 35860 279460 35866 279472
rect 60642 279460 60648 279472
rect 35860 279432 60648 279460
rect 35860 279420 35866 279432
rect 60642 279420 60648 279432
rect 60700 279460 60706 279472
rect 66806 279460 66812 279472
rect 60700 279432 66812 279460
rect 60700 279420 60706 279432
rect 66806 279420 66812 279432
rect 66864 279420 66870 279472
rect 123478 279420 123484 279472
rect 123536 279460 123542 279472
rect 153930 279460 153936 279472
rect 123536 279432 153936 279460
rect 123536 279420 123542 279432
rect 153930 279420 153936 279432
rect 153988 279420 153994 279472
rect 158714 278740 158720 278792
rect 158772 278780 158778 278792
rect 160186 278780 160192 278792
rect 158772 278752 160192 278780
rect 158772 278740 158778 278752
rect 160186 278740 160192 278752
rect 160244 278780 160250 278792
rect 191742 278780 191748 278792
rect 160244 278752 191748 278780
rect 160244 278740 160250 278752
rect 191742 278740 191748 278752
rect 191800 278740 191806 278792
rect 255406 278672 255412 278724
rect 255464 278712 255470 278724
rect 280338 278712 280344 278724
rect 255464 278684 280344 278712
rect 255464 278672 255470 278684
rect 280338 278672 280344 278684
rect 280396 278672 280402 278724
rect 255498 278604 255504 278656
rect 255556 278644 255562 278656
rect 263594 278644 263600 278656
rect 255556 278616 263600 278644
rect 255556 278604 255562 278616
rect 263594 278604 263600 278616
rect 263652 278604 263658 278656
rect 65886 278264 65892 278316
rect 65944 278304 65950 278316
rect 67542 278304 67548 278316
rect 65944 278276 67548 278304
rect 65944 278264 65950 278276
rect 67542 278264 67548 278276
rect 67600 278264 67606 278316
rect 99374 277992 99380 278044
rect 99432 278032 99438 278044
rect 118878 278032 118884 278044
rect 99432 278004 118884 278032
rect 99432 277992 99438 278004
rect 118878 277992 118884 278004
rect 118936 277992 118942 278044
rect 138658 277992 138664 278044
rect 138716 278032 138722 278044
rect 158438 278032 158444 278044
rect 138716 278004 158444 278032
rect 138716 277992 138722 278004
rect 158438 277992 158444 278004
rect 158496 278032 158502 278044
rect 183370 278032 183376 278044
rect 158496 278004 183376 278032
rect 158496 277992 158502 278004
rect 183370 277992 183376 278004
rect 183428 277992 183434 278044
rect 183370 277380 183376 277432
rect 183428 277420 183434 277432
rect 191558 277420 191564 277432
rect 183428 277392 191564 277420
rect 183428 277380 183434 277392
rect 191558 277380 191564 277392
rect 191616 277380 191622 277432
rect 52270 277312 52276 277364
rect 52328 277352 52334 277364
rect 66898 277352 66904 277364
rect 52328 277324 66904 277352
rect 52328 277312 52334 277324
rect 66898 277312 66904 277324
rect 66956 277312 66962 277364
rect 100202 277312 100208 277364
rect 100260 277352 100266 277364
rect 184658 277352 184664 277364
rect 100260 277324 184664 277352
rect 100260 277312 100266 277324
rect 184658 277312 184664 277324
rect 184716 277312 184722 277364
rect 255590 277312 255596 277364
rect 255648 277352 255654 277364
rect 278958 277352 278964 277364
rect 255648 277324 278964 277352
rect 255648 277312 255654 277324
rect 278958 277312 278964 277324
rect 279016 277312 279022 277364
rect 255406 276632 255412 276684
rect 255464 276672 255470 276684
rect 276290 276672 276296 276684
rect 255464 276644 276296 276672
rect 255464 276632 255470 276644
rect 276290 276632 276296 276644
rect 276348 276632 276354 276684
rect 184658 276088 184664 276140
rect 184716 276128 184722 276140
rect 189810 276128 189816 276140
rect 184716 276100 189816 276128
rect 184716 276088 184722 276100
rect 189810 276088 189816 276100
rect 189868 276088 189874 276140
rect 100754 276020 100760 276072
rect 100812 276060 100818 276072
rect 129090 276060 129096 276072
rect 100812 276032 129096 276060
rect 100812 276020 100818 276032
rect 129090 276020 129096 276032
rect 129148 276020 129154 276072
rect 151262 276020 151268 276072
rect 151320 276060 151326 276072
rect 191742 276060 191748 276072
rect 151320 276032 191748 276060
rect 151320 276020 151326 276032
rect 191742 276020 191748 276032
rect 191800 276020 191806 276072
rect 276106 276020 276112 276072
rect 276164 276060 276170 276072
rect 276290 276060 276296 276072
rect 276164 276032 276296 276060
rect 276164 276020 276170 276032
rect 276290 276020 276296 276032
rect 276348 276020 276354 276072
rect 61838 275952 61844 276004
rect 61896 275992 61902 276004
rect 66898 275992 66904 276004
rect 61896 275964 66904 275992
rect 61896 275952 61902 275964
rect 66898 275952 66904 275964
rect 66956 275952 66962 276004
rect 255498 275952 255504 276004
rect 255556 275992 255562 276004
rect 277670 275992 277676 276004
rect 255556 275964 277676 275992
rect 255556 275952 255562 275964
rect 277670 275952 277676 275964
rect 277728 275952 277734 276004
rect 100938 275272 100944 275324
rect 100996 275312 101002 275324
rect 155402 275312 155408 275324
rect 100996 275284 155408 275312
rect 100996 275272 101002 275284
rect 155402 275272 155408 275284
rect 155460 275272 155466 275324
rect 177942 275272 177948 275324
rect 178000 275312 178006 275324
rect 184198 275312 184204 275324
rect 178000 275284 184204 275312
rect 178000 275272 178006 275284
rect 184198 275272 184204 275284
rect 184256 275272 184262 275324
rect 100754 274660 100760 274712
rect 100812 274700 100818 274712
rect 136082 274700 136088 274712
rect 100812 274672 136088 274700
rect 100812 274660 100818 274672
rect 136082 274660 136088 274672
rect 136140 274660 136146 274712
rect 255406 274660 255412 274712
rect 255464 274700 255470 274712
rect 270678 274700 270684 274712
rect 255464 274672 270684 274700
rect 255464 274660 255470 274672
rect 270678 274660 270684 274672
rect 270736 274700 270742 274712
rect 272242 274700 272248 274712
rect 270736 274672 272248 274700
rect 270736 274660 270742 274672
rect 272242 274660 272248 274672
rect 272300 274660 272306 274712
rect 100846 274592 100852 274644
rect 100904 274632 100910 274644
rect 160738 274632 160744 274644
rect 100904 274604 160744 274632
rect 100904 274592 100910 274604
rect 160738 274592 160744 274604
rect 160796 274592 160802 274644
rect 163590 274592 163596 274644
rect 163648 274632 163654 274644
rect 182910 274632 182916 274644
rect 163648 274604 182916 274632
rect 163648 274592 163654 274604
rect 182910 274592 182916 274604
rect 182968 274592 182974 274644
rect 255498 274592 255504 274644
rect 255556 274632 255562 274644
rect 281718 274632 281724 274644
rect 255556 274604 281724 274632
rect 255556 274592 255562 274604
rect 281718 274592 281724 274604
rect 281776 274592 281782 274644
rect 255406 274252 255412 274304
rect 255464 274292 255470 274304
rect 259546 274292 259552 274304
rect 255464 274264 259552 274292
rect 255464 274252 255470 274264
rect 259546 274252 259552 274264
rect 259604 274252 259610 274304
rect 60642 273232 60648 273284
rect 60700 273272 60706 273284
rect 63310 273272 63316 273284
rect 60700 273244 63316 273272
rect 60700 273232 60706 273244
rect 63310 273232 63316 273244
rect 63368 273272 63374 273284
rect 66898 273272 66904 273284
rect 63368 273244 66904 273272
rect 63368 273232 63374 273244
rect 66898 273232 66904 273244
rect 66956 273232 66962 273284
rect 67266 273232 67272 273284
rect 67324 273272 67330 273284
rect 68278 273272 68284 273284
rect 67324 273244 68284 273272
rect 67324 273232 67330 273244
rect 68278 273232 68284 273244
rect 68336 273232 68342 273284
rect 156690 273232 156696 273284
rect 156748 273272 156754 273284
rect 160830 273272 160836 273284
rect 156748 273244 160836 273272
rect 156748 273232 156754 273244
rect 160830 273232 160836 273244
rect 160888 273232 160894 273284
rect 162762 273232 162768 273284
rect 162820 273272 162826 273284
rect 163590 273272 163596 273284
rect 162820 273244 163596 273272
rect 162820 273232 162826 273244
rect 163590 273232 163596 273244
rect 163648 273232 163654 273284
rect 185578 273232 185584 273284
rect 185636 273272 185642 273284
rect 188890 273272 188896 273284
rect 185636 273244 188896 273272
rect 185636 273232 185642 273244
rect 188890 273232 188896 273244
rect 188948 273272 188954 273284
rect 191742 273272 191748 273284
rect 188948 273244 191748 273272
rect 188948 273232 188954 273244
rect 191742 273232 191748 273244
rect 191800 273232 191806 273284
rect 100846 273164 100852 273216
rect 100904 273204 100910 273216
rect 107010 273204 107016 273216
rect 100904 273176 107016 273204
rect 100904 273164 100910 273176
rect 107010 273164 107016 273176
rect 107068 273164 107074 273216
rect 255406 273164 255412 273216
rect 255464 273204 255470 273216
rect 259454 273204 259460 273216
rect 255464 273176 259460 273204
rect 255464 273164 255470 273176
rect 259454 273164 259460 273176
rect 259512 273164 259518 273216
rect 291286 273164 291292 273216
rect 291344 273204 291350 273216
rect 580166 273204 580172 273216
rect 291344 273176 580172 273204
rect 291344 273164 291350 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 135990 272552 135996 272604
rect 136048 272592 136054 272604
rect 155218 272592 155224 272604
rect 136048 272564 155224 272592
rect 136048 272552 136054 272564
rect 155218 272552 155224 272564
rect 155276 272552 155282 272604
rect 100754 272484 100760 272536
rect 100812 272524 100818 272536
rect 113174 272524 113180 272536
rect 100812 272496 113180 272524
rect 100812 272484 100818 272496
rect 113174 272484 113180 272496
rect 113232 272524 113238 272536
rect 141694 272524 141700 272536
rect 113232 272496 141700 272524
rect 113232 272484 113238 272496
rect 141694 272484 141700 272496
rect 141752 272484 141758 272536
rect 281994 272484 282000 272536
rect 282052 272524 282058 272536
rect 290090 272524 290096 272536
rect 282052 272496 290096 272524
rect 282052 272484 282058 272496
rect 290090 272484 290096 272496
rect 290148 272484 290154 272536
rect 60550 271940 60556 271992
rect 60608 271980 60614 271992
rect 61746 271980 61752 271992
rect 60608 271952 61752 271980
rect 60608 271940 60614 271952
rect 61746 271940 61752 271952
rect 61804 271980 61810 271992
rect 66898 271980 66904 271992
rect 61804 271952 66904 271980
rect 61804 271940 61810 271952
rect 66898 271940 66904 271952
rect 66956 271940 66962 271992
rect 191282 271912 191288 271924
rect 161446 271884 191288 271912
rect 136542 271804 136548 271856
rect 136600 271844 136606 271856
rect 160094 271844 160100 271856
rect 136600 271816 160100 271844
rect 136600 271804 136606 271816
rect 160094 271804 160100 271816
rect 160152 271844 160158 271856
rect 161446 271844 161474 271884
rect 191282 271872 191288 271884
rect 191340 271872 191346 271924
rect 255406 271872 255412 271924
rect 255464 271912 255470 271924
rect 281718 271912 281724 271924
rect 255464 271884 281724 271912
rect 255464 271872 255470 271884
rect 281718 271872 281724 271884
rect 281776 271912 281782 271924
rect 281994 271912 282000 271924
rect 281776 271884 282000 271912
rect 281776 271872 281782 271884
rect 281994 271872 282000 271884
rect 282052 271872 282058 271924
rect 184290 271844 184296 271856
rect 160152 271816 161474 271844
rect 171106 271816 184296 271844
rect 160152 271804 160158 271816
rect 158622 271736 158628 271788
rect 158680 271776 158686 271788
rect 161474 271776 161480 271788
rect 158680 271748 161480 271776
rect 158680 271736 158686 271748
rect 161474 271736 161480 271748
rect 161532 271776 161538 271788
rect 171106 271776 171134 271816
rect 184290 271804 184296 271816
rect 184348 271804 184354 271856
rect 255498 271804 255504 271856
rect 255556 271844 255562 271856
rect 261570 271844 261576 271856
rect 255556 271816 261576 271844
rect 255556 271804 255562 271816
rect 261570 271804 261576 271816
rect 261628 271804 261634 271856
rect 161532 271748 171134 271776
rect 161532 271736 161538 271748
rect 100754 271192 100760 271244
rect 100812 271232 100818 271244
rect 114554 271232 114560 271244
rect 100812 271204 114560 271232
rect 100812 271192 100818 271204
rect 114554 271192 114560 271204
rect 114612 271192 114618 271244
rect 101214 271124 101220 271176
rect 101272 271164 101278 271176
rect 102042 271164 102048 271176
rect 101272 271136 102048 271164
rect 101272 271124 101278 271136
rect 102042 271124 102048 271136
rect 102100 271164 102106 271176
rect 133690 271164 133696 271176
rect 102100 271136 133696 271164
rect 102100 271124 102106 271136
rect 133690 271124 133696 271136
rect 133748 271124 133754 271176
rect 259362 271124 259368 271176
rect 259420 271164 259426 271176
rect 280430 271164 280436 271176
rect 259420 271136 280436 271164
rect 259420 271124 259426 271136
rect 280430 271124 280436 271136
rect 280488 271124 280494 271176
rect 184382 270648 184388 270700
rect 184440 270688 184446 270700
rect 186222 270688 186228 270700
rect 184440 270660 186228 270688
rect 184440 270648 184446 270660
rect 186222 270648 186228 270660
rect 186280 270688 186286 270700
rect 191742 270688 191748 270700
rect 186280 270660 191748 270688
rect 186280 270648 186286 270660
rect 191742 270648 191748 270660
rect 191800 270648 191806 270700
rect 64690 270580 64696 270632
rect 64748 270620 64754 270632
rect 66898 270620 66904 270632
rect 64748 270592 66904 270620
rect 64748 270580 64754 270592
rect 66898 270580 66904 270592
rect 66956 270580 66962 270632
rect 56502 270444 56508 270496
rect 56560 270484 56566 270496
rect 59078 270484 59084 270496
rect 56560 270456 59084 270484
rect 56560 270444 56566 270456
rect 59078 270444 59084 270456
rect 59136 270444 59142 270496
rect 133690 270444 133696 270496
rect 133748 270484 133754 270496
rect 151354 270484 151360 270496
rect 133748 270456 151360 270484
rect 133748 270444 133754 270456
rect 151354 270444 151360 270456
rect 151412 270444 151418 270496
rect 162118 270444 162124 270496
rect 162176 270484 162182 270496
rect 169570 270484 169576 270496
rect 162176 270456 169576 270484
rect 162176 270444 162182 270456
rect 169570 270444 169576 270456
rect 169628 270484 169634 270496
rect 191190 270484 191196 270496
rect 169628 270456 191196 270484
rect 169628 270444 169634 270456
rect 191190 270444 191196 270456
rect 191248 270444 191254 270496
rect 255406 270240 255412 270292
rect 255464 270280 255470 270292
rect 259362 270280 259368 270292
rect 255464 270252 259368 270280
rect 255464 270240 255470 270252
rect 259362 270240 259368 270252
rect 259420 270240 259426 270292
rect 41322 269764 41328 269816
rect 41380 269804 41386 269816
rect 50798 269804 50804 269816
rect 41380 269776 50804 269804
rect 41380 269764 41386 269776
rect 50798 269764 50804 269776
rect 50856 269764 50862 269816
rect 59078 269764 59084 269816
rect 59136 269804 59142 269816
rect 66898 269804 66904 269816
rect 59136 269776 66904 269804
rect 59136 269764 59142 269776
rect 66898 269764 66904 269776
rect 66956 269764 66962 269816
rect 98822 269764 98828 269816
rect 98880 269804 98886 269816
rect 159634 269804 159640 269816
rect 98880 269776 159640 269804
rect 98880 269764 98886 269776
rect 159634 269764 159640 269776
rect 159692 269764 159698 269816
rect 261018 269764 261024 269816
rect 261076 269804 261082 269816
rect 273254 269804 273260 269816
rect 261076 269776 273260 269804
rect 261076 269764 261082 269776
rect 273254 269764 273260 269776
rect 273312 269764 273318 269816
rect 255406 269152 255412 269204
rect 255464 269192 255470 269204
rect 261018 269192 261024 269204
rect 255464 269164 261024 269192
rect 255464 269152 255470 269164
rect 261018 269152 261024 269164
rect 261076 269152 261082 269204
rect 100754 269084 100760 269136
rect 100812 269124 100818 269136
rect 115474 269124 115480 269136
rect 100812 269096 115480 269124
rect 100812 269084 100818 269096
rect 115474 269084 115480 269096
rect 115532 269084 115538 269136
rect 178770 269084 178776 269136
rect 178828 269124 178834 269136
rect 193398 269124 193404 269136
rect 178828 269096 193404 269124
rect 178828 269084 178834 269096
rect 193398 269084 193404 269096
rect 193456 269084 193462 269136
rect 259362 269084 259368 269136
rect 259420 269124 259426 269136
rect 291286 269124 291292 269136
rect 259420 269096 291292 269124
rect 259420 269084 259426 269096
rect 291286 269084 291292 269096
rect 291344 269084 291350 269136
rect 52270 269016 52276 269068
rect 52328 269056 52334 269068
rect 53742 269056 53748 269068
rect 52328 269028 53748 269056
rect 52328 269016 52334 269028
rect 53742 269016 53748 269028
rect 53800 269056 53806 269068
rect 66714 269056 66720 269068
rect 53800 269028 66720 269056
rect 53800 269016 53806 269028
rect 66714 269016 66720 269028
rect 66772 269016 66778 269068
rect 166258 269016 166264 269068
rect 166316 269056 166322 269068
rect 167730 269056 167736 269068
rect 166316 269028 167736 269056
rect 166316 269016 166322 269028
rect 167730 269016 167736 269028
rect 167788 269016 167794 269068
rect 267826 269016 267832 269068
rect 267884 269056 267890 269068
rect 270770 269056 270776 269068
rect 267884 269028 270776 269056
rect 267884 269016 267890 269028
rect 270770 269016 270776 269028
rect 270828 269016 270834 269068
rect 100018 268336 100024 268388
rect 100076 268376 100082 268388
rect 115290 268376 115296 268388
rect 100076 268348 115296 268376
rect 100076 268336 100082 268348
rect 115290 268336 115296 268348
rect 115348 268336 115354 268388
rect 120810 268336 120816 268388
rect 120868 268376 120874 268388
rect 133138 268376 133144 268388
rect 120868 268348 133144 268376
rect 120868 268336 120874 268348
rect 133138 268336 133144 268348
rect 133196 268336 133202 268388
rect 181898 268336 181904 268388
rect 181956 268376 181962 268388
rect 192570 268376 192576 268388
rect 181956 268348 192576 268376
rect 181956 268336 181962 268348
rect 192570 268336 192576 268348
rect 192628 268336 192634 268388
rect 255406 268336 255412 268388
rect 255464 268376 255470 268388
rect 271138 268376 271144 268388
rect 255464 268348 271144 268376
rect 255464 268336 255470 268348
rect 271138 268336 271144 268348
rect 271196 268376 271202 268388
rect 271782 268376 271788 268388
rect 271196 268348 271788 268376
rect 271196 268336 271202 268348
rect 271782 268336 271788 268348
rect 271840 268336 271846 268388
rect 99006 267996 99012 268048
rect 99064 268036 99070 268048
rect 104250 268036 104256 268048
rect 99064 268008 104256 268036
rect 99064 267996 99070 268008
rect 104250 267996 104256 268008
rect 104308 267996 104314 268048
rect 255406 267724 255412 267776
rect 255464 267764 255470 267776
rect 267826 267764 267832 267776
rect 255464 267736 267832 267764
rect 255464 267724 255470 267736
rect 267826 267724 267832 267736
rect 267884 267724 267890 267776
rect 271782 267724 271788 267776
rect 271840 267764 271846 267776
rect 280430 267764 280436 267776
rect 271840 267736 280436 267764
rect 271840 267724 271846 267736
rect 280430 267724 280436 267736
rect 280488 267724 280494 267776
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 37918 267696 37924 267708
rect 3568 267668 37924 267696
rect 3568 267656 3574 267668
rect 37918 267656 37924 267668
rect 37976 267656 37982 267708
rect 50982 267656 50988 267708
rect 51040 267696 51046 267708
rect 60734 267696 60740 267708
rect 51040 267668 60740 267696
rect 51040 267656 51046 267668
rect 60734 267656 60740 267668
rect 60792 267656 60798 267708
rect 98730 267656 98736 267708
rect 98788 267696 98794 267708
rect 146202 267696 146208 267708
rect 98788 267668 146208 267696
rect 98788 267656 98794 267668
rect 146202 267656 146208 267668
rect 146260 267656 146266 267708
rect 100754 267044 100760 267096
rect 100812 267084 100818 267096
rect 106090 267084 106096 267096
rect 100812 267056 106096 267084
rect 100812 267044 100818 267056
rect 106090 267044 106096 267056
rect 106148 267044 106154 267096
rect 146202 267044 146208 267096
rect 146260 267084 146266 267096
rect 177390 267084 177396 267096
rect 146260 267056 177396 267084
rect 146260 267044 146266 267056
rect 177390 267044 177396 267056
rect 177448 267044 177454 267096
rect 118050 266976 118056 267028
rect 118108 267016 118114 267028
rect 182910 267016 182916 267028
rect 118108 266988 182916 267016
rect 118108 266976 118114 266988
rect 182910 266976 182916 266988
rect 182968 266976 182974 267028
rect 265618 266976 265624 267028
rect 265676 267016 265682 267028
rect 277486 267016 277492 267028
rect 265676 266988 277492 267016
rect 265676 266976 265682 266988
rect 277486 266976 277492 266988
rect 277544 266976 277550 267028
rect 62022 266364 62028 266416
rect 62080 266404 62086 266416
rect 64598 266404 64604 266416
rect 62080 266376 64604 266404
rect 62080 266364 62086 266376
rect 64598 266364 64604 266376
rect 64656 266404 64662 266416
rect 66898 266404 66904 266416
rect 64656 266376 66904 266404
rect 64656 266364 64662 266376
rect 66898 266364 66904 266376
rect 66956 266364 66962 266416
rect 106182 266364 106188 266416
rect 106240 266404 106246 266416
rect 112530 266404 112536 266416
rect 106240 266376 112536 266404
rect 106240 266364 106246 266376
rect 112530 266364 112536 266376
rect 112588 266364 112594 266416
rect 255406 266364 255412 266416
rect 255464 266404 255470 266416
rect 258350 266404 258356 266416
rect 255464 266376 258356 266404
rect 255464 266364 255470 266376
rect 258350 266364 258356 266376
rect 258408 266364 258414 266416
rect 270402 266364 270408 266416
rect 270460 266404 270466 266416
rect 270770 266404 270776 266416
rect 270460 266376 270776 266404
rect 270460 266364 270466 266376
rect 270770 266364 270776 266376
rect 270828 266364 270834 266416
rect 100754 265616 100760 265668
rect 100812 265656 100818 265668
rect 148594 265656 148600 265668
rect 100812 265628 148600 265656
rect 100812 265616 100818 265628
rect 148594 265616 148600 265628
rect 148652 265616 148658 265668
rect 163590 265616 163596 265668
rect 163648 265656 163654 265668
rect 191558 265656 191564 265668
rect 163648 265628 191564 265656
rect 163648 265616 163654 265628
rect 191558 265616 191564 265628
rect 191616 265616 191622 265668
rect 255314 265616 255320 265668
rect 255372 265656 255378 265668
rect 265066 265656 265072 265668
rect 255372 265628 265072 265656
rect 255372 265616 255378 265628
rect 265066 265616 265072 265628
rect 265124 265616 265130 265668
rect 63402 264936 63408 264988
rect 63460 264976 63466 264988
rect 66254 264976 66260 264988
rect 63460 264948 66260 264976
rect 63460 264936 63466 264948
rect 66254 264936 66260 264948
rect 66312 264936 66318 264988
rect 105630 264936 105636 264988
rect 105688 264976 105694 264988
rect 109678 264976 109684 264988
rect 105688 264948 109684 264976
rect 105688 264936 105694 264948
rect 109678 264936 109684 264948
rect 109736 264936 109742 264988
rect 170306 264936 170312 264988
rect 170364 264976 170370 264988
rect 191742 264976 191748 264988
rect 170364 264948 191748 264976
rect 170364 264936 170370 264948
rect 191742 264936 191748 264948
rect 191800 264936 191806 264988
rect 253842 264936 253848 264988
rect 253900 264976 253906 264988
rect 273254 264976 273260 264988
rect 253900 264948 273260 264976
rect 253900 264936 253906 264948
rect 273254 264936 273260 264948
rect 273312 264936 273318 264988
rect 3418 264868 3424 264920
rect 3476 264908 3482 264920
rect 32398 264908 32404 264920
rect 3476 264880 32404 264908
rect 3476 264868 3482 264880
rect 32398 264868 32404 264880
rect 32456 264868 32462 264920
rect 104434 264188 104440 264240
rect 104492 264228 104498 264240
rect 173342 264228 173348 264240
rect 104492 264200 173348 264228
rect 104492 264188 104498 264200
rect 173342 264188 173348 264200
rect 173400 264188 173406 264240
rect 255406 264188 255412 264240
rect 255464 264228 255470 264240
rect 255464 264200 258074 264228
rect 255464 264188 255470 264200
rect 184750 264120 184756 264172
rect 184808 264160 184814 264172
rect 191742 264160 191748 264172
rect 184808 264132 191748 264160
rect 184808 264120 184814 264132
rect 191742 264120 191748 264132
rect 191800 264120 191806 264172
rect 258046 264092 258074 264200
rect 263778 264092 263784 264104
rect 258046 264064 263784 264092
rect 263778 264052 263784 264064
rect 263836 264092 263842 264104
rect 264330 264092 264336 264104
rect 263836 264064 264336 264092
rect 263836 264052 263842 264064
rect 264330 264052 264336 264064
rect 264388 264052 264394 264104
rect 60550 263848 60556 263900
rect 60608 263888 60614 263900
rect 61654 263888 61660 263900
rect 60608 263860 61660 263888
rect 60608 263848 60614 263860
rect 61654 263848 61660 263860
rect 61712 263888 61718 263900
rect 66254 263888 66260 263900
rect 61712 263860 66260 263888
rect 61712 263848 61718 263860
rect 66254 263848 66260 263860
rect 66312 263848 66318 263900
rect 100754 263576 100760 263628
rect 100812 263616 100818 263628
rect 113818 263616 113824 263628
rect 100812 263588 113824 263616
rect 100812 263576 100818 263588
rect 113818 263576 113824 263588
rect 113876 263576 113882 263628
rect 255498 263576 255504 263628
rect 255556 263616 255562 263628
rect 259730 263616 259736 263628
rect 255556 263588 259736 263616
rect 255556 263576 255562 263588
rect 259730 263576 259736 263588
rect 259788 263576 259794 263628
rect 100662 263508 100668 263560
rect 100720 263548 100726 263560
rect 113082 263548 113088 263560
rect 100720 263520 113088 263548
rect 100720 263508 100726 263520
rect 113082 263508 113088 263520
rect 113140 263548 113146 263560
rect 155494 263548 155500 263560
rect 113140 263520 155500 263548
rect 113140 263508 113146 263520
rect 155494 263508 155500 263520
rect 155552 263508 155558 263560
rect 255406 263508 255412 263560
rect 255464 263548 255470 263560
rect 274726 263548 274732 263560
rect 255464 263520 274732 263548
rect 255464 263508 255470 263520
rect 274726 263508 274732 263520
rect 274784 263548 274790 263560
rect 277394 263548 277400 263560
rect 274784 263520 277400 263548
rect 274784 263508 274790 263520
rect 277394 263508 277400 263520
rect 277452 263508 277458 263560
rect 255498 262828 255504 262880
rect 255556 262868 255562 262880
rect 287238 262868 287244 262880
rect 255556 262840 287244 262868
rect 255556 262828 255562 262840
rect 287238 262828 287244 262840
rect 287296 262828 287302 262880
rect 7558 262216 7564 262268
rect 7616 262256 7622 262268
rect 49510 262256 49516 262268
rect 7616 262228 49516 262256
rect 7616 262216 7622 262228
rect 49510 262216 49516 262228
rect 49568 262256 49574 262268
rect 66254 262256 66260 262268
rect 49568 262228 66260 262256
rect 49568 262216 49574 262228
rect 66254 262216 66260 262228
rect 66312 262216 66318 262268
rect 191742 262256 191748 262268
rect 165540 262228 191748 262256
rect 99282 262148 99288 262200
rect 99340 262188 99346 262200
rect 104342 262188 104348 262200
rect 99340 262160 104348 262188
rect 99340 262148 99346 262160
rect 104342 262148 104348 262160
rect 104400 262148 104406 262200
rect 133782 262080 133788 262132
rect 133840 262120 133846 262132
rect 164234 262120 164240 262132
rect 133840 262092 164240 262120
rect 133840 262080 133846 262092
rect 164234 262080 164240 262092
rect 164292 262120 164298 262132
rect 165540 262120 165568 262228
rect 191742 262216 191748 262228
rect 191800 262216 191806 262268
rect 191558 262188 191564 262200
rect 164292 262092 165568 262120
rect 171106 262160 191564 262188
rect 164292 262080 164298 262092
rect 165522 262012 165528 262064
rect 165580 262052 165586 262064
rect 171106 262052 171134 262160
rect 191558 262148 191564 262160
rect 191616 262148 191622 262200
rect 165580 262024 171134 262052
rect 165580 262012 165586 262024
rect 104802 261944 104808 261996
rect 104860 261984 104866 261996
rect 110598 261984 110604 261996
rect 104860 261956 110604 261984
rect 104860 261944 104866 261956
rect 110598 261944 110604 261956
rect 110656 261944 110662 261996
rect 50890 261536 50896 261588
rect 50948 261576 50954 261588
rect 66254 261576 66260 261588
rect 50948 261548 66260 261576
rect 50948 261536 50954 261548
rect 66254 261536 66260 261548
rect 66312 261536 66318 261588
rect 4062 261468 4068 261520
rect 4120 261508 4126 261520
rect 66162 261508 66168 261520
rect 4120 261480 66168 261508
rect 4120 261468 4126 261480
rect 66162 261468 66168 261480
rect 66220 261468 66226 261520
rect 111794 261468 111800 261520
rect 111852 261508 111858 261520
rect 129182 261508 129188 261520
rect 111852 261480 129188 261508
rect 111852 261468 111858 261480
rect 129182 261468 129188 261480
rect 129240 261468 129246 261520
rect 149882 261468 149888 261520
rect 149940 261508 149946 261520
rect 166258 261508 166264 261520
rect 149940 261480 166264 261508
rect 149940 261468 149946 261480
rect 166258 261468 166264 261480
rect 166316 261468 166322 261520
rect 255498 261468 255504 261520
rect 255556 261508 255562 261520
rect 278314 261508 278320 261520
rect 255556 261480 278320 261508
rect 255556 261468 255562 261480
rect 278314 261468 278320 261480
rect 278372 261468 278378 261520
rect 266446 260788 266452 260840
rect 266504 260828 266510 260840
rect 279418 260828 279424 260840
rect 266504 260800 279424 260828
rect 266504 260788 266510 260800
rect 279418 260788 279424 260800
rect 279476 260788 279482 260840
rect 188982 260176 188988 260228
rect 189040 260216 189046 260228
rect 193214 260216 193220 260228
rect 189040 260188 193220 260216
rect 189040 260176 189046 260188
rect 193214 260176 193220 260188
rect 193272 260176 193278 260228
rect 43990 260108 43996 260160
rect 44048 260148 44054 260160
rect 66254 260148 66260 260160
rect 44048 260120 66260 260148
rect 44048 260108 44054 260120
rect 66254 260108 66260 260120
rect 66312 260108 66318 260160
rect 173250 260108 173256 260160
rect 173308 260148 173314 260160
rect 191742 260148 191748 260160
rect 173308 260120 191748 260148
rect 173308 260108 173314 260120
rect 191742 260108 191748 260120
rect 191800 260108 191806 260160
rect 255406 260108 255412 260160
rect 255464 260148 255470 260160
rect 266446 260148 266452 260160
rect 255464 260120 266452 260148
rect 255464 260108 255470 260120
rect 266446 260108 266452 260120
rect 266504 260108 266510 260160
rect 100754 259496 100760 259548
rect 100812 259536 100818 259548
rect 137554 259536 137560 259548
rect 100812 259508 137560 259536
rect 100812 259496 100818 259508
rect 137554 259496 137560 259508
rect 137612 259496 137618 259548
rect 100846 259428 100852 259480
rect 100904 259468 100910 259480
rect 163774 259468 163780 259480
rect 100904 259440 163780 259468
rect 100904 259428 100910 259440
rect 163774 259428 163780 259440
rect 163832 259428 163838 259480
rect 255406 259428 255412 259480
rect 255464 259468 255470 259480
rect 263594 259468 263600 259480
rect 255464 259440 263600 259468
rect 255464 259428 255470 259440
rect 263594 259428 263600 259440
rect 263652 259428 263658 259480
rect 61930 259360 61936 259412
rect 61988 259400 61994 259412
rect 66622 259400 66628 259412
rect 61988 259372 66628 259400
rect 61988 259360 61994 259372
rect 66622 259360 66628 259372
rect 66680 259360 66686 259412
rect 255590 259360 255596 259412
rect 255648 259400 255654 259412
rect 294138 259400 294144 259412
rect 255648 259372 294144 259400
rect 255648 259360 255654 259372
rect 294138 259360 294144 259372
rect 294196 259360 294202 259412
rect 55122 258680 55128 258732
rect 55180 258720 55186 258732
rect 58986 258720 58992 258732
rect 55180 258692 58992 258720
rect 55180 258680 55186 258692
rect 58986 258680 58992 258692
rect 59044 258720 59050 258732
rect 66346 258720 66352 258732
rect 59044 258692 66352 258720
rect 59044 258680 59050 258692
rect 66346 258680 66352 258692
rect 66404 258680 66410 258732
rect 100754 258680 100760 258732
rect 100812 258720 100818 258732
rect 155310 258720 155316 258732
rect 100812 258692 155316 258720
rect 100812 258680 100818 258692
rect 155310 258680 155316 258692
rect 155368 258680 155374 258732
rect 255498 258680 255504 258732
rect 255556 258720 255562 258732
rect 266446 258720 266452 258732
rect 255556 258692 266452 258720
rect 255556 258680 255562 258692
rect 266446 258680 266452 258692
rect 266504 258680 266510 258732
rect 285950 258068 285956 258120
rect 286008 258108 286014 258120
rect 287330 258108 287336 258120
rect 286008 258080 287336 258108
rect 286008 258068 286014 258080
rect 287330 258068 287336 258080
rect 287388 258068 287394 258120
rect 66346 258000 66352 258052
rect 66404 258040 66410 258052
rect 68186 258040 68192 258052
rect 66404 258012 68192 258040
rect 66404 258000 66410 258012
rect 68186 258000 68192 258012
rect 68244 258000 68250 258052
rect 101674 258000 101680 258052
rect 101732 258040 101738 258052
rect 111058 258040 111064 258052
rect 101732 258012 111064 258040
rect 101732 258000 101738 258012
rect 111058 258000 111064 258012
rect 111116 258000 111122 258052
rect 44082 257320 44088 257372
rect 44140 257360 44146 257372
rect 53834 257360 53840 257372
rect 44140 257332 53840 257360
rect 44140 257320 44146 257332
rect 53834 257320 53840 257332
rect 53892 257320 53898 257372
rect 102042 257320 102048 257372
rect 102100 257360 102106 257372
rect 126422 257360 126428 257372
rect 102100 257332 126428 257360
rect 102100 257320 102106 257332
rect 126422 257320 126428 257332
rect 126480 257320 126486 257372
rect 136082 257320 136088 257372
rect 136140 257360 136146 257372
rect 178862 257360 178868 257372
rect 136140 257332 178868 257360
rect 136140 257320 136146 257332
rect 178862 257320 178868 257332
rect 178920 257320 178926 257372
rect 255406 256776 255412 256828
rect 255464 256816 255470 256828
rect 262582 256816 262588 256828
rect 255464 256788 262588 256816
rect 255464 256776 255470 256788
rect 262582 256776 262588 256788
rect 262640 256816 262646 256828
rect 262766 256816 262772 256828
rect 262640 256788 262772 256816
rect 262640 256776 262646 256788
rect 262766 256776 262772 256788
rect 262824 256776 262830 256828
rect 53834 256708 53840 256760
rect 53892 256748 53898 256760
rect 54938 256748 54944 256760
rect 53892 256720 54944 256748
rect 53892 256708 53898 256720
rect 54938 256708 54944 256720
rect 54996 256748 55002 256760
rect 66254 256748 66260 256760
rect 54996 256720 66260 256748
rect 54996 256708 55002 256720
rect 66254 256708 66260 256720
rect 66312 256708 66318 256760
rect 174538 256640 174544 256692
rect 174596 256680 174602 256692
rect 183462 256680 183468 256692
rect 174596 256652 183468 256680
rect 174596 256640 174602 256652
rect 183462 256640 183468 256652
rect 183520 256680 183526 256692
rect 190638 256680 190644 256692
rect 183520 256652 190644 256680
rect 183520 256640 183526 256652
rect 190638 256640 190644 256652
rect 190696 256640 190702 256692
rect 49602 255960 49608 256012
rect 49660 256000 49666 256012
rect 64598 256000 64604 256012
rect 49660 255972 64604 256000
rect 49660 255960 49666 255972
rect 64598 255960 64604 255972
rect 64656 256000 64662 256012
rect 66898 256000 66904 256012
rect 64656 255972 66904 256000
rect 64656 255960 64662 255972
rect 66898 255960 66904 255972
rect 66956 255960 66962 256012
rect 100846 255960 100852 256012
rect 100904 256000 100910 256012
rect 137370 256000 137376 256012
rect 100904 255972 137376 256000
rect 100904 255960 100910 255972
rect 137370 255960 137376 255972
rect 137428 255960 137434 256012
rect 283098 255960 283104 256012
rect 283156 256000 283162 256012
rect 580718 256000 580724 256012
rect 283156 255972 580724 256000
rect 283156 255960 283162 255972
rect 580718 255960 580724 255972
rect 580776 255960 580782 256012
rect 255406 255348 255412 255400
rect 255464 255388 255470 255400
rect 278958 255388 278964 255400
rect 255464 255360 278964 255388
rect 255464 255348 255470 255360
rect 278958 255348 278964 255360
rect 279016 255348 279022 255400
rect 100754 255280 100760 255332
rect 100812 255320 100818 255332
rect 188522 255320 188528 255332
rect 100812 255292 188528 255320
rect 100812 255280 100818 255292
rect 188522 255280 188528 255292
rect 188580 255280 188586 255332
rect 254578 255280 254584 255332
rect 254636 255320 254642 255332
rect 255590 255320 255596 255332
rect 254636 255292 255596 255320
rect 254636 255280 254642 255292
rect 255590 255280 255596 255292
rect 255648 255320 255654 255332
rect 283098 255320 283104 255332
rect 255648 255292 283104 255320
rect 255648 255280 255654 255292
rect 283098 255280 283104 255292
rect 283156 255280 283162 255332
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 43438 255252 43444 255264
rect 3476 255224 43444 255252
rect 3476 255212 3482 255224
rect 43438 255212 43444 255224
rect 43496 255212 43502 255264
rect 57882 254668 57888 254720
rect 57940 254708 57946 254720
rect 66898 254708 66904 254720
rect 57940 254680 66904 254708
rect 57940 254668 57946 254680
rect 66898 254668 66904 254680
rect 66956 254668 66962 254720
rect 272334 254600 272340 254652
rect 272392 254640 272398 254652
rect 280246 254640 280252 254652
rect 272392 254612 280252 254640
rect 272392 254600 272398 254612
rect 280246 254600 280252 254612
rect 280304 254600 280310 254652
rect 46842 254532 46848 254584
rect 46900 254572 46906 254584
rect 66714 254572 66720 254584
rect 46900 254544 66720 254572
rect 46900 254532 46906 254544
rect 66714 254532 66720 254544
rect 66772 254532 66778 254584
rect 126882 254532 126888 254584
rect 126940 254572 126946 254584
rect 162210 254572 162216 254584
rect 126940 254544 162216 254572
rect 126940 254532 126946 254544
rect 162210 254532 162216 254544
rect 162268 254532 162274 254584
rect 255406 254532 255412 254584
rect 255464 254572 255470 254584
rect 285950 254572 285956 254584
rect 255464 254544 285956 254572
rect 255464 254532 255470 254544
rect 285950 254532 285956 254544
rect 286008 254532 286014 254584
rect 100754 253988 100760 254040
rect 100812 254028 100818 254040
rect 111058 254028 111064 254040
rect 100812 254000 111064 254028
rect 100812 253988 100818 254000
rect 111058 253988 111064 254000
rect 111116 253988 111122 254040
rect 167822 253988 167828 254040
rect 167880 254028 167886 254040
rect 170766 254028 170772 254040
rect 167880 254000 170772 254028
rect 167880 253988 167886 254000
rect 170766 253988 170772 254000
rect 170824 254028 170830 254040
rect 184290 254028 184296 254040
rect 170824 254000 184296 254028
rect 170824 253988 170830 254000
rect 184290 253988 184296 254000
rect 184348 253988 184354 254040
rect 56594 253920 56600 253972
rect 56652 253960 56658 253972
rect 57882 253960 57888 253972
rect 56652 253932 57888 253960
rect 56652 253920 56658 253932
rect 57882 253920 57888 253932
rect 57940 253920 57946 253972
rect 102962 253920 102968 253972
rect 103020 253960 103026 253972
rect 103330 253960 103336 253972
rect 103020 253932 103336 253960
rect 103020 253920 103026 253932
rect 103330 253920 103336 253932
rect 103388 253960 103394 253972
rect 125594 253960 125600 253972
rect 103388 253932 125600 253960
rect 103388 253920 103394 253932
rect 125594 253920 125600 253932
rect 125652 253960 125658 253972
rect 126882 253960 126888 253972
rect 125652 253932 126888 253960
rect 125652 253920 125658 253932
rect 126882 253920 126888 253932
rect 126940 253920 126946 253972
rect 190638 253960 190644 253972
rect 161446 253932 190644 253960
rect 161446 253904 161474 253932
rect 190638 253920 190644 253932
rect 190696 253920 190702 253972
rect 255498 253920 255504 253972
rect 255556 253960 255562 253972
rect 271874 253960 271880 253972
rect 255556 253932 271880 253960
rect 255556 253920 255562 253932
rect 271874 253920 271880 253932
rect 271932 253960 271938 253972
rect 272334 253960 272340 253972
rect 271932 253932 272340 253960
rect 271932 253920 271938 253932
rect 272334 253920 272340 253932
rect 272392 253920 272398 253972
rect 63218 253852 63224 253904
rect 63276 253892 63282 253904
rect 66622 253892 66628 253904
rect 63276 253864 66628 253892
rect 63276 253852 63282 253864
rect 66622 253852 66628 253864
rect 66680 253852 66686 253904
rect 131022 253852 131028 253904
rect 131080 253892 131086 253904
rect 161446 253892 161480 253904
rect 131080 253864 161480 253892
rect 131080 253852 131086 253864
rect 161474 253852 161480 253864
rect 161532 253852 161538 253904
rect 163682 253240 163688 253292
rect 163740 253280 163746 253292
rect 174630 253280 174636 253292
rect 163740 253252 174636 253280
rect 163740 253240 163746 253252
rect 174630 253240 174636 253252
rect 174688 253240 174694 253292
rect 32398 253172 32404 253224
rect 32456 253212 32462 253224
rect 66898 253212 66904 253224
rect 32456 253184 66904 253212
rect 32456 253172 32462 253184
rect 66898 253172 66904 253184
rect 66956 253212 66962 253224
rect 67266 253212 67272 253224
rect 66956 253184 67272 253212
rect 66956 253172 66962 253184
rect 67266 253172 67272 253184
rect 67324 253172 67330 253224
rect 102870 253172 102876 253224
rect 102928 253212 102934 253224
rect 173802 253212 173808 253224
rect 102928 253184 173808 253212
rect 102928 253172 102934 253184
rect 173802 253172 173808 253184
rect 173860 253212 173866 253224
rect 174722 253212 174728 253224
rect 173860 253184 174728 253212
rect 173860 253172 173866 253184
rect 174722 253172 174728 253184
rect 174780 253172 174786 253224
rect 179322 253172 179328 253224
rect 179380 253212 179386 253224
rect 192662 253212 192668 253224
rect 179380 253184 192668 253212
rect 179380 253172 179386 253184
rect 192662 253172 192668 253184
rect 192720 253172 192726 253224
rect 255406 253172 255412 253224
rect 255464 253212 255470 253224
rect 262490 253212 262496 253224
rect 255464 253184 262496 253212
rect 255464 253172 255470 253184
rect 262490 253172 262496 253184
rect 262548 253172 262554 253224
rect 281626 252764 281632 252816
rect 281684 252804 281690 252816
rect 285858 252804 285864 252816
rect 281684 252776 285864 252804
rect 281684 252764 281690 252776
rect 285858 252764 285864 252776
rect 285916 252764 285922 252816
rect 101582 252492 101588 252544
rect 101640 252532 101646 252544
rect 104802 252532 104808 252544
rect 101640 252504 104808 252532
rect 101640 252492 101646 252504
rect 104802 252492 104808 252504
rect 104860 252532 104866 252544
rect 128262 252532 128268 252544
rect 104860 252504 128268 252532
rect 104860 252492 104866 252504
rect 128262 252492 128268 252504
rect 128320 252532 128326 252544
rect 129734 252532 129740 252544
rect 128320 252504 129740 252532
rect 128320 252492 128326 252504
rect 129734 252492 129740 252504
rect 129792 252492 129798 252544
rect 255498 251880 255504 251932
rect 255556 251920 255562 251932
rect 266446 251920 266452 251932
rect 255556 251892 266452 251920
rect 255556 251880 255562 251892
rect 266446 251880 266452 251892
rect 266504 251880 266510 251932
rect 55030 251812 55036 251864
rect 55088 251852 55094 251864
rect 66070 251852 66076 251864
rect 55088 251824 66076 251852
rect 55088 251812 55094 251824
rect 66070 251812 66076 251824
rect 66128 251852 66134 251864
rect 66622 251852 66628 251864
rect 66128 251824 66628 251852
rect 66128 251812 66134 251824
rect 66622 251812 66628 251824
rect 66680 251812 66686 251864
rect 164142 251812 164148 251864
rect 164200 251852 164206 251864
rect 191742 251852 191748 251864
rect 164200 251824 191748 251852
rect 164200 251812 164206 251824
rect 191742 251812 191748 251824
rect 191800 251812 191806 251864
rect 255406 251812 255412 251864
rect 255464 251852 255470 251864
rect 281626 251852 281632 251864
rect 255464 251824 281632 251852
rect 255464 251812 255470 251824
rect 281626 251812 281632 251824
rect 281684 251812 281690 251864
rect 64874 251132 64880 251184
rect 64932 251172 64938 251184
rect 66254 251172 66260 251184
rect 64932 251144 66260 251172
rect 64932 251132 64938 251144
rect 66254 251132 66260 251144
rect 66312 251132 66318 251184
rect 106090 251132 106096 251184
rect 106148 251172 106154 251184
rect 106918 251172 106924 251184
rect 106148 251144 106924 251172
rect 106148 251132 106154 251144
rect 106918 251132 106924 251144
rect 106976 251132 106982 251184
rect 169570 251132 169576 251184
rect 169628 251172 169634 251184
rect 191558 251172 191564 251184
rect 169628 251144 191564 251172
rect 169628 251132 169634 251144
rect 191558 251132 191564 251144
rect 191616 251132 191622 251184
rect 48130 250452 48136 250504
rect 48188 250492 48194 250504
rect 66990 250492 66996 250504
rect 48188 250464 66996 250492
rect 48188 250452 48194 250464
rect 66990 250452 66996 250464
rect 67048 250452 67054 250504
rect 100754 250452 100760 250504
rect 100812 250492 100818 250504
rect 106090 250492 106096 250504
rect 100812 250464 106096 250492
rect 100812 250452 100818 250464
rect 106090 250452 106096 250464
rect 106148 250452 106154 250504
rect 122190 250452 122196 250504
rect 122248 250492 122254 250504
rect 167822 250492 167828 250504
rect 122248 250464 167828 250492
rect 122248 250452 122254 250464
rect 167822 250452 167828 250464
rect 167880 250452 167886 250504
rect 274910 250452 274916 250504
rect 274968 250492 274974 250504
rect 582650 250492 582656 250504
rect 274968 250464 582656 250492
rect 274968 250452 274974 250464
rect 582650 250452 582656 250464
rect 582708 250452 582714 250504
rect 255498 249772 255504 249824
rect 255556 249812 255562 249824
rect 274910 249812 274916 249824
rect 255556 249784 274916 249812
rect 255556 249772 255562 249784
rect 274910 249772 274916 249784
rect 274968 249772 274974 249824
rect 165522 249568 165528 249620
rect 165580 249608 165586 249620
rect 168374 249608 168380 249620
rect 165580 249580 168380 249608
rect 165580 249568 165586 249580
rect 168374 249568 168380 249580
rect 168432 249568 168438 249620
rect 151262 249132 151268 249144
rect 132466 249104 151268 249132
rect 53650 249024 53656 249076
rect 53708 249064 53714 249076
rect 64782 249064 64788 249076
rect 53708 249036 64788 249064
rect 53708 249024 53714 249036
rect 64782 249024 64788 249036
rect 64840 249064 64846 249076
rect 66898 249064 66904 249076
rect 64840 249036 66904 249064
rect 64840 249024 64846 249036
rect 66898 249024 66904 249036
rect 66956 249024 66962 249076
rect 100846 249024 100852 249076
rect 100904 249064 100910 249076
rect 106182 249064 106188 249076
rect 100904 249036 106188 249064
rect 100904 249024 100910 249036
rect 106182 249024 106188 249036
rect 106240 249064 106246 249076
rect 129182 249064 129188 249076
rect 106240 249036 129188 249064
rect 106240 249024 106246 249036
rect 129182 249024 129188 249036
rect 129240 249064 129246 249076
rect 132466 249064 132494 249104
rect 151262 249092 151268 249104
rect 151320 249092 151326 249144
rect 129240 249036 132494 249064
rect 129240 249024 129246 249036
rect 137462 249024 137468 249076
rect 137520 249064 137526 249076
rect 160278 249064 160284 249076
rect 137520 249036 160284 249064
rect 137520 249024 137526 249036
rect 160278 249024 160284 249036
rect 160336 249024 160342 249076
rect 182818 249024 182824 249076
rect 182876 249064 182882 249076
rect 191650 249064 191656 249076
rect 182876 249036 191656 249064
rect 182876 249024 182882 249036
rect 191650 249024 191656 249036
rect 191708 249024 191714 249076
rect 187510 248820 187516 248872
rect 187568 248860 187574 248872
rect 191282 248860 191288 248872
rect 187568 248832 191288 248860
rect 187568 248820 187574 248832
rect 191282 248820 191288 248832
rect 191340 248820 191346 248872
rect 255406 248480 255412 248532
rect 255464 248520 255470 248532
rect 278038 248520 278044 248532
rect 255464 248492 278044 248520
rect 255464 248480 255470 248492
rect 278038 248480 278044 248492
rect 278096 248480 278102 248532
rect 255498 248412 255504 248464
rect 255556 248452 255562 248464
rect 292666 248452 292672 248464
rect 255556 248424 292672 248452
rect 255556 248412 255562 248424
rect 292666 248412 292672 248424
rect 292724 248452 292730 248464
rect 582466 248452 582472 248464
rect 292724 248424 582472 248452
rect 292724 248412 292730 248424
rect 582466 248412 582472 248424
rect 582524 248412 582530 248464
rect 148594 247664 148600 247716
rect 148652 247704 148658 247716
rect 180334 247704 180340 247716
rect 148652 247676 180340 247704
rect 148652 247664 148658 247676
rect 180334 247664 180340 247676
rect 180392 247664 180398 247716
rect 255498 247664 255504 247716
rect 255556 247704 255562 247716
rect 259546 247704 259552 247716
rect 255556 247676 259552 247704
rect 255556 247664 255562 247676
rect 259546 247664 259552 247676
rect 259604 247704 259610 247716
rect 271966 247704 271972 247716
rect 259604 247676 271972 247704
rect 259604 247664 259610 247676
rect 271966 247664 271972 247676
rect 272024 247664 272030 247716
rect 53650 247052 53656 247104
rect 53708 247092 53714 247104
rect 66622 247092 66628 247104
rect 53708 247064 66628 247092
rect 53708 247052 53714 247064
rect 66622 247052 66628 247064
rect 66680 247052 66686 247104
rect 181530 247052 181536 247104
rect 181588 247092 181594 247104
rect 191742 247092 191748 247104
rect 181588 247064 191748 247092
rect 181588 247052 181594 247064
rect 191742 247052 191748 247064
rect 191800 247052 191806 247104
rect 254118 247052 254124 247104
rect 254176 247092 254182 247104
rect 259638 247092 259644 247104
rect 254176 247064 259644 247092
rect 254176 247052 254182 247064
rect 259638 247052 259644 247064
rect 259696 247052 259702 247104
rect 59170 246984 59176 247036
rect 59228 247024 59234 247036
rect 64874 247024 64880 247036
rect 59228 246996 64880 247024
rect 59228 246984 59234 246996
rect 64874 246984 64880 246996
rect 64932 246984 64938 247036
rect 101030 246304 101036 246356
rect 101088 246344 101094 246356
rect 101398 246344 101404 246356
rect 101088 246316 101404 246344
rect 101088 246304 101094 246316
rect 101398 246304 101404 246316
rect 101456 246344 101462 246356
rect 159542 246344 159548 246356
rect 101456 246316 159548 246344
rect 101456 246304 101462 246316
rect 159542 246304 159548 246316
rect 159600 246304 159606 246356
rect 183370 246304 183376 246356
rect 183428 246344 183434 246356
rect 192478 246344 192484 246356
rect 183428 246316 192484 246344
rect 183428 246304 183434 246316
rect 192478 246304 192484 246316
rect 192536 246304 192542 246356
rect 280062 246304 280068 246356
rect 280120 246344 280126 246356
rect 298370 246344 298376 246356
rect 280120 246316 298376 246344
rect 280120 246304 280126 246316
rect 298370 246304 298376 246316
rect 298428 246304 298434 246356
rect 254670 246168 254676 246220
rect 254728 246208 254734 246220
rect 258350 246208 258356 246220
rect 254728 246180 258356 246208
rect 254728 246168 254734 246180
rect 258350 246168 258356 246180
rect 258408 246168 258414 246220
rect 166350 245624 166356 245676
rect 166408 245664 166414 245676
rect 169846 245664 169852 245676
rect 166408 245636 169852 245664
rect 166408 245624 166414 245636
rect 169846 245624 169852 245636
rect 169904 245624 169910 245676
rect 255682 245624 255688 245676
rect 255740 245664 255746 245676
rect 279418 245664 279424 245676
rect 255740 245636 279424 245664
rect 255740 245624 255746 245636
rect 279418 245624 279424 245636
rect 279476 245664 279482 245676
rect 280062 245664 280068 245676
rect 279476 245636 280068 245664
rect 279476 245624 279482 245636
rect 280062 245624 280068 245636
rect 280120 245624 280126 245676
rect 100938 245556 100944 245608
rect 100996 245596 101002 245608
rect 165614 245596 165620 245608
rect 100996 245568 165620 245596
rect 100996 245556 101002 245568
rect 165614 245556 165620 245568
rect 165672 245556 165678 245608
rect 255498 245556 255504 245608
rect 255556 245596 255562 245608
rect 289814 245596 289820 245608
rect 255556 245568 289820 245596
rect 255556 245556 255562 245568
rect 289814 245556 289820 245568
rect 289872 245556 289878 245608
rect 100846 245148 100852 245200
rect 100904 245188 100910 245200
rect 105630 245188 105636 245200
rect 100904 245160 105636 245188
rect 100904 245148 100910 245160
rect 105630 245148 105636 245160
rect 105688 245148 105694 245200
rect 184198 244944 184204 244996
rect 184256 244984 184262 244996
rect 193674 244984 193680 244996
rect 184256 244956 193680 244984
rect 184256 244944 184262 244956
rect 193674 244944 193680 244956
rect 193732 244944 193738 244996
rect 165614 244876 165620 244928
rect 165672 244916 165678 244928
rect 193122 244916 193128 244928
rect 165672 244888 193128 244916
rect 165672 244876 165678 244888
rect 193122 244876 193128 244888
rect 193180 244876 193186 244928
rect 255590 244876 255596 244928
rect 255648 244916 255654 244928
rect 258534 244916 258540 244928
rect 255648 244888 258540 244916
rect 255648 244876 255654 244888
rect 258534 244876 258540 244888
rect 258592 244916 258598 244928
rect 284294 244916 284300 244928
rect 258592 244888 284300 244916
rect 258592 244876 258598 244888
rect 284294 244876 284300 244888
rect 284352 244876 284358 244928
rect 289814 244264 289820 244316
rect 289872 244304 289878 244316
rect 294046 244304 294052 244316
rect 289872 244276 294052 244304
rect 289872 244264 289878 244276
rect 294046 244264 294052 244276
rect 294104 244264 294110 244316
rect 57698 244196 57704 244248
rect 57756 244236 57762 244248
rect 66898 244236 66904 244248
rect 57756 244208 66904 244236
rect 57756 244196 57762 244208
rect 66898 244196 66904 244208
rect 66956 244196 66962 244248
rect 98546 243516 98552 243568
rect 98604 243556 98610 243568
rect 106274 243556 106280 243568
rect 98604 243528 106280 243556
rect 98604 243516 98610 243528
rect 106274 243516 106280 243528
rect 106332 243516 106338 243568
rect 106918 243516 106924 243568
rect 106976 243556 106982 243568
rect 125042 243556 125048 243568
rect 106976 243528 125048 243556
rect 106976 243516 106982 243528
rect 125042 243516 125048 243528
rect 125100 243516 125106 243568
rect 153838 243516 153844 243568
rect 153896 243556 153902 243568
rect 189074 243556 189080 243568
rect 153896 243528 189080 243556
rect 153896 243516 153902 243528
rect 189074 243516 189080 243528
rect 189132 243516 189138 243568
rect 255498 243516 255504 243568
rect 255556 243556 255562 243568
rect 277486 243556 277492 243568
rect 255556 243528 277492 243556
rect 255556 243516 255562 243528
rect 277486 243516 277492 243528
rect 277544 243556 277550 243568
rect 280246 243556 280252 243568
rect 277544 243528 280252 243556
rect 277544 243516 277550 243528
rect 280246 243516 280252 243528
rect 280304 243516 280310 243568
rect 100846 243448 100852 243500
rect 100904 243488 100910 243500
rect 102778 243488 102784 243500
rect 100904 243460 102784 243488
rect 100904 243448 100910 243460
rect 102778 243448 102784 243460
rect 102836 243448 102842 243500
rect 185670 243448 185676 243500
rect 185728 243488 185734 243500
rect 258166 243488 258172 243500
rect 185728 243460 198136 243488
rect 185728 243448 185734 243460
rect 173802 243176 173808 243228
rect 173860 243216 173866 243228
rect 176654 243216 176660 243228
rect 173860 243188 176660 243216
rect 173860 243176 173866 243188
rect 176654 243176 176660 243188
rect 176712 243176 176718 243228
rect 57698 242904 57704 242956
rect 57756 242944 57762 242956
rect 66530 242944 66536 242956
rect 57756 242916 66536 242944
rect 57756 242904 57762 242916
rect 66530 242904 66536 242916
rect 66588 242904 66594 242956
rect 189074 242904 189080 242956
rect 189132 242944 189138 242956
rect 191742 242944 191748 242956
rect 189132 242916 191748 242944
rect 189132 242904 189138 242916
rect 191742 242904 191748 242916
rect 191800 242904 191806 242956
rect 141694 242836 141700 242888
rect 141752 242876 141758 242888
rect 141752 242848 180794 242876
rect 141752 242836 141758 242848
rect 180766 242808 180794 242848
rect 184842 242836 184848 242888
rect 184900 242876 184906 242888
rect 191098 242876 191104 242888
rect 184900 242848 191104 242876
rect 184900 242836 184906 242848
rect 191098 242836 191104 242848
rect 191156 242836 191162 242888
rect 186314 242808 186320 242820
rect 180766 242780 186320 242808
rect 186314 242768 186320 242780
rect 186372 242768 186378 242820
rect 100846 242224 100852 242276
rect 100904 242264 100910 242276
rect 103606 242264 103612 242276
rect 100904 242236 103612 242264
rect 100904 242224 100910 242236
rect 103606 242224 103612 242236
rect 103664 242224 103670 242276
rect 186314 242224 186320 242276
rect 186372 242264 186378 242276
rect 187602 242264 187608 242276
rect 186372 242236 187608 242264
rect 186372 242224 186378 242236
rect 187602 242224 187608 242236
rect 187660 242264 187666 242276
rect 193582 242264 193588 242276
rect 187660 242236 193588 242264
rect 187660 242224 187666 242236
rect 193582 242224 193588 242236
rect 193640 242224 193646 242276
rect 69014 242156 69020 242208
rect 69072 242196 69078 242208
rect 98178 242196 98184 242208
rect 69072 242168 98184 242196
rect 69072 242156 69078 242168
rect 98178 242156 98184 242168
rect 98236 242156 98242 242208
rect 198108 242072 198136 243460
rect 248386 243460 258172 243488
rect 248386 242944 248414 243460
rect 258166 243448 258172 243460
rect 258224 243448 258230 243500
rect 243004 242916 248414 242944
rect 243004 242072 243032 242916
rect 255682 242836 255688 242888
rect 255740 242876 255746 242888
rect 258350 242876 258356 242888
rect 255740 242848 258356 242876
rect 255740 242836 255746 242848
rect 258350 242836 258356 242848
rect 258408 242876 258414 242888
rect 259270 242876 259276 242888
rect 258408 242848 259276 242876
rect 258408 242836 258414 242848
rect 259270 242836 259276 242848
rect 259328 242836 259334 242888
rect 252370 242292 252376 242344
rect 252428 242332 252434 242344
rect 252922 242332 252928 242344
rect 252428 242304 252928 242332
rect 252428 242292 252434 242304
rect 252922 242292 252928 242304
rect 252980 242292 252986 242344
rect 259270 242224 259276 242276
rect 259328 242264 259334 242276
rect 278774 242264 278780 242276
rect 259328 242236 278780 242264
rect 259328 242224 259334 242236
rect 278774 242224 278780 242236
rect 278832 242224 278838 242276
rect 255498 242156 255504 242208
rect 255556 242196 255562 242208
rect 284386 242196 284392 242208
rect 255556 242168 284392 242196
rect 255556 242156 255562 242168
rect 284386 242156 284392 242168
rect 284444 242156 284450 242208
rect 192662 242020 192668 242072
rect 192720 242060 192726 242072
rect 197998 242060 198004 242072
rect 192720 242032 198004 242060
rect 192720 242020 192726 242032
rect 197998 242020 198004 242032
rect 198056 242020 198062 242072
rect 198090 242020 198096 242072
rect 198148 242020 198154 242072
rect 242986 242020 242992 242072
rect 243044 242020 243050 242072
rect 95418 241748 95424 241800
rect 95476 241788 95482 241800
rect 102962 241788 102968 241800
rect 95476 241760 102968 241788
rect 95476 241748 95482 241760
rect 102962 241748 102968 241760
rect 103020 241748 103026 241800
rect 57882 241476 57888 241528
rect 57940 241516 57946 241528
rect 66898 241516 66904 241528
rect 57940 241488 66904 241516
rect 57940 241476 57946 241488
rect 66898 241476 66904 241488
rect 66956 241476 66962 241528
rect 193674 241476 193680 241528
rect 193732 241516 193738 241528
rect 215294 241516 215300 241528
rect 193732 241488 215300 241516
rect 193732 241476 193738 241488
rect 215294 241476 215300 241488
rect 215352 241516 215358 241528
rect 216306 241516 216312 241528
rect 215352 241488 216312 241516
rect 215352 241476 215358 241488
rect 216306 241476 216312 241488
rect 216364 241476 216370 241528
rect 22830 241408 22836 241460
rect 22888 241448 22894 241460
rect 93440 241448 93446 241460
rect 22888 241420 93446 241448
rect 22888 241408 22894 241420
rect 93440 241408 93446 241420
rect 93498 241408 93504 241460
rect 255590 241408 255596 241460
rect 255648 241448 255654 241460
rect 268102 241448 268108 241460
rect 255648 241420 268108 241448
rect 255648 241408 255654 241420
rect 268102 241408 268108 241420
rect 268160 241448 268166 241460
rect 283006 241448 283012 241460
rect 268160 241420 283012 241448
rect 268160 241408 268166 241420
rect 283006 241408 283012 241420
rect 283064 241408 283070 241460
rect 3418 241068 3424 241120
rect 3476 241108 3482 241120
rect 7558 241108 7564 241120
rect 3476 241080 7564 241108
rect 3476 241068 3482 241080
rect 7558 241068 7564 241080
rect 7616 241068 7622 241120
rect 94038 240796 94044 240848
rect 94096 240836 94102 240848
rect 126974 240836 126980 240848
rect 94096 240808 126980 240836
rect 94096 240796 94102 240808
rect 126974 240796 126980 240808
rect 127032 240796 127038 240848
rect 110598 240728 110604 240780
rect 110656 240768 110662 240780
rect 180702 240768 180708 240780
rect 110656 240740 180708 240768
rect 110656 240728 110662 240740
rect 180702 240728 180708 240740
rect 180760 240728 180766 240780
rect 193122 240728 193128 240780
rect 193180 240768 193186 240780
rect 207290 240768 207296 240780
rect 193180 240740 207296 240768
rect 193180 240728 193186 240740
rect 207290 240728 207296 240740
rect 207348 240728 207354 240780
rect 250438 240728 250444 240780
rect 250496 240768 250502 240780
rect 266630 240768 266636 240780
rect 250496 240740 266636 240768
rect 250496 240728 250502 240740
rect 266630 240728 266636 240740
rect 266688 240728 266694 240780
rect 68646 240592 68652 240644
rect 68704 240632 68710 240644
rect 76650 240632 76656 240644
rect 68704 240604 76656 240632
rect 68704 240592 68710 240604
rect 76650 240592 76656 240604
rect 76708 240592 76714 240644
rect 249058 240592 249064 240644
rect 249116 240632 249122 240644
rect 254118 240632 254124 240644
rect 249116 240604 254124 240632
rect 249116 240592 249122 240604
rect 254118 240592 254124 240604
rect 254176 240592 254182 240644
rect 69014 240116 69020 240168
rect 69072 240156 69078 240168
rect 69934 240156 69940 240168
rect 69072 240128 69940 240156
rect 69072 240116 69078 240128
rect 69934 240116 69940 240128
rect 69992 240116 69998 240168
rect 73154 240116 73160 240168
rect 73212 240156 73218 240168
rect 73798 240156 73804 240168
rect 73212 240128 73804 240156
rect 73212 240116 73218 240128
rect 73798 240116 73804 240128
rect 73856 240116 73862 240168
rect 74534 240116 74540 240168
rect 74592 240156 74598 240168
rect 75454 240156 75460 240168
rect 74592 240128 75460 240156
rect 74592 240116 74598 240128
rect 75454 240116 75460 240128
rect 75512 240116 75518 240168
rect 78674 240116 78680 240168
rect 78732 240156 78738 240168
rect 79318 240156 79324 240168
rect 78732 240128 79324 240156
rect 78732 240116 78738 240128
rect 79318 240116 79324 240128
rect 79376 240116 79382 240168
rect 89714 240116 89720 240168
rect 89772 240156 89778 240168
rect 90358 240156 90364 240168
rect 89772 240128 90364 240156
rect 89772 240116 89778 240128
rect 90358 240116 90364 240128
rect 90416 240116 90422 240168
rect 126974 240116 126980 240168
rect 127032 240156 127038 240168
rect 225598 240156 225604 240168
rect 127032 240128 225604 240156
rect 127032 240116 127038 240128
rect 225598 240116 225604 240128
rect 225656 240116 225662 240168
rect 48222 240048 48228 240100
rect 48280 240088 48286 240100
rect 76006 240088 76012 240100
rect 48280 240060 76012 240088
rect 48280 240048 48286 240060
rect 76006 240048 76012 240060
rect 76064 240048 76070 240100
rect 76558 240048 76564 240100
rect 76616 240088 76622 240100
rect 78214 240088 78220 240100
rect 76616 240060 78220 240088
rect 76616 240048 76622 240060
rect 78214 240048 78220 240060
rect 78272 240048 78278 240100
rect 80974 240048 80980 240100
rect 81032 240088 81038 240100
rect 81802 240088 81808 240100
rect 81032 240060 81808 240088
rect 81032 240048 81038 240060
rect 81802 240048 81808 240060
rect 81860 240048 81866 240100
rect 182082 240048 182088 240100
rect 182140 240088 182146 240100
rect 211522 240088 211528 240100
rect 182140 240060 211528 240088
rect 182140 240048 182146 240060
rect 211522 240048 211528 240060
rect 211580 240088 211586 240100
rect 213178 240088 213184 240100
rect 211580 240060 213184 240088
rect 211580 240048 211586 240060
rect 213178 240048 213184 240060
rect 213236 240048 213242 240100
rect 70486 239980 70492 240032
rect 70544 240020 70550 240032
rect 71314 240020 71320 240032
rect 70544 239992 71320 240020
rect 70544 239980 70550 239992
rect 71314 239980 71320 239992
rect 71372 239980 71378 240032
rect 98546 239980 98552 240032
rect 98604 240020 98610 240032
rect 166902 240020 166908 240032
rect 98604 239992 166908 240020
rect 98604 239980 98610 239992
rect 166902 239980 166908 239992
rect 166960 240020 166966 240032
rect 195330 240020 195336 240032
rect 166960 239992 195336 240020
rect 166960 239980 166966 239992
rect 195330 239980 195336 239992
rect 195388 239980 195394 240032
rect 89622 239912 89628 239964
rect 89680 239952 89686 239964
rect 182082 239952 182088 239964
rect 89680 239924 182088 239952
rect 89680 239912 89686 239924
rect 182082 239912 182088 239924
rect 182140 239912 182146 239964
rect 71774 239776 71780 239828
rect 71832 239816 71838 239828
rect 72694 239816 72700 239828
rect 71832 239788 72700 239816
rect 71832 239776 71838 239788
rect 72694 239776 72700 239788
rect 72752 239776 72758 239828
rect 75178 239640 75184 239692
rect 75236 239680 75242 239692
rect 77294 239680 77300 239692
rect 75236 239652 77300 239680
rect 75236 239640 75242 239652
rect 77294 239640 77300 239652
rect 77352 239640 77358 239692
rect 82630 239504 82636 239556
rect 82688 239544 82694 239556
rect 88426 239544 88432 239556
rect 82688 239516 88432 239544
rect 82688 239504 82694 239516
rect 88426 239504 88432 239516
rect 88484 239504 88490 239556
rect 83642 239436 83648 239488
rect 83700 239476 83706 239488
rect 91002 239476 91008 239488
rect 83700 239448 91008 239476
rect 83700 239436 83706 239448
rect 91002 239436 91008 239448
rect 91060 239436 91066 239488
rect 224218 239368 224224 239420
rect 224276 239408 224282 239420
rect 235534 239408 235540 239420
rect 224276 239380 235540 239408
rect 224276 239368 224282 239380
rect 235534 239368 235540 239380
rect 235592 239368 235598 239420
rect 252462 239368 252468 239420
rect 252520 239408 252526 239420
rect 261478 239408 261484 239420
rect 252520 239380 261484 239408
rect 252520 239368 252526 239380
rect 261478 239368 261484 239380
rect 261536 239368 261542 239420
rect 91278 239300 91284 239352
rect 91336 239340 91342 239352
rect 93946 239340 93952 239352
rect 91336 239312 93952 239340
rect 91336 239300 91342 239312
rect 93946 239300 93952 239312
rect 94004 239300 94010 239352
rect 252094 239164 252100 239216
rect 252152 239204 252158 239216
rect 254026 239204 254032 239216
rect 252152 239176 254032 239204
rect 252152 239164 252158 239176
rect 254026 239164 254032 239176
rect 254084 239164 254090 239216
rect 224862 238960 224868 239012
rect 224920 239000 224926 239012
rect 225966 239000 225972 239012
rect 224920 238972 225972 239000
rect 224920 238960 224926 238972
rect 225966 238960 225972 238972
rect 226024 238960 226030 239012
rect 84930 238756 84936 238808
rect 84988 238796 84994 238808
rect 85482 238796 85488 238808
rect 84988 238768 85488 238796
rect 84988 238756 84994 238768
rect 85482 238756 85488 238768
rect 85540 238756 85546 238808
rect 46750 238688 46756 238740
rect 46808 238728 46814 238740
rect 74994 238728 75000 238740
rect 46808 238700 75000 238728
rect 46808 238688 46814 238700
rect 74994 238688 75000 238700
rect 75052 238688 75058 238740
rect 160002 238688 160008 238740
rect 160060 238728 160066 238740
rect 261018 238728 261024 238740
rect 160060 238700 261024 238728
rect 160060 238688 160066 238700
rect 261018 238688 261024 238700
rect 261076 238688 261082 238740
rect 80790 238620 80796 238672
rect 80848 238660 80854 238672
rect 164878 238660 164884 238672
rect 80848 238632 164884 238660
rect 80848 238620 80854 238632
rect 164878 238620 164884 238632
rect 164936 238620 164942 238672
rect 222102 238620 222108 238672
rect 222160 238660 222166 238672
rect 270770 238660 270776 238672
rect 222160 238632 270776 238660
rect 222160 238620 222166 238632
rect 270770 238620 270776 238632
rect 270828 238620 270834 238672
rect 193766 238484 193772 238536
rect 193824 238524 193830 238536
rect 193824 238496 200114 238524
rect 193824 238484 193830 238496
rect 200086 238388 200114 238496
rect 201494 238388 201500 238400
rect 200086 238360 201500 238388
rect 201494 238348 201500 238360
rect 201552 238388 201558 238400
rect 201954 238388 201960 238400
rect 201552 238360 201960 238388
rect 201552 238348 201558 238360
rect 201954 238348 201960 238360
rect 202012 238348 202018 238400
rect 93854 238008 93860 238060
rect 93912 238048 93918 238060
rect 113174 238048 113180 238060
rect 93912 238020 113180 238048
rect 93912 238008 93918 238020
rect 113174 238008 113180 238020
rect 113232 238048 113238 238060
rect 122834 238048 122840 238060
rect 113232 238020 122840 238048
rect 113232 238008 113238 238020
rect 122834 238008 122840 238020
rect 122892 238008 122898 238060
rect 68554 237940 68560 237992
rect 68612 237980 68618 237992
rect 76742 237980 76748 237992
rect 68612 237952 76748 237980
rect 68612 237940 68618 237952
rect 76742 237940 76748 237952
rect 76800 237940 76806 237992
rect 221090 237668 221096 237720
rect 221148 237708 221154 237720
rect 222102 237708 222108 237720
rect 221148 237680 222108 237708
rect 221148 237668 221154 237680
rect 222102 237668 222108 237680
rect 222160 237668 222166 237720
rect 78582 237396 78588 237448
rect 78640 237436 78646 237448
rect 78766 237436 78772 237448
rect 78640 237408 78772 237436
rect 78640 237396 78646 237408
rect 78766 237396 78772 237408
rect 78824 237396 78830 237448
rect 67818 237328 67824 237380
rect 67876 237368 67882 237380
rect 166350 237368 166356 237380
rect 67876 237340 166356 237368
rect 67876 237328 67882 237340
rect 166350 237328 166356 237340
rect 166408 237328 166414 237380
rect 193674 237328 193680 237380
rect 193732 237368 193738 237380
rect 213914 237368 213920 237380
rect 193732 237340 213920 237368
rect 193732 237328 193738 237340
rect 213914 237328 213920 237340
rect 213972 237328 213978 237380
rect 164878 237260 164884 237312
rect 164936 237300 164942 237312
rect 196618 237300 196624 237312
rect 164936 237272 196624 237300
rect 164936 237260 164942 237272
rect 196618 237260 196624 237272
rect 196676 237260 196682 237312
rect 86954 237124 86960 237176
rect 87012 237164 87018 237176
rect 87598 237164 87604 237176
rect 87012 237136 87604 237164
rect 87012 237124 87018 237136
rect 87598 237124 87604 237136
rect 87656 237124 87662 237176
rect 196618 236716 196624 236768
rect 196676 236756 196682 236768
rect 197170 236756 197176 236768
rect 196676 236728 197176 236756
rect 196676 236716 196682 236728
rect 197170 236716 197176 236728
rect 197228 236716 197234 236768
rect 214650 236716 214656 236768
rect 214708 236756 214714 236768
rect 252370 236756 252376 236768
rect 214708 236728 252376 236756
rect 214708 236716 214714 236728
rect 252370 236716 252376 236728
rect 252428 236716 252434 236768
rect 50982 236648 50988 236700
rect 51040 236688 51046 236700
rect 71866 236688 71872 236700
rect 51040 236660 71872 236688
rect 51040 236648 51046 236660
rect 71866 236648 71872 236660
rect 71924 236648 71930 236700
rect 93946 236648 93952 236700
rect 94004 236688 94010 236700
rect 116670 236688 116676 236700
rect 94004 236660 116676 236688
rect 94004 236648 94010 236660
rect 116670 236648 116676 236660
rect 116728 236688 116734 236700
rect 118694 236688 118700 236700
rect 116728 236660 118700 236688
rect 116728 236648 116734 236660
rect 118694 236648 118700 236660
rect 118752 236648 118758 236700
rect 197354 236648 197360 236700
rect 197412 236688 197418 236700
rect 259730 236688 259736 236700
rect 197412 236660 259736 236688
rect 197412 236648 197418 236660
rect 259730 236648 259736 236660
rect 259788 236648 259794 236700
rect 118970 236240 118976 236292
rect 119028 236280 119034 236292
rect 124950 236280 124956 236292
rect 119028 236252 124956 236280
rect 119028 236240 119034 236252
rect 124950 236240 124956 236252
rect 125008 236240 125014 236292
rect 89530 235968 89536 236020
rect 89588 236008 89594 236020
rect 89806 236008 89812 236020
rect 89588 235980 89812 236008
rect 89588 235968 89594 235980
rect 89806 235968 89812 235980
rect 89864 235968 89870 236020
rect 213914 235968 213920 236020
rect 213972 236008 213978 236020
rect 214558 236008 214564 236020
rect 213972 235980 214564 236008
rect 213972 235968 213978 235980
rect 214558 235968 214564 235980
rect 214616 235968 214622 236020
rect 89346 235900 89352 235952
rect 89404 235940 89410 235952
rect 110506 235940 110512 235952
rect 89404 235912 110512 235940
rect 89404 235900 89410 235912
rect 110506 235900 110512 235912
rect 110564 235900 110570 235952
rect 115474 235900 115480 235952
rect 115532 235940 115538 235952
rect 259546 235940 259552 235952
rect 115532 235912 259552 235940
rect 115532 235900 115538 235912
rect 259546 235900 259552 235912
rect 259604 235940 259610 235952
rect 259822 235940 259828 235952
rect 259604 235912 259828 235940
rect 259604 235900 259610 235912
rect 259822 235900 259828 235912
rect 259880 235900 259886 235952
rect 182910 235832 182916 235884
rect 182968 235872 182974 235884
rect 265250 235872 265256 235884
rect 182968 235844 265256 235872
rect 182968 235832 182974 235844
rect 265250 235832 265256 235844
rect 265308 235832 265314 235884
rect 280154 235220 280160 235272
rect 280212 235260 280218 235272
rect 580258 235260 580264 235272
rect 280212 235232 580264 235260
rect 280212 235220 280218 235232
rect 580258 235220 580264 235232
rect 580316 235220 580322 235272
rect 182910 235016 182916 235068
rect 182968 235056 182974 235068
rect 183462 235056 183468 235068
rect 182968 235028 183468 235056
rect 182968 235016 182974 235028
rect 183462 235016 183468 235028
rect 183520 235016 183526 235068
rect 43438 234608 43444 234660
rect 43496 234648 43502 234660
rect 96890 234648 96896 234660
rect 43496 234620 96896 234648
rect 43496 234608 43502 234620
rect 96890 234608 96896 234620
rect 96948 234648 96954 234660
rect 97350 234648 97356 234660
rect 96948 234620 97356 234648
rect 96948 234608 96954 234620
rect 97350 234608 97356 234620
rect 97408 234608 97414 234660
rect 97902 234608 97908 234660
rect 97960 234648 97966 234660
rect 99466 234648 99472 234660
rect 97960 234620 99472 234648
rect 97960 234608 97966 234620
rect 99466 234608 99472 234620
rect 99524 234608 99530 234660
rect 88334 234540 88340 234592
rect 88392 234580 88398 234592
rect 120718 234580 120724 234592
rect 88392 234552 120724 234580
rect 88392 234540 88398 234552
rect 120718 234540 120724 234552
rect 120776 234580 120782 234592
rect 122926 234580 122932 234592
rect 120776 234552 122932 234580
rect 120776 234540 120782 234552
rect 122926 234540 122932 234552
rect 122984 234540 122990 234592
rect 167730 234540 167736 234592
rect 167788 234580 167794 234592
rect 256786 234580 256792 234592
rect 167788 234552 256792 234580
rect 167788 234540 167794 234552
rect 256786 234540 256792 234552
rect 256844 234540 256850 234592
rect 137830 234472 137836 234524
rect 137888 234512 137894 234524
rect 181530 234512 181536 234524
rect 137888 234484 181536 234512
rect 137888 234472 137894 234484
rect 181530 234472 181536 234484
rect 181588 234472 181594 234524
rect 192570 234472 192576 234524
rect 192628 234512 192634 234524
rect 205634 234512 205640 234524
rect 192628 234484 205640 234512
rect 192628 234472 192634 234484
rect 205634 234472 205640 234484
rect 205692 234472 205698 234524
rect 207658 234472 207664 234524
rect 207716 234512 207722 234524
rect 266538 234512 266544 234524
rect 207716 234484 266544 234512
rect 207716 234472 207722 234484
rect 266538 234472 266544 234484
rect 266596 234472 266602 234524
rect 205634 234064 205640 234116
rect 205692 234104 205698 234116
rect 206738 234104 206744 234116
rect 205692 234076 206744 234104
rect 205692 234064 205698 234076
rect 206738 234064 206744 234076
rect 206796 234064 206802 234116
rect 97258 233860 97264 233912
rect 97316 233900 97322 233912
rect 98086 233900 98092 233912
rect 97316 233872 98092 233900
rect 97316 233860 97322 233872
rect 98086 233860 98092 233872
rect 98144 233860 98150 233912
rect 69106 233180 69112 233232
rect 69164 233220 69170 233232
rect 171042 233220 171048 233232
rect 69164 233192 171048 233220
rect 69164 233180 69170 233192
rect 171042 233180 171048 233192
rect 171100 233180 171106 233232
rect 207290 233180 207296 233232
rect 207348 233220 207354 233232
rect 237374 233220 237380 233232
rect 207348 233192 237380 233220
rect 207348 233180 207354 233192
rect 237374 233180 237380 233192
rect 237432 233220 237438 233232
rect 237926 233220 237932 233232
rect 237432 233192 237932 233220
rect 237432 233180 237438 233192
rect 237926 233180 237932 233192
rect 237984 233180 237990 233232
rect 54846 233112 54852 233164
rect 54904 233152 54910 233164
rect 87046 233152 87052 233164
rect 54904 233124 87052 233152
rect 54904 233112 54910 233124
rect 87046 233112 87052 233124
rect 87104 233152 87110 233164
rect 88242 233152 88248 233164
rect 87104 233124 88248 233152
rect 87104 233112 87110 233124
rect 88242 233112 88248 233124
rect 88300 233112 88306 233164
rect 89714 233112 89720 233164
rect 89772 233152 89778 233164
rect 116578 233152 116584 233164
rect 89772 233124 116584 233152
rect 89772 233112 89778 233124
rect 116578 233112 116584 233124
rect 116636 233152 116642 233164
rect 122190 233152 122196 233164
rect 116636 233124 122196 233152
rect 116636 233112 116642 233124
rect 122190 233112 122196 233124
rect 122248 233112 122254 233164
rect 247678 232568 247684 232620
rect 247736 232608 247742 232620
rect 262306 232608 262312 232620
rect 247736 232580 262312 232608
rect 247736 232568 247742 232580
rect 262306 232568 262312 232580
rect 262364 232568 262370 232620
rect 242158 232500 242164 232552
rect 242216 232540 242222 232552
rect 268010 232540 268016 232552
rect 242216 232512 268016 232540
rect 242216 232500 242222 232512
rect 268010 232500 268016 232512
rect 268068 232500 268074 232552
rect 278038 232500 278044 232552
rect 278096 232540 278102 232552
rect 580166 232540 580172 232552
rect 278096 232512 580172 232540
rect 278096 232500 278102 232512
rect 580166 232500 580172 232512
rect 580224 232500 580230 232552
rect 85482 231752 85488 231804
rect 85540 231792 85546 231804
rect 140866 231792 140872 231804
rect 85540 231764 140872 231792
rect 85540 231752 85546 231764
rect 140866 231752 140872 231764
rect 140924 231792 140930 231804
rect 141510 231792 141516 231804
rect 140924 231764 141516 231792
rect 140924 231752 140930 231764
rect 141510 231752 141516 231764
rect 141568 231752 141574 231804
rect 171042 231752 171048 231804
rect 171100 231792 171106 231804
rect 209130 231792 209136 231804
rect 171100 231764 209136 231792
rect 171100 231752 171106 231764
rect 209130 231752 209136 231764
rect 209188 231752 209194 231804
rect 225598 231752 225604 231804
rect 225656 231792 225662 231804
rect 292574 231792 292580 231804
rect 225656 231764 292580 231792
rect 225656 231752 225662 231764
rect 292574 231752 292580 231764
rect 292632 231752 292638 231804
rect 80054 231072 80060 231124
rect 80112 231112 80118 231124
rect 114646 231112 114652 231124
rect 80112 231084 114652 231112
rect 80112 231072 80118 231084
rect 114646 231072 114652 231084
rect 114704 231112 114710 231124
rect 123478 231112 123484 231124
rect 114704 231084 123484 231112
rect 114704 231072 114710 231084
rect 123478 231072 123484 231084
rect 123536 231072 123542 231124
rect 140866 231072 140872 231124
rect 140924 231112 140930 231124
rect 178862 231112 178868 231124
rect 140924 231084 178868 231112
rect 140924 231072 140930 231084
rect 178862 231072 178868 231084
rect 178920 231072 178926 231124
rect 246298 231072 246304 231124
rect 246356 231112 246362 231124
rect 267918 231112 267924 231124
rect 246356 231084 267924 231112
rect 246356 231072 246362 231084
rect 267918 231072 267924 231084
rect 267976 231072 267982 231124
rect 78674 230392 78680 230444
rect 78732 230432 78738 230444
rect 108942 230432 108948 230444
rect 78732 230404 108948 230432
rect 78732 230392 78738 230404
rect 108942 230392 108948 230404
rect 109000 230432 109006 230444
rect 111886 230432 111892 230444
rect 109000 230404 111892 230432
rect 109000 230392 109006 230404
rect 111886 230392 111892 230404
rect 111944 230392 111950 230444
rect 163774 230392 163780 230444
rect 163832 230432 163838 230444
rect 262398 230432 262404 230444
rect 163832 230404 262404 230432
rect 163832 230392 163838 230404
rect 262398 230392 262404 230404
rect 262456 230392 262462 230444
rect 268378 229984 268384 230036
rect 268436 230024 268442 230036
rect 272058 230024 272064 230036
rect 268436 229996 272064 230024
rect 268436 229984 268442 229996
rect 272058 229984 272064 229996
rect 272116 229984 272122 230036
rect 74534 229712 74540 229764
rect 74592 229752 74598 229764
rect 87598 229752 87604 229764
rect 74592 229724 87604 229752
rect 74592 229712 74598 229724
rect 87598 229712 87604 229724
rect 87656 229712 87662 229764
rect 88242 229712 88248 229764
rect 88300 229752 88306 229764
rect 103514 229752 103520 229764
rect 88300 229724 103520 229752
rect 88300 229712 88306 229724
rect 103514 229712 103520 229724
rect 103572 229712 103578 229764
rect 111058 229712 111064 229764
rect 111116 229752 111122 229764
rect 119338 229752 119344 229764
rect 111116 229724 119344 229752
rect 111116 229712 111122 229724
rect 119338 229712 119344 229724
rect 119396 229712 119402 229764
rect 152642 229712 152648 229764
rect 152700 229752 152706 229764
rect 219434 229752 219440 229764
rect 152700 229724 219440 229752
rect 152700 229712 152706 229724
rect 219434 229712 219440 229724
rect 219492 229752 219498 229764
rect 258350 229752 258356 229764
rect 219492 229724 258356 229752
rect 219492 229712 219498 229724
rect 258350 229712 258356 229724
rect 258408 229712 258414 229764
rect 278682 229576 278688 229628
rect 278740 229616 278746 229628
rect 284478 229616 284484 229628
rect 278740 229588 284484 229616
rect 278740 229576 278746 229588
rect 284478 229576 284484 229588
rect 284536 229576 284542 229628
rect 178862 229032 178868 229084
rect 178920 229072 178926 229084
rect 214650 229072 214656 229084
rect 178920 229044 214656 229072
rect 178920 229032 178926 229044
rect 214650 229032 214656 229044
rect 214708 229032 214714 229084
rect 223482 229032 223488 229084
rect 223540 229072 223546 229084
rect 289906 229072 289912 229084
rect 223540 229044 289912 229072
rect 223540 229032 223546 229044
rect 289906 229032 289912 229044
rect 289964 229032 289970 229084
rect 238018 228352 238024 228404
rect 238076 228392 238082 228404
rect 263778 228392 263784 228404
rect 238076 228364 263784 228392
rect 238076 228352 238082 228364
rect 263778 228352 263784 228364
rect 263836 228352 263842 228404
rect 49510 227740 49516 227792
rect 49568 227780 49574 227792
rect 55122 227780 55128 227792
rect 49568 227752 55128 227780
rect 49568 227740 49574 227752
rect 55122 227740 55128 227752
rect 55180 227780 55186 227792
rect 169938 227780 169944 227792
rect 55180 227752 169944 227780
rect 55180 227740 55186 227752
rect 169938 227740 169944 227752
rect 169996 227780 170002 227792
rect 170490 227780 170496 227792
rect 169996 227752 170496 227780
rect 169996 227740 170002 227752
rect 170490 227740 170496 227752
rect 170548 227740 170554 227792
rect 178862 227740 178868 227792
rect 178920 227780 178926 227792
rect 179322 227780 179328 227792
rect 178920 227752 179328 227780
rect 178920 227740 178926 227752
rect 179322 227740 179328 227752
rect 179380 227740 179386 227792
rect 222930 227740 222936 227792
rect 222988 227780 222994 227792
rect 223482 227780 223488 227792
rect 222988 227752 223488 227780
rect 222988 227740 222994 227752
rect 223482 227740 223488 227752
rect 223540 227740 223546 227792
rect 189718 227060 189724 227112
rect 189776 227100 189782 227112
rect 209038 227100 209044 227112
rect 189776 227072 209044 227100
rect 189776 227060 189782 227072
rect 209038 227060 209044 227072
rect 209096 227060 209102 227112
rect 108482 226992 108488 227044
rect 108540 227032 108546 227044
rect 229094 227032 229100 227044
rect 108540 227004 229100 227032
rect 108540 226992 108546 227004
rect 229094 226992 229100 227004
rect 229152 227032 229158 227044
rect 229922 227032 229928 227044
rect 229152 227004 229928 227032
rect 229152 226992 229158 227004
rect 229922 226992 229928 227004
rect 229980 226992 229986 227044
rect 256050 226788 256056 226840
rect 256108 226828 256114 226840
rect 259638 226828 259644 226840
rect 256108 226800 259644 226828
rect 256108 226788 256114 226800
rect 259638 226788 259644 226800
rect 259696 226788 259702 226840
rect 229922 226312 229928 226364
rect 229980 226352 229986 226364
rect 256050 226352 256056 226364
rect 229980 226324 256056 226352
rect 229980 226312 229986 226324
rect 256050 226312 256056 226324
rect 256108 226312 256114 226364
rect 137554 226244 137560 226296
rect 137612 226284 137618 226296
rect 280430 226284 280436 226296
rect 137612 226256 280436 226284
rect 137612 226244 137618 226256
rect 280430 226244 280436 226256
rect 280488 226244 280494 226296
rect 210510 226176 210516 226228
rect 210568 226216 210574 226228
rect 262490 226216 262496 226228
rect 210568 226188 262496 226216
rect 210568 226176 210574 226188
rect 262490 226176 262496 226188
rect 262548 226176 262554 226228
rect 280154 225020 280160 225072
rect 280212 225060 280218 225072
rect 280430 225060 280436 225072
rect 280212 225032 280436 225060
rect 280212 225020 280218 225032
rect 280430 225020 280436 225032
rect 280488 225020 280494 225072
rect 67358 224952 67364 225004
rect 67416 224992 67422 225004
rect 204162 224992 204168 225004
rect 67416 224964 204168 224992
rect 67416 224952 67422 224964
rect 204162 224952 204168 224964
rect 204220 224952 204226 225004
rect 210510 224952 210516 225004
rect 210568 224992 210574 225004
rect 210970 224992 210976 225004
rect 210568 224964 210976 224992
rect 210568 224952 210574 224964
rect 210970 224952 210976 224964
rect 211028 224952 211034 225004
rect 166350 224884 166356 224936
rect 166408 224924 166414 224936
rect 166902 224924 166908 224936
rect 166408 224896 166908 224924
rect 166408 224884 166414 224896
rect 166902 224884 166908 224896
rect 166960 224924 166966 224936
rect 204346 224924 204352 224936
rect 166960 224896 204352 224924
rect 166960 224884 166966 224896
rect 204346 224884 204352 224896
rect 204404 224884 204410 224936
rect 50798 224204 50804 224256
rect 50856 224244 50862 224256
rect 160738 224244 160744 224256
rect 50856 224216 160744 224244
rect 50856 224204 50862 224216
rect 160738 224204 160744 224216
rect 160796 224204 160802 224256
rect 191282 224204 191288 224256
rect 191340 224244 191346 224256
rect 194594 224244 194600 224256
rect 191340 224216 194600 224244
rect 191340 224204 191346 224216
rect 194594 224204 194600 224216
rect 194652 224204 194658 224256
rect 206278 224204 206284 224256
rect 206336 224244 206342 224256
rect 252554 224244 252560 224256
rect 206336 224216 252560 224244
rect 206336 224204 206342 224216
rect 252554 224204 252560 224216
rect 252612 224204 252618 224256
rect 253198 224204 253204 224256
rect 253256 224244 253262 224256
rect 270586 224244 270592 224256
rect 253256 224216 270592 224244
rect 253256 224204 253262 224216
rect 270586 224204 270592 224216
rect 270644 224204 270650 224256
rect 165522 223524 165528 223576
rect 165580 223564 165586 223576
rect 274910 223564 274916 223576
rect 165580 223536 274916 223564
rect 165580 223524 165586 223536
rect 274910 223524 274916 223536
rect 274968 223524 274974 223576
rect 56502 222844 56508 222896
rect 56560 222884 56566 222896
rect 163682 222884 163688 222896
rect 56560 222856 163688 222884
rect 56560 222844 56566 222856
rect 163682 222844 163688 222856
rect 163740 222884 163746 222896
rect 164142 222884 164148 222896
rect 163740 222856 164148 222884
rect 163740 222844 163746 222856
rect 164142 222844 164148 222856
rect 164200 222844 164206 222896
rect 220078 222844 220084 222896
rect 220136 222884 220142 222896
rect 252738 222884 252744 222896
rect 220136 222856 252744 222884
rect 220136 222844 220142 222856
rect 252738 222844 252744 222856
rect 252796 222844 252802 222896
rect 64598 222096 64604 222148
rect 64656 222136 64662 222148
rect 153102 222136 153108 222148
rect 64656 222108 153108 222136
rect 64656 222096 64662 222108
rect 153102 222096 153108 222108
rect 153160 222096 153166 222148
rect 204162 222096 204168 222148
rect 204220 222136 204226 222148
rect 265158 222136 265164 222148
rect 204220 222108 265164 222136
rect 204220 222096 204226 222108
rect 265158 222096 265164 222108
rect 265216 222096 265222 222148
rect 153102 221416 153108 221468
rect 153160 221456 153166 221468
rect 187602 221456 187608 221468
rect 153160 221428 187608 221456
rect 153160 221416 153166 221428
rect 187602 221416 187608 221428
rect 187660 221456 187666 221468
rect 195974 221456 195980 221468
rect 187660 221428 195980 221456
rect 187660 221416 187666 221428
rect 195974 221416 195980 221428
rect 196032 221416 196038 221468
rect 252554 221416 252560 221468
rect 252612 221456 252618 221468
rect 274818 221456 274824 221468
rect 252612 221428 274824 221456
rect 252612 221416 252618 221428
rect 274818 221416 274824 221428
rect 274876 221416 274882 221468
rect 102778 220736 102784 220788
rect 102836 220776 102842 220788
rect 263686 220776 263692 220788
rect 102836 220748 263692 220776
rect 102836 220736 102842 220748
rect 263686 220736 263692 220748
rect 263744 220736 263750 220788
rect 53650 220056 53656 220108
rect 53708 220096 53714 220108
rect 171870 220096 171876 220108
rect 53708 220068 171876 220096
rect 53708 220056 53714 220068
rect 171870 220056 171876 220068
rect 171928 220056 171934 220108
rect 222838 220056 222844 220108
rect 222896 220096 222902 220108
rect 252646 220096 252652 220108
rect 222896 220068 252652 220096
rect 222896 220056 222902 220068
rect 252646 220056 252652 220068
rect 252704 220056 252710 220108
rect 256050 220056 256056 220108
rect 256108 220096 256114 220108
rect 580350 220096 580356 220108
rect 256108 220068 580356 220096
rect 256108 220056 256114 220068
rect 580350 220056 580356 220068
rect 580408 220056 580414 220108
rect 160738 219376 160744 219428
rect 160796 219416 160802 219428
rect 161382 219416 161388 219428
rect 160796 219388 161388 219416
rect 160796 219376 160802 219388
rect 161382 219376 161388 219388
rect 161440 219416 161446 219428
rect 278038 219416 278044 219428
rect 161440 219388 278044 219416
rect 161440 219376 161446 219388
rect 278038 219376 278044 219388
rect 278096 219376 278102 219428
rect 47578 218764 47584 218816
rect 47636 218804 47642 218816
rect 106918 218804 106924 218816
rect 47636 218776 106924 218804
rect 47636 218764 47642 218776
rect 106918 218764 106924 218776
rect 106976 218764 106982 218816
rect 92566 218696 92572 218748
rect 92624 218736 92630 218748
rect 153838 218736 153844 218748
rect 92624 218708 153844 218736
rect 92624 218696 92630 218708
rect 153838 218696 153844 218708
rect 153896 218696 153902 218748
rect 154022 218696 154028 218748
rect 154080 218736 154086 218748
rect 256602 218736 256608 218748
rect 154080 218708 256608 218736
rect 154080 218696 154086 218708
rect 256602 218696 256608 218708
rect 256660 218736 256666 218748
rect 258534 218736 258540 218748
rect 256660 218708 258540 218736
rect 256660 218696 256666 218708
rect 258534 218696 258540 218708
rect 258592 218696 258598 218748
rect 71774 217948 71780 218000
rect 71832 217988 71838 218000
rect 73062 217988 73068 218000
rect 71832 217960 73068 217988
rect 71832 217948 71838 217960
rect 73062 217948 73068 217960
rect 73120 217988 73126 218000
rect 166994 217988 167000 218000
rect 73120 217960 167000 217988
rect 73120 217948 73126 217960
rect 166994 217948 167000 217960
rect 167052 217988 167058 218000
rect 271874 217988 271880 218000
rect 167052 217960 271880 217988
rect 167052 217948 167058 217960
rect 271874 217948 271880 217960
rect 271932 217948 271938 218000
rect 172054 217880 172060 217932
rect 172112 217920 172118 217932
rect 224218 217920 224224 217932
rect 172112 217892 224224 217920
rect 172112 217880 172118 217892
rect 224218 217880 224224 217892
rect 224276 217880 224282 217932
rect 106090 217268 106096 217320
rect 106148 217308 106154 217320
rect 120166 217308 120172 217320
rect 106148 217280 120172 217308
rect 106148 217268 106154 217280
rect 120166 217268 120172 217280
rect 120224 217268 120230 217320
rect 239398 217268 239404 217320
rect 239456 217308 239462 217320
rect 249150 217308 249156 217320
rect 239456 217280 249156 217308
rect 239456 217268 239462 217280
rect 249150 217268 249156 217280
rect 249208 217268 249214 217320
rect 171870 216656 171876 216708
rect 171928 216696 171934 216708
rect 172054 216696 172060 216708
rect 171928 216668 172060 216696
rect 171928 216656 171934 216668
rect 172054 216656 172060 216668
rect 172112 216656 172118 216708
rect 98730 216588 98736 216640
rect 98788 216628 98794 216640
rect 103606 216628 103612 216640
rect 98788 216600 103612 216628
rect 98788 216588 98794 216600
rect 103606 216588 103612 216600
rect 103664 216628 103670 216640
rect 264974 216628 264980 216640
rect 103664 216600 264980 216628
rect 103664 216588 103670 216600
rect 264974 216588 264980 216600
rect 265032 216588 265038 216640
rect 184290 216520 184296 216572
rect 184348 216560 184354 216572
rect 247770 216560 247776 216572
rect 184348 216532 247776 216560
rect 184348 216520 184354 216532
rect 247770 216520 247776 216532
rect 247828 216520 247834 216572
rect 119338 215908 119344 215960
rect 119396 215948 119402 215960
rect 159542 215948 159548 215960
rect 119396 215920 159548 215948
rect 119396 215908 119402 215920
rect 159542 215908 159548 215920
rect 159600 215908 159606 215960
rect 258718 215908 258724 215960
rect 258776 215948 258782 215960
rect 273254 215948 273260 215960
rect 258776 215920 273260 215948
rect 258776 215908 258782 215920
rect 273254 215908 273260 215920
rect 273312 215908 273318 215960
rect 184290 215636 184296 215688
rect 184348 215676 184354 215688
rect 184842 215676 184848 215688
rect 184348 215648 184848 215676
rect 184348 215636 184354 215648
rect 184842 215636 184848 215648
rect 184900 215636 184906 215688
rect 3970 214888 3976 214940
rect 4028 214928 4034 214940
rect 7558 214928 7564 214940
rect 4028 214900 7564 214928
rect 4028 214888 4034 214900
rect 7558 214888 7564 214900
rect 7616 214888 7622 214940
rect 105630 214548 105636 214600
rect 105688 214588 105694 214600
rect 244918 214588 244924 214600
rect 105688 214560 244924 214588
rect 105688 214548 105694 214560
rect 244918 214548 244924 214560
rect 244976 214548 244982 214600
rect 95234 213188 95240 213240
rect 95292 213228 95298 213240
rect 117406 213228 117412 213240
rect 95292 213200 117412 213228
rect 95292 213188 95298 213200
rect 117406 213188 117412 213200
rect 117464 213188 117470 213240
rect 117406 212508 117412 212560
rect 117464 212548 117470 212560
rect 258074 212548 258080 212560
rect 117464 212520 258080 212548
rect 117464 212508 117470 212520
rect 258074 212508 258080 212520
rect 258132 212548 258138 212560
rect 258626 212548 258632 212560
rect 258132 212520 258632 212548
rect 258132 212508 258138 212520
rect 258626 212508 258632 212520
rect 258684 212508 258690 212560
rect 50982 212440 50988 212492
rect 51040 212480 51046 212492
rect 269390 212480 269396 212492
rect 51040 212452 269396 212480
rect 51040 212440 51046 212452
rect 269390 212440 269396 212452
rect 269448 212440 269454 212492
rect 149790 212372 149796 212424
rect 149848 212412 149854 212424
rect 222378 212412 222384 212424
rect 149848 212384 222384 212412
rect 149848 212372 149854 212384
rect 222378 212372 222384 212384
rect 222436 212412 222442 212424
rect 222930 212412 222936 212424
rect 222436 212384 222936 212412
rect 222436 212372 222442 212384
rect 222930 212372 222936 212384
rect 222988 212372 222994 212424
rect 142982 210468 142988 210520
rect 143040 210508 143046 210520
rect 235994 210508 236000 210520
rect 143040 210480 236000 210508
rect 143040 210468 143046 210480
rect 235994 210468 236000 210480
rect 236052 210468 236058 210520
rect 78582 210400 78588 210452
rect 78640 210440 78646 210452
rect 106918 210440 106924 210452
rect 78640 210412 106924 210440
rect 78640 210400 78646 210412
rect 106918 210400 106924 210412
rect 106976 210440 106982 210452
rect 257338 210440 257344 210452
rect 106976 210412 257344 210440
rect 106976 210400 106982 210412
rect 257338 210400 257344 210412
rect 257396 210400 257402 210452
rect 173802 209720 173808 209772
rect 173860 209760 173866 209772
rect 278958 209760 278964 209772
rect 173860 209732 278964 209760
rect 173860 209720 173866 209732
rect 278958 209720 278964 209732
rect 279016 209720 279022 209772
rect 97350 209108 97356 209160
rect 97408 209148 97414 209160
rect 108114 209148 108120 209160
rect 97408 209120 108120 209148
rect 97408 209108 97414 209120
rect 108114 209108 108120 209120
rect 108172 209108 108178 209160
rect 57698 209040 57704 209092
rect 57756 209080 57762 209092
rect 173802 209080 173808 209092
rect 57756 209052 173808 209080
rect 57756 209040 57762 209052
rect 173802 209040 173808 209052
rect 173860 209040 173866 209092
rect 107746 208360 107752 208412
rect 107804 208400 107810 208412
rect 108114 208400 108120 208412
rect 107804 208372 108120 208400
rect 107804 208360 107810 208372
rect 108114 208360 108120 208372
rect 108172 208400 108178 208412
rect 263594 208400 263600 208412
rect 108172 208372 263600 208400
rect 108172 208360 108178 208372
rect 263594 208360 263600 208372
rect 263652 208400 263658 208412
rect 263962 208400 263968 208412
rect 263652 208372 263968 208400
rect 263652 208360 263658 208372
rect 263962 208360 263968 208372
rect 264020 208360 264026 208412
rect 86954 207680 86960 207732
rect 87012 207720 87018 207732
rect 103606 207720 103612 207732
rect 87012 207692 103612 207720
rect 87012 207680 87018 207692
rect 103606 207680 103612 207692
rect 103664 207720 103670 207732
rect 104802 207720 104808 207732
rect 103664 207692 104808 207720
rect 103664 207680 103670 207692
rect 104802 207680 104808 207692
rect 104860 207680 104866 207732
rect 13814 207612 13820 207664
rect 13872 207652 13878 207664
rect 189074 207652 189080 207664
rect 13872 207624 189080 207652
rect 13872 207612 13878 207624
rect 189074 207612 189080 207624
rect 189132 207612 189138 207664
rect 104802 207000 104808 207052
rect 104860 207040 104866 207052
rect 269298 207040 269304 207052
rect 104860 207012 269304 207040
rect 104860 207000 104866 207012
rect 269298 207000 269304 207012
rect 269356 207000 269362 207052
rect 96614 206320 96620 206372
rect 96672 206360 96678 206372
rect 109218 206360 109224 206372
rect 96672 206332 109224 206360
rect 96672 206320 96678 206332
rect 109218 206320 109224 206332
rect 109276 206320 109282 206372
rect 84102 206252 84108 206304
rect 84160 206292 84166 206304
rect 113266 206292 113272 206304
rect 84160 206264 113272 206292
rect 84160 206252 84166 206264
rect 113266 206252 113272 206264
rect 113324 206292 113330 206304
rect 113910 206292 113916 206304
rect 113324 206264 113916 206292
rect 113324 206252 113330 206264
rect 113910 206252 113916 206264
rect 113968 206252 113974 206304
rect 227714 206252 227720 206304
rect 227772 206292 227778 206304
rect 270678 206292 270684 206304
rect 227772 206264 270684 206292
rect 227772 206252 227778 206264
rect 270678 206252 270684 206264
rect 270736 206252 270742 206304
rect 109218 205708 109224 205760
rect 109276 205748 109282 205760
rect 227714 205748 227720 205760
rect 109276 205720 227720 205748
rect 109276 205708 109282 205720
rect 227714 205708 227720 205720
rect 227772 205708 227778 205760
rect 113910 205640 113916 205692
rect 113968 205680 113974 205692
rect 260926 205680 260932 205692
rect 113968 205652 260932 205680
rect 113968 205640 113974 205652
rect 260926 205640 260932 205652
rect 260984 205640 260990 205692
rect 77294 204892 77300 204944
rect 77352 204932 77358 204944
rect 109126 204932 109132 204944
rect 77352 204904 109132 204932
rect 77352 204892 77358 204904
rect 109126 204892 109132 204904
rect 109184 204892 109190 204944
rect 255958 204892 255964 204944
rect 256016 204932 256022 204944
rect 265066 204932 265072 204944
rect 256016 204904 265072 204932
rect 256016 204892 256022 204904
rect 265066 204892 265072 204904
rect 265124 204892 265130 204944
rect 159542 204212 159548 204264
rect 159600 204252 159606 204264
rect 292666 204252 292672 204264
rect 159600 204224 292672 204252
rect 159600 204212 159606 204224
rect 292666 204212 292672 204224
rect 292724 204212 292730 204264
rect 203518 203532 203524 203584
rect 203576 203572 203582 203584
rect 281810 203572 281816 203584
rect 203576 203544 281816 203572
rect 203576 203532 203582 203544
rect 281810 203532 281816 203544
rect 281868 203532 281874 203584
rect 98086 202784 98092 202836
rect 98144 202824 98150 202836
rect 98822 202824 98828 202836
rect 98144 202796 98828 202824
rect 98144 202784 98150 202796
rect 98822 202784 98828 202796
rect 98880 202784 98886 202836
rect 3326 202172 3332 202224
rect 3384 202212 3390 202224
rect 98086 202212 98092 202224
rect 3384 202184 98092 202212
rect 3384 202172 3390 202184
rect 98086 202172 98092 202184
rect 98144 202172 98150 202224
rect 175090 202172 175096 202224
rect 175148 202212 175154 202224
rect 209130 202212 209136 202224
rect 175148 202184 209136 202212
rect 175148 202172 175154 202184
rect 209130 202172 209136 202184
rect 209188 202172 209194 202224
rect 38654 202104 38660 202156
rect 38712 202144 38718 202156
rect 182818 202144 182824 202156
rect 38712 202116 182824 202144
rect 38712 202104 38718 202116
rect 182818 202104 182824 202116
rect 182876 202104 182882 202156
rect 192570 202104 192576 202156
rect 192628 202144 192634 202156
rect 228358 202144 228364 202156
rect 192628 202116 228364 202144
rect 192628 202104 192634 202116
rect 228358 202104 228364 202116
rect 228416 202104 228422 202156
rect 54938 201424 54944 201476
rect 54996 201464 55002 201476
rect 291286 201464 291292 201476
rect 54996 201436 291292 201464
rect 54996 201424 55002 201436
rect 291286 201424 291292 201436
rect 291344 201424 291350 201476
rect 243538 200744 243544 200796
rect 243596 200784 243602 200796
rect 268378 200784 268384 200796
rect 243596 200756 268384 200784
rect 243596 200744 243602 200756
rect 268378 200744 268384 200756
rect 268436 200744 268442 200796
rect 249702 199384 249708 199436
rect 249760 199424 249766 199436
rect 293954 199424 293960 199436
rect 249760 199396 293960 199424
rect 249760 199384 249766 199396
rect 293954 199384 293960 199396
rect 294012 199384 294018 199436
rect 129090 198636 129096 198688
rect 129148 198676 129154 198688
rect 256694 198676 256700 198688
rect 129148 198648 256700 198676
rect 129148 198636 129154 198648
rect 256694 198636 256700 198648
rect 256752 198636 256758 198688
rect 195238 197956 195244 198008
rect 195296 197996 195302 198008
rect 280338 197996 280344 198008
rect 195296 197968 280344 197996
rect 195296 197956 195302 197968
rect 280338 197956 280344 197968
rect 280396 197956 280402 198008
rect 23474 196596 23480 196648
rect 23532 196636 23538 196648
rect 187050 196636 187056 196648
rect 23532 196608 187056 196636
rect 23532 196596 23538 196608
rect 187050 196596 187056 196608
rect 187108 196596 187114 196648
rect 200022 196596 200028 196648
rect 200080 196636 200086 196648
rect 582466 196636 582472 196648
rect 200080 196608 582472 196636
rect 200080 196596 200086 196608
rect 582466 196596 582472 196608
rect 582524 196596 582530 196648
rect 244918 195916 244924 195968
rect 244976 195956 244982 195968
rect 272518 195956 272524 195968
rect 244976 195928 272524 195956
rect 244976 195916 244982 195928
rect 272518 195916 272524 195928
rect 272576 195916 272582 195968
rect 90358 195236 90364 195288
rect 90416 195276 90422 195288
rect 129090 195276 129096 195288
rect 90416 195248 129096 195276
rect 90416 195236 90422 195248
rect 129090 195236 129096 195248
rect 129148 195236 129154 195288
rect 137370 195236 137376 195288
rect 137428 195276 137434 195288
rect 150434 195276 150440 195288
rect 137428 195248 150440 195276
rect 137428 195236 137434 195248
rect 150434 195236 150440 195248
rect 150492 195236 150498 195288
rect 164970 195236 164976 195288
rect 165028 195276 165034 195288
rect 196618 195276 196624 195288
rect 165028 195248 196624 195276
rect 165028 195236 165034 195248
rect 196618 195236 196624 195248
rect 196676 195236 196682 195288
rect 272518 195236 272524 195288
rect 272576 195276 272582 195288
rect 579982 195276 579988 195288
rect 272576 195248 579988 195276
rect 272576 195236 272582 195248
rect 579982 195236 579988 195248
rect 580040 195236 580046 195288
rect 162670 194488 162676 194540
rect 162728 194528 162734 194540
rect 170398 194528 170404 194540
rect 162728 194500 170404 194528
rect 162728 194488 162734 194500
rect 170398 194488 170404 194500
rect 170456 194488 170462 194540
rect 131758 193876 131764 193928
rect 131816 193916 131822 193928
rect 145558 193916 145564 193928
rect 131816 193888 145564 193916
rect 131816 193876 131822 193888
rect 145558 193876 145564 193888
rect 145616 193876 145622 193928
rect 61838 193808 61844 193860
rect 61896 193848 61902 193860
rect 69014 193848 69020 193860
rect 61896 193820 69020 193848
rect 61896 193808 61902 193820
rect 69014 193808 69020 193820
rect 69072 193808 69078 193860
rect 123478 193808 123484 193860
rect 123536 193848 123542 193860
rect 137462 193848 137468 193860
rect 123536 193820 137468 193848
rect 123536 193808 123542 193820
rect 137462 193808 137468 193820
rect 137520 193808 137526 193860
rect 138658 193808 138664 193860
rect 138716 193848 138722 193860
rect 148502 193848 148508 193860
rect 138716 193820 148508 193848
rect 138716 193808 138722 193820
rect 148502 193808 148508 193820
rect 148560 193808 148566 193860
rect 170490 193808 170496 193860
rect 170548 193848 170554 193860
rect 189718 193848 189724 193860
rect 170548 193820 189724 193848
rect 170548 193808 170554 193820
rect 189718 193808 189724 193820
rect 189776 193808 189782 193860
rect 49694 189728 49700 189780
rect 49752 189768 49758 189780
rect 193306 189768 193312 189780
rect 49752 189740 193312 189768
rect 49752 189728 49758 189740
rect 193306 189728 193312 189740
rect 193364 189728 193370 189780
rect 213178 189728 213184 189780
rect 213236 189768 213242 189780
rect 295426 189768 295432 189780
rect 213236 189740 295432 189768
rect 213236 189728 213242 189740
rect 295426 189728 295432 189740
rect 295484 189728 295490 189780
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 43438 189020 43444 189032
rect 3476 188992 43444 189020
rect 3476 188980 3482 188992
rect 43438 188980 43444 188992
rect 43496 188980 43502 189032
rect 232498 188300 232504 188352
rect 232556 188340 232562 188352
rect 276290 188340 276296 188352
rect 232556 188312 276296 188340
rect 232556 188300 232562 188312
rect 276290 188300 276296 188312
rect 276348 188300 276354 188352
rect 48314 186940 48320 186992
rect 48372 186980 48378 186992
rect 120810 186980 120816 186992
rect 48372 186952 120816 186980
rect 48372 186940 48378 186952
rect 120810 186940 120816 186952
rect 120868 186940 120874 186992
rect 195330 186940 195336 186992
rect 195388 186980 195394 186992
rect 226334 186980 226340 186992
rect 195388 186952 226340 186980
rect 195388 186940 195394 186952
rect 226334 186940 226340 186952
rect 226392 186940 226398 186992
rect 133138 185648 133144 185700
rect 133196 185688 133202 185700
rect 147122 185688 147128 185700
rect 133196 185660 147128 185688
rect 133196 185648 133202 185660
rect 147122 185648 147128 185660
rect 147180 185648 147186 185700
rect 45462 185580 45468 185632
rect 45520 185620 45526 185632
rect 73430 185620 73436 185632
rect 45520 185592 73436 185620
rect 45520 185580 45526 185592
rect 73430 185580 73436 185592
rect 73488 185580 73494 185632
rect 118786 185580 118792 185632
rect 118844 185620 118850 185632
rect 138750 185620 138756 185632
rect 118844 185592 138756 185620
rect 118844 185580 118850 185592
rect 138750 185580 138756 185592
rect 138808 185580 138814 185632
rect 145558 184968 145564 185020
rect 145616 185008 145622 185020
rect 153930 185008 153936 185020
rect 145616 184980 153936 185008
rect 145616 184968 145622 184980
rect 153930 184968 153936 184980
rect 153988 184968 153994 185020
rect 195330 184152 195336 184204
rect 195388 184192 195394 184204
rect 249058 184192 249064 184204
rect 195388 184164 249064 184192
rect 195388 184152 195394 184164
rect 249058 184152 249064 184164
rect 249116 184152 249122 184204
rect 122098 182860 122104 182912
rect 122156 182900 122162 182912
rect 134702 182900 134708 182912
rect 122156 182872 134708 182900
rect 122156 182860 122162 182872
rect 134702 182860 134708 182872
rect 134760 182860 134766 182912
rect 89530 182792 89536 182844
rect 89588 182832 89594 182844
rect 124306 182832 124312 182844
rect 89588 182804 124312 182832
rect 89588 182792 89594 182804
rect 124306 182792 124312 182804
rect 124364 182792 124370 182844
rect 69658 180820 69664 180872
rect 69716 180860 69722 180872
rect 175918 180860 175924 180872
rect 69716 180832 175924 180860
rect 69716 180820 69722 180832
rect 175918 180820 175924 180832
rect 175976 180820 175982 180872
rect 214558 180140 214564 180192
rect 214616 180180 214622 180192
rect 224954 180180 224960 180192
rect 214616 180152 224960 180180
rect 214616 180140 214622 180152
rect 224954 180140 224960 180152
rect 225012 180140 225018 180192
rect 91002 180072 91008 180124
rect 91060 180112 91066 180124
rect 107654 180112 107660 180124
rect 91060 180084 107660 180112
rect 91060 180072 91066 180084
rect 107654 180072 107660 180084
rect 107712 180072 107718 180124
rect 122834 180072 122840 180124
rect 122892 180112 122898 180124
rect 140130 180112 140136 180124
rect 122892 180084 140136 180112
rect 122892 180072 122898 180084
rect 140130 180072 140136 180084
rect 140188 180072 140194 180124
rect 207750 180072 207756 180124
rect 207808 180112 207814 180124
rect 287238 180112 287244 180124
rect 207808 180084 287244 180112
rect 207808 180072 207814 180084
rect 287238 180072 287244 180084
rect 287296 180072 287302 180124
rect 191098 179732 191104 179784
rect 191156 179772 191162 179784
rect 198918 179772 198924 179784
rect 191156 179744 198924 179772
rect 191156 179732 191162 179744
rect 198918 179732 198924 179744
rect 198976 179732 198982 179784
rect 1394 178644 1400 178696
rect 1452 178684 1458 178696
rect 145650 178684 145656 178696
rect 1452 178656 145656 178684
rect 1452 178644 1458 178656
rect 145650 178644 145656 178656
rect 145708 178644 145714 178696
rect 197998 178644 198004 178696
rect 198056 178684 198062 178696
rect 234614 178684 234620 178696
rect 198056 178656 234620 178684
rect 198056 178644 198062 178656
rect 234614 178644 234620 178656
rect 234672 178644 234678 178696
rect 241422 178644 241428 178696
rect 241480 178684 241486 178696
rect 580166 178684 580172 178696
rect 241480 178656 580172 178684
rect 241480 178644 241486 178656
rect 580166 178644 580172 178656
rect 580224 178644 580230 178696
rect 240778 178032 240784 178084
rect 240836 178072 240842 178084
rect 241422 178072 241428 178084
rect 240836 178044 241428 178072
rect 240836 178032 240842 178044
rect 241422 178032 241428 178044
rect 241480 178032 241486 178084
rect 85482 177284 85488 177336
rect 85540 177324 85546 177336
rect 213178 177324 213184 177336
rect 85540 177296 213184 177324
rect 85540 177284 85546 177296
rect 213178 177284 213184 177296
rect 213236 177284 213242 177336
rect 228358 177284 228364 177336
rect 228416 177324 228422 177336
rect 251818 177324 251824 177336
rect 228416 177296 251824 177324
rect 228416 177284 228422 177296
rect 251818 177284 251824 177296
rect 251876 177284 251882 177336
rect 84194 176672 84200 176724
rect 84252 176712 84258 176724
rect 85482 176712 85488 176724
rect 84252 176684 85488 176712
rect 84252 176672 84258 176684
rect 85482 176672 85488 176684
rect 85540 176672 85546 176724
rect 93118 176672 93124 176724
rect 93176 176712 93182 176724
rect 93670 176712 93676 176724
rect 93176 176684 93676 176712
rect 93176 176672 93182 176684
rect 93670 176672 93676 176684
rect 93728 176712 93734 176724
rect 220078 176712 220084 176724
rect 93728 176684 220084 176712
rect 93728 176672 93734 176684
rect 220078 176672 220084 176684
rect 220136 176672 220142 176724
rect 88978 175924 88984 175976
rect 89036 175964 89042 175976
rect 121546 175964 121552 175976
rect 89036 175936 121552 175964
rect 89036 175924 89042 175936
rect 121546 175924 121552 175936
rect 121604 175964 121610 175976
rect 214006 175964 214012 175976
rect 121604 175936 214012 175964
rect 121604 175924 121610 175936
rect 214006 175924 214012 175936
rect 214064 175924 214070 175976
rect 214006 175244 214012 175296
rect 214064 175284 214070 175296
rect 247678 175284 247684 175296
rect 214064 175256 247684 175284
rect 214064 175244 214070 175256
rect 247678 175244 247684 175256
rect 247736 175244 247742 175296
rect 255314 175244 255320 175296
rect 255372 175284 255378 175296
rect 256602 175284 256608 175296
rect 255372 175256 256608 175284
rect 255372 175244 255378 175256
rect 256602 175244 256608 175256
rect 256660 175284 256666 175296
rect 583018 175284 583024 175296
rect 256660 175256 583024 175284
rect 256660 175244 256666 175256
rect 583018 175244 583024 175256
rect 583076 175244 583082 175296
rect 196066 175176 196072 175228
rect 196124 175216 196130 175228
rect 196802 175216 196808 175228
rect 196124 175188 196808 175216
rect 196124 175176 196130 175188
rect 196802 175176 196808 175188
rect 196860 175176 196866 175228
rect 205726 174700 205732 174752
rect 205784 174740 205790 174752
rect 206278 174740 206284 174752
rect 205784 174712 206284 174740
rect 205784 174700 205790 174712
rect 206278 174700 206284 174712
rect 206336 174700 206342 174752
rect 82078 174496 82084 174548
rect 82136 174536 82142 174548
rect 82722 174536 82728 174548
rect 82136 174508 82728 174536
rect 82136 174496 82142 174508
rect 82722 174496 82728 174508
rect 82780 174536 82786 174548
rect 205726 174536 205732 174548
rect 82780 174508 205732 174536
rect 82780 174496 82786 174508
rect 205726 174496 205732 174508
rect 205784 174496 205790 174548
rect 88334 173884 88340 173936
rect 88392 173924 88398 173936
rect 196802 173924 196808 173936
rect 88392 173896 196808 173924
rect 88392 173884 88398 173896
rect 196802 173884 196808 173896
rect 196860 173884 196866 173936
rect 137462 172592 137468 172644
rect 137520 172632 137526 172644
rect 228358 172632 228364 172644
rect 137520 172604 228364 172632
rect 137520 172592 137526 172604
rect 228358 172592 228364 172604
rect 228416 172592 228422 172644
rect 205726 172524 205732 172576
rect 205784 172564 205790 172576
rect 320174 172564 320180 172576
rect 205784 172536 320180 172564
rect 205784 172524 205790 172536
rect 320174 172524 320180 172536
rect 320232 172524 320238 172576
rect 85574 171844 85580 171896
rect 85632 171884 85638 171896
rect 106274 171884 106280 171896
rect 85632 171856 106280 171884
rect 85632 171844 85638 171856
rect 106274 171844 106280 171856
rect 106332 171844 106338 171896
rect 91002 171776 91008 171828
rect 91060 171816 91066 171828
rect 180150 171816 180156 171828
rect 91060 171788 180156 171816
rect 91060 171776 91066 171788
rect 180150 171776 180156 171788
rect 180208 171816 180214 171828
rect 221458 171816 221464 171828
rect 180208 171788 221464 171816
rect 180208 171776 180214 171788
rect 221458 171776 221464 171788
rect 221516 171776 221522 171828
rect 237374 171776 237380 171828
rect 237432 171816 237438 171828
rect 256694 171816 256700 171828
rect 237432 171788 256700 171816
rect 237432 171776 237438 171788
rect 256694 171776 256700 171788
rect 256752 171776 256758 171828
rect 112438 171096 112444 171148
rect 112496 171136 112502 171148
rect 230566 171136 230572 171148
rect 112496 171108 230572 171136
rect 112496 171096 112502 171108
rect 230566 171096 230572 171108
rect 230624 171096 230630 171148
rect 194870 170620 194876 170672
rect 194928 170660 194934 170672
rect 195330 170660 195336 170672
rect 194928 170632 195336 170660
rect 194928 170620 194934 170632
rect 195330 170620 195336 170632
rect 195388 170620 195394 170672
rect 56318 170348 56324 170400
rect 56376 170388 56382 170400
rect 194870 170388 194876 170400
rect 56376 170360 194876 170388
rect 56376 170348 56382 170360
rect 194870 170348 194876 170360
rect 194928 170348 194934 170400
rect 196710 170348 196716 170400
rect 196768 170388 196774 170400
rect 205634 170388 205640 170400
rect 196768 170360 205640 170388
rect 196768 170348 196774 170360
rect 205634 170348 205640 170360
rect 205692 170348 205698 170400
rect 215386 170348 215392 170400
rect 215444 170388 215450 170400
rect 259454 170388 259460 170400
rect 215444 170360 259460 170388
rect 215444 170348 215450 170360
rect 259454 170348 259460 170360
rect 259512 170348 259518 170400
rect 115290 169736 115296 169788
rect 115348 169776 115354 169788
rect 204714 169776 204720 169788
rect 115348 169748 204720 169776
rect 115348 169736 115354 169748
rect 204714 169736 204720 169748
rect 204772 169736 204778 169788
rect 262674 168988 262680 169040
rect 262732 169028 262738 169040
rect 276198 169028 276204 169040
rect 262732 169000 276204 169028
rect 262732 168988 262738 169000
rect 276198 168988 276204 169000
rect 276256 168988 276262 169040
rect 87690 168444 87696 168496
rect 87748 168484 87754 168496
rect 200666 168484 200672 168496
rect 87748 168456 200672 168484
rect 87748 168444 87754 168456
rect 200666 168444 200672 168456
rect 200724 168444 200730 168496
rect 204254 168444 204260 168496
rect 204312 168484 204318 168496
rect 204714 168484 204720 168496
rect 204312 168456 204720 168484
rect 204312 168444 204318 168456
rect 204714 168444 204720 168456
rect 204772 168484 204778 168496
rect 262306 168484 262312 168496
rect 204772 168456 262312 168484
rect 204772 168444 204778 168456
rect 262306 168444 262312 168456
rect 262364 168484 262370 168496
rect 262674 168484 262680 168496
rect 262364 168456 262680 168484
rect 262364 168444 262370 168456
rect 262674 168444 262680 168456
rect 262732 168444 262738 168496
rect 92658 168376 92664 168428
rect 92716 168416 92722 168428
rect 222194 168416 222200 168428
rect 92716 168388 222200 168416
rect 92716 168376 92722 168388
rect 222194 168376 222200 168388
rect 222252 168416 222258 168428
rect 222838 168416 222844 168428
rect 222252 168388 222844 168416
rect 222252 168376 222258 168388
rect 222838 168376 222844 168388
rect 222896 168376 222902 168428
rect 76742 167628 76748 167680
rect 76800 167668 76806 167680
rect 202874 167668 202880 167680
rect 76800 167640 202880 167668
rect 76800 167628 76806 167640
rect 202874 167628 202880 167640
rect 202932 167668 202938 167680
rect 203518 167668 203524 167680
rect 202932 167640 203524 167668
rect 202932 167628 202938 167640
rect 203518 167628 203524 167640
rect 203576 167628 203582 167680
rect 222286 167628 222292 167680
rect 222344 167668 222350 167680
rect 238018 167668 238024 167680
rect 222344 167640 238024 167668
rect 222344 167628 222350 167640
rect 238018 167628 238024 167640
rect 238076 167628 238082 167680
rect 75914 167016 75920 167068
rect 75972 167056 75978 167068
rect 76742 167056 76748 167068
rect 75972 167028 76748 167056
rect 75972 167016 75978 167028
rect 76742 167016 76748 167028
rect 76800 167016 76806 167068
rect 195974 167016 195980 167068
rect 196032 167056 196038 167068
rect 196618 167056 196624 167068
rect 196032 167028 196624 167056
rect 196032 167016 196038 167028
rect 196618 167016 196624 167028
rect 196676 167056 196682 167068
rect 303614 167056 303620 167068
rect 196676 167028 303620 167056
rect 196676 167016 196682 167028
rect 303614 167016 303620 167028
rect 303672 167016 303678 167068
rect 169110 165656 169116 165708
rect 169168 165696 169174 165708
rect 224218 165696 224224 165708
rect 169168 165668 224224 165696
rect 169168 165656 169174 165668
rect 224218 165656 224224 165668
rect 224276 165656 224282 165708
rect 82906 165588 82912 165640
rect 82964 165628 82970 165640
rect 204990 165628 204996 165640
rect 82964 165600 204996 165628
rect 82964 165588 82970 165600
rect 204990 165588 204996 165600
rect 205048 165588 205054 165640
rect 199378 164840 199384 164892
rect 199436 164880 199442 164892
rect 260834 164880 260840 164892
rect 199436 164852 260840 164880
rect 199436 164840 199442 164852
rect 260834 164840 260840 164852
rect 260892 164840 260898 164892
rect 65886 164296 65892 164348
rect 65944 164336 65950 164348
rect 154022 164336 154028 164348
rect 65944 164308 154028 164336
rect 65944 164296 65950 164308
rect 154022 164296 154028 164308
rect 154080 164296 154086 164348
rect 82170 164228 82176 164280
rect 82228 164268 82234 164280
rect 208394 164268 208400 164280
rect 82228 164240 208400 164268
rect 82228 164228 82234 164240
rect 208394 164228 208400 164240
rect 208452 164228 208458 164280
rect 224770 163480 224776 163532
rect 224828 163520 224834 163532
rect 283098 163520 283104 163532
rect 224828 163492 283104 163520
rect 224828 163480 224834 163492
rect 283098 163480 283104 163492
rect 283156 163480 283162 163532
rect 60550 162936 60556 162988
rect 60608 162976 60614 162988
rect 152642 162976 152648 162988
rect 60608 162948 152648 162976
rect 60608 162936 60614 162948
rect 152642 162936 152648 162948
rect 152700 162936 152706 162988
rect 2866 162868 2872 162920
rect 2924 162908 2930 162920
rect 4798 162908 4804 162920
rect 2924 162880 4804 162908
rect 2924 162868 2930 162880
rect 4798 162868 4804 162880
rect 4856 162868 4862 162920
rect 92474 162868 92480 162920
rect 92532 162908 92538 162920
rect 222286 162908 222292 162920
rect 92532 162880 222292 162908
rect 92532 162868 92538 162880
rect 222286 162868 222292 162880
rect 222344 162868 222350 162920
rect 133230 161984 133236 162036
rect 133288 162024 133294 162036
rect 133690 162024 133696 162036
rect 133288 161996 133696 162024
rect 133288 161984 133294 161996
rect 133690 161984 133696 161996
rect 133748 161984 133754 162036
rect 133230 161508 133236 161560
rect 133288 161548 133294 161560
rect 226518 161548 226524 161560
rect 133288 161520 226524 161548
rect 133288 161508 133294 161520
rect 226518 161508 226524 161520
rect 226576 161508 226582 161560
rect 87138 161440 87144 161492
rect 87196 161480 87202 161492
rect 215386 161480 215392 161492
rect 87196 161452 215392 161480
rect 87196 161440 87202 161452
rect 215386 161440 215392 161452
rect 215444 161440 215450 161492
rect 231118 160760 231124 160812
rect 231176 160800 231182 160812
rect 274726 160800 274732 160812
rect 231176 160772 274732 160800
rect 231176 160760 231182 160772
rect 274726 160760 274732 160772
rect 274784 160760 274790 160812
rect 97902 160692 97908 160744
rect 97960 160732 97966 160744
rect 249794 160732 249800 160744
rect 97960 160704 249800 160732
rect 97960 160692 97966 160704
rect 249794 160692 249800 160704
rect 249852 160692 249858 160744
rect 97350 160148 97356 160200
rect 97408 160188 97414 160200
rect 97902 160188 97908 160200
rect 97408 160160 97908 160188
rect 97408 160148 97414 160160
rect 97902 160148 97908 160160
rect 97960 160148 97966 160200
rect 91738 160080 91744 160132
rect 91796 160120 91802 160132
rect 92290 160120 92296 160132
rect 91796 160092 92296 160120
rect 91796 160080 91802 160092
rect 92290 160080 92296 160092
rect 92348 160120 92354 160132
rect 218790 160120 218796 160132
rect 92348 160092 218796 160120
rect 92348 160080 92354 160092
rect 218790 160080 218796 160092
rect 218848 160080 218854 160132
rect 249610 159400 249616 159452
rect 249668 159440 249674 159452
rect 249668 159412 277394 159440
rect 249668 159400 249674 159412
rect 202782 159332 202788 159384
rect 202840 159372 202846 159384
rect 269206 159372 269212 159384
rect 202840 159344 269212 159372
rect 202840 159332 202846 159344
rect 269206 159332 269212 159344
rect 269264 159332 269270 159384
rect 277366 159372 277394 159412
rect 278866 159372 278872 159384
rect 277366 159344 278872 159372
rect 278866 159332 278872 159344
rect 278924 159372 278930 159384
rect 338758 159372 338764 159384
rect 278924 159344 338764 159372
rect 278924 159332 278930 159344
rect 338758 159332 338764 159344
rect 338816 159332 338822 159384
rect 198734 159196 198740 159248
rect 198792 159236 198798 159248
rect 199378 159236 199384 159248
rect 198792 159208 199384 159236
rect 198792 159196 198798 159208
rect 199378 159196 199384 159208
rect 199436 159196 199442 159248
rect 72970 158788 72976 158840
rect 73028 158828 73034 158840
rect 198734 158828 198740 158840
rect 73028 158800 198740 158828
rect 73028 158788 73034 158800
rect 198734 158788 198740 158800
rect 198792 158788 198798 158840
rect 91830 158720 91836 158772
rect 91888 158760 91894 158772
rect 92382 158760 92388 158772
rect 91888 158732 92388 158760
rect 91888 158720 91894 158732
rect 92382 158720 92388 158732
rect 92440 158760 92446 158772
rect 220998 158760 221004 158772
rect 92440 158732 221004 158760
rect 92440 158720 92446 158732
rect 220998 158720 221004 158732
rect 221056 158720 221062 158772
rect 192478 158652 192484 158704
rect 192536 158692 192542 158704
rect 249610 158692 249616 158704
rect 192536 158664 249616 158692
rect 192536 158652 192542 158664
rect 249610 158652 249616 158664
rect 249668 158652 249674 158704
rect 56410 157972 56416 158024
rect 56468 158012 56474 158024
rect 74626 158012 74632 158024
rect 56468 157984 74632 158012
rect 56468 157972 56474 157984
rect 74626 157972 74632 157984
rect 74684 157972 74690 158024
rect 76558 157972 76564 158024
rect 76616 158012 76622 158024
rect 107010 158012 107016 158024
rect 76616 157984 107016 158012
rect 76616 157972 76622 157984
rect 107010 157972 107016 157984
rect 107068 157972 107074 158024
rect 154022 157972 154028 158024
rect 154080 158012 154086 158024
rect 187694 158012 187700 158024
rect 154080 157984 187700 158012
rect 154080 157972 154086 157984
rect 187694 157972 187700 157984
rect 187752 157972 187758 158024
rect 97994 157360 98000 157412
rect 98052 157400 98058 157412
rect 98822 157400 98828 157412
rect 98052 157372 98828 157400
rect 98052 157360 98058 157372
rect 98822 157360 98828 157372
rect 98880 157400 98886 157412
rect 227714 157400 227720 157412
rect 98880 157372 227720 157400
rect 98880 157360 98886 157372
rect 227714 157360 227720 157372
rect 227772 157360 227778 157412
rect 187694 157292 187700 157344
rect 187752 157332 187758 157344
rect 188890 157332 188896 157344
rect 187752 157304 188896 157332
rect 187752 157292 187758 157304
rect 188890 157292 188896 157304
rect 188948 157332 188954 157344
rect 214650 157332 214656 157344
rect 188948 157304 214656 157332
rect 188948 157292 188954 157304
rect 214650 157292 214656 157304
rect 214708 157292 214714 157344
rect 35802 156612 35808 156664
rect 35860 156652 35866 156664
rect 67726 156652 67732 156664
rect 35860 156624 67732 156652
rect 35860 156612 35866 156624
rect 67726 156612 67732 156624
rect 67784 156652 67790 156664
rect 68922 156652 68928 156664
rect 67784 156624 68928 156652
rect 67784 156612 67790 156624
rect 68922 156612 68928 156624
rect 68980 156612 68986 156664
rect 68922 156000 68928 156052
rect 68980 156040 68986 156052
rect 188430 156040 188436 156052
rect 68980 156012 188436 156040
rect 68980 156000 68986 156012
rect 188430 156000 188436 156012
rect 188488 156000 188494 156052
rect 210510 156000 210516 156052
rect 210568 156040 210574 156052
rect 210970 156040 210976 156052
rect 210568 156012 210976 156040
rect 210568 156000 210574 156012
rect 210970 156000 210976 156012
rect 211028 156040 211034 156052
rect 229094 156040 229100 156052
rect 211028 156012 229100 156040
rect 211028 156000 211034 156012
rect 229094 156000 229100 156012
rect 229152 156000 229158 156052
rect 75178 155932 75184 155984
rect 75236 155972 75242 155984
rect 201678 155972 201684 155984
rect 75236 155944 201684 155972
rect 75236 155932 75242 155944
rect 201678 155932 201684 155944
rect 201736 155972 201742 155984
rect 202782 155972 202788 155984
rect 201736 155944 202788 155972
rect 201736 155932 201742 155944
rect 202782 155932 202788 155944
rect 202840 155932 202846 155984
rect 218054 155932 218060 155984
rect 218112 155972 218118 155984
rect 218882 155972 218888 155984
rect 218112 155944 218888 155972
rect 218112 155932 218118 155944
rect 218882 155932 218888 155944
rect 218940 155972 218946 155984
rect 246390 155972 246396 155984
rect 218940 155944 246396 155972
rect 218940 155932 218946 155944
rect 246390 155932 246396 155944
rect 246448 155932 246454 155984
rect 60458 155864 60464 155916
rect 60516 155904 60522 155916
rect 60642 155904 60648 155916
rect 60516 155876 60648 155904
rect 60516 155864 60522 155876
rect 60642 155864 60648 155876
rect 60700 155864 60706 155916
rect 294690 155184 294696 155236
rect 294748 155224 294754 155236
rect 583110 155224 583116 155236
rect 294748 155196 583116 155224
rect 294748 155184 294754 155196
rect 583110 155184 583116 155196
rect 583168 155184 583174 155236
rect 60458 154640 60464 154692
rect 60516 154680 60522 154692
rect 154022 154680 154028 154692
rect 60516 154652 154028 154680
rect 60516 154640 60522 154652
rect 154022 154640 154028 154652
rect 154080 154640 154086 154692
rect 158714 154640 158720 154692
rect 158772 154680 158778 154692
rect 160002 154680 160008 154692
rect 158772 154652 160008 154680
rect 158772 154640 158778 154652
rect 160002 154640 160008 154652
rect 160060 154680 160066 154692
rect 186958 154680 186964 154692
rect 160060 154652 186964 154680
rect 160060 154640 160066 154652
rect 186958 154640 186964 154652
rect 187016 154640 187022 154692
rect 187694 154640 187700 154692
rect 187752 154680 187758 154692
rect 224954 154680 224960 154692
rect 187752 154652 224960 154680
rect 187752 154640 187758 154652
rect 224954 154640 224960 154652
rect 225012 154640 225018 154692
rect 88610 154572 88616 154624
rect 88668 154612 88674 154624
rect 218698 154612 218704 154624
rect 88668 154584 218704 154612
rect 88668 154572 88674 154584
rect 218698 154572 218704 154584
rect 218756 154572 218762 154624
rect 93854 153892 93860 153944
rect 93912 153932 93918 153944
rect 131114 153932 131120 153944
rect 93912 153904 131120 153932
rect 93912 153892 93918 153904
rect 131114 153892 131120 153904
rect 131172 153932 131178 153944
rect 223666 153932 223672 153944
rect 131172 153904 223672 153932
rect 131172 153892 131178 153904
rect 223666 153892 223672 153904
rect 223724 153892 223730 153944
rect 65978 153824 65984 153876
rect 66036 153864 66042 153876
rect 158714 153864 158720 153876
rect 66036 153836 158720 153864
rect 66036 153824 66042 153836
rect 158714 153824 158720 153836
rect 158772 153824 158778 153876
rect 192478 153824 192484 153876
rect 192536 153864 192542 153876
rect 218054 153864 218060 153876
rect 192536 153836 218060 153864
rect 192536 153824 192542 153836
rect 218054 153824 218060 153836
rect 218112 153824 218118 153876
rect 187510 153212 187516 153264
rect 187568 153252 187574 153264
rect 191834 153252 191840 153264
rect 187568 153224 191840 153252
rect 187568 153212 187574 153224
rect 191834 153212 191840 153224
rect 191892 153212 191898 153264
rect 222378 152464 222384 152516
rect 222436 152504 222442 152516
rect 222838 152504 222844 152516
rect 222436 152476 222844 152504
rect 222436 152464 222442 152476
rect 222838 152464 222844 152476
rect 222896 152464 222902 152516
rect 182910 151920 182916 151972
rect 182968 151960 182974 151972
rect 222838 151960 222844 151972
rect 182968 151932 222844 151960
rect 182968 151920 182974 151932
rect 222838 151920 222844 151932
rect 222896 151920 222902 151972
rect 62022 151852 62028 151904
rect 62080 151892 62086 151904
rect 131850 151892 131856 151904
rect 62080 151864 131856 151892
rect 62080 151852 62086 151864
rect 131850 151852 131856 151864
rect 131908 151852 131914 151904
rect 151262 151852 151268 151904
rect 151320 151892 151326 151904
rect 208486 151892 208492 151904
rect 151320 151864 208492 151892
rect 151320 151852 151326 151864
rect 208486 151852 208492 151864
rect 208544 151852 208550 151904
rect 69750 151784 69756 151836
rect 69808 151824 69814 151836
rect 160186 151824 160192 151836
rect 69808 151796 160192 151824
rect 69808 151784 69814 151796
rect 160186 151784 160192 151796
rect 160244 151824 160250 151836
rect 160738 151824 160744 151836
rect 160244 151796 160744 151824
rect 160244 151784 160250 151796
rect 160738 151784 160744 151796
rect 160796 151784 160802 151836
rect 220814 151784 220820 151836
rect 220872 151824 220878 151836
rect 222102 151824 222108 151836
rect 220872 151796 222108 151824
rect 220872 151784 220878 151796
rect 222102 151784 222108 151796
rect 222160 151824 222166 151836
rect 302234 151824 302240 151836
rect 222160 151796 302240 151824
rect 222160 151784 222166 151796
rect 302234 151784 302240 151796
rect 302292 151784 302298 151836
rect 74810 151104 74816 151156
rect 74868 151144 74874 151156
rect 177942 151144 177948 151156
rect 74868 151116 177948 151144
rect 74868 151104 74874 151116
rect 177942 151104 177948 151116
rect 178000 151144 178006 151156
rect 178000 151116 180794 151144
rect 178000 151104 178006 151116
rect 63402 151036 63408 151088
rect 63460 151076 63466 151088
rect 167638 151076 167644 151088
rect 63460 151048 167644 151076
rect 63460 151036 63466 151048
rect 167638 151036 167644 151048
rect 167696 151036 167702 151088
rect 180766 151076 180794 151116
rect 189626 151104 189632 151156
rect 189684 151144 189690 151156
rect 201494 151144 201500 151156
rect 189684 151116 201500 151144
rect 189684 151104 189690 151116
rect 201494 151104 201500 151116
rect 201552 151104 201558 151156
rect 201586 151076 201592 151088
rect 180766 151048 201592 151076
rect 201586 151036 201592 151048
rect 201644 151036 201650 151088
rect 207842 151036 207848 151088
rect 207900 151076 207906 151088
rect 220814 151076 220820 151088
rect 207900 151048 220820 151076
rect 207900 151036 207906 151048
rect 220814 151036 220820 151048
rect 220872 151036 220878 151088
rect 204162 150424 204168 150476
rect 204220 150464 204226 150476
rect 230658 150464 230664 150476
rect 204220 150436 230664 150464
rect 204220 150424 204226 150436
rect 230658 150424 230664 150436
rect 230716 150424 230722 150476
rect 148594 149744 148600 149796
rect 148652 149784 148658 149796
rect 204162 149784 204168 149796
rect 148652 149756 204168 149784
rect 148652 149744 148658 149756
rect 204162 149744 204168 149756
rect 204220 149744 204226 149796
rect 206370 149744 206376 149796
rect 206428 149784 206434 149796
rect 252462 149784 252468 149796
rect 206428 149756 252468 149784
rect 206428 149744 206434 149756
rect 252462 149744 252468 149756
rect 252520 149744 252526 149796
rect 86862 149676 86868 149728
rect 86920 149716 86926 149728
rect 124858 149716 124864 149728
rect 86920 149688 124864 149716
rect 86920 149676 86926 149688
rect 124858 149676 124864 149688
rect 124916 149716 124922 149728
rect 216766 149716 216772 149728
rect 124916 149688 216772 149716
rect 124916 149676 124922 149688
rect 216766 149676 216772 149688
rect 216824 149676 216830 149728
rect 252462 149132 252468 149184
rect 252520 149172 252526 149184
rect 256050 149172 256056 149184
rect 252520 149144 256056 149172
rect 252520 149132 252526 149144
rect 256050 149132 256056 149144
rect 256108 149132 256114 149184
rect 67542 149064 67548 149116
rect 67600 149104 67606 149116
rect 111150 149104 111156 149116
rect 67600 149076 111156 149104
rect 67600 149064 67606 149076
rect 111150 149064 111156 149076
rect 111208 149064 111214 149116
rect 216858 149064 216864 149116
rect 216916 149104 216922 149116
rect 217318 149104 217324 149116
rect 216916 149076 217324 149104
rect 216916 149064 216922 149076
rect 217318 149064 217324 149076
rect 217376 149104 217382 149116
rect 582742 149104 582748 149116
rect 217376 149076 582748 149104
rect 217376 149064 217382 149076
rect 582742 149064 582748 149076
rect 582800 149064 582806 149116
rect 193030 148996 193036 149048
rect 193088 149036 193094 149048
rect 211062 149036 211068 149048
rect 193088 149008 211068 149036
rect 193088 148996 193094 149008
rect 211062 148996 211068 149008
rect 211120 148996 211126 149048
rect 218514 148996 218520 149048
rect 218572 149036 218578 149048
rect 218698 149036 218704 149048
rect 218572 149008 218704 149036
rect 218572 148996 218578 149008
rect 218698 148996 218704 149008
rect 218756 149036 218762 149048
rect 267826 149036 267832 149048
rect 218756 149008 267832 149036
rect 218756 148996 218762 149008
rect 267826 148996 267832 149008
rect 267884 148996 267890 149048
rect 190362 148384 190368 148436
rect 190420 148424 190426 148436
rect 193214 148424 193220 148436
rect 190420 148396 193220 148424
rect 190420 148384 190426 148396
rect 193214 148384 193220 148396
rect 193272 148384 193278 148436
rect 64690 148316 64696 148368
rect 64748 148356 64754 148368
rect 192478 148356 192484 148368
rect 64748 148328 192484 148356
rect 64748 148316 64754 148328
rect 192478 148316 192484 148328
rect 192536 148316 192542 148368
rect 48222 147636 48228 147688
rect 48280 147676 48286 147688
rect 104158 147676 104164 147688
rect 48280 147648 104164 147676
rect 48280 147636 48286 147648
rect 104158 147636 104164 147648
rect 104216 147636 104222 147688
rect 212994 147636 213000 147688
rect 213052 147676 213058 147688
rect 233878 147676 233884 147688
rect 213052 147648 233884 147676
rect 213052 147636 213058 147648
rect 233878 147636 233884 147648
rect 233936 147636 233942 147688
rect 214006 147568 214012 147620
rect 214064 147608 214070 147620
rect 216858 147608 216864 147620
rect 214064 147580 216864 147608
rect 214064 147568 214070 147580
rect 216858 147568 216864 147580
rect 216916 147568 216922 147620
rect 208394 146956 208400 147008
rect 208452 146996 208458 147008
rect 209130 146996 209136 147008
rect 208452 146968 209136 146996
rect 208452 146956 208458 146968
rect 209130 146956 209136 146968
rect 209188 146956 209194 147008
rect 3142 146888 3148 146940
rect 3200 146928 3206 146940
rect 95418 146928 95424 146940
rect 3200 146900 95424 146928
rect 3200 146888 3206 146900
rect 95418 146888 95424 146900
rect 95476 146928 95482 146940
rect 153930 146928 153936 146940
rect 95476 146900 153936 146928
rect 95476 146888 95482 146900
rect 153930 146888 153936 146900
rect 153988 146888 153994 146940
rect 154022 146888 154028 146940
rect 154080 146928 154086 146940
rect 187694 146928 187700 146940
rect 154080 146900 187700 146928
rect 154080 146888 154086 146900
rect 187694 146888 187700 146900
rect 187752 146888 187758 146940
rect 252186 146888 252192 146940
rect 252244 146928 252250 146940
rect 288710 146928 288716 146940
rect 252244 146900 288716 146928
rect 252244 146888 252250 146900
rect 288710 146888 288716 146900
rect 288768 146928 288774 146940
rect 327074 146928 327080 146940
rect 288768 146900 327080 146928
rect 288768 146888 288774 146900
rect 327074 146888 327080 146900
rect 327132 146888 327138 146940
rect 221458 146344 221464 146396
rect 221516 146384 221522 146396
rect 256142 146384 256148 146396
rect 221516 146356 256148 146384
rect 221516 146344 221522 146356
rect 256142 146344 256148 146356
rect 256200 146344 256206 146396
rect 67266 146276 67272 146328
rect 67324 146316 67330 146328
rect 97442 146316 97448 146328
rect 67324 146288 97448 146316
rect 67324 146276 67330 146288
rect 97442 146276 97448 146288
rect 97500 146276 97506 146328
rect 100018 146276 100024 146328
rect 100076 146316 100082 146328
rect 100570 146316 100576 146328
rect 100076 146288 100576 146316
rect 100076 146276 100082 146288
rect 100570 146276 100576 146288
rect 100628 146316 100634 146328
rect 224954 146316 224960 146328
rect 100628 146288 224960 146316
rect 100628 146276 100634 146288
rect 224954 146276 224960 146288
rect 225012 146276 225018 146328
rect 4798 146208 4804 146260
rect 4856 146248 4862 146260
rect 86862 146248 86868 146260
rect 4856 146220 86868 146248
rect 4856 146208 4862 146220
rect 86862 146208 86868 146220
rect 86920 146248 86926 146260
rect 87598 146248 87604 146260
rect 86920 146220 87604 146248
rect 86920 146208 86926 146220
rect 87598 146208 87604 146220
rect 87656 146208 87662 146260
rect 89622 146208 89628 146260
rect 89680 146248 89686 146260
rect 95234 146248 95240 146260
rect 89680 146220 95240 146248
rect 89680 146208 89686 146220
rect 95234 146208 95240 146220
rect 95292 146208 95298 146260
rect 218790 146208 218796 146260
rect 218848 146248 218854 146260
rect 221090 146248 221096 146260
rect 218848 146220 221096 146248
rect 218848 146208 218854 146220
rect 221090 146208 221096 146220
rect 221148 146208 221154 146260
rect 204898 145528 204904 145580
rect 204956 145568 204962 145580
rect 234706 145568 234712 145580
rect 204956 145540 234712 145568
rect 204956 145528 204962 145540
rect 234706 145528 234712 145540
rect 234764 145528 234770 145580
rect 259362 145528 259368 145580
rect 259420 145568 259426 145580
rect 277578 145568 277584 145580
rect 259420 145540 277584 145568
rect 259420 145528 259426 145540
rect 277578 145528 277584 145540
rect 277636 145528 277642 145580
rect 177850 144984 177856 145036
rect 177908 145024 177914 145036
rect 209866 145024 209872 145036
rect 177908 144996 209872 145024
rect 177908 144984 177914 144996
rect 209866 144984 209872 144996
rect 209924 144984 209930 145036
rect 71774 144916 71780 144968
rect 71832 144956 71838 144968
rect 72878 144956 72884 144968
rect 71832 144928 72884 144956
rect 71832 144916 71838 144928
rect 72878 144916 72884 144928
rect 72936 144956 72942 144968
rect 198366 144956 198372 144968
rect 72936 144928 198372 144956
rect 72936 144916 72942 144928
rect 198366 144916 198372 144928
rect 198424 144916 198430 144968
rect 228358 144916 228364 144968
rect 228416 144956 228422 144968
rect 349798 144956 349804 144968
rect 228416 144928 349804 144956
rect 228416 144916 228422 144928
rect 349798 144916 349804 144928
rect 349856 144916 349862 144968
rect 85574 144712 85580 144764
rect 85632 144752 85638 144764
rect 88978 144752 88984 144764
rect 85632 144724 88984 144752
rect 85632 144712 85638 144724
rect 88978 144712 88984 144724
rect 89036 144712 89042 144764
rect 90082 144712 90088 144764
rect 90140 144752 90146 144764
rect 93118 144752 93124 144764
rect 90140 144724 93124 144752
rect 90140 144712 90146 144724
rect 93118 144712 93124 144724
rect 93176 144712 93182 144764
rect 186958 144372 186964 144424
rect 187016 144412 187022 144424
rect 193582 144412 193588 144424
rect 187016 144384 193588 144412
rect 187016 144372 187022 144384
rect 193582 144372 193588 144384
rect 193640 144372 193646 144424
rect 175918 144236 175924 144288
rect 175976 144276 175982 144288
rect 194134 144276 194140 144288
rect 175976 144248 194140 144276
rect 175976 144236 175982 144248
rect 194134 144236 194140 144248
rect 194192 144236 194198 144288
rect 102134 144168 102140 144220
rect 102192 144208 102198 144220
rect 178770 144208 178776 144220
rect 102192 144180 178776 144208
rect 102192 144168 102198 144180
rect 178770 144168 178776 144180
rect 178828 144168 178834 144220
rect 224494 144168 224500 144220
rect 224552 144208 224558 144220
rect 224862 144208 224868 144220
rect 224552 144180 224868 144208
rect 224552 144168 224558 144180
rect 224862 144168 224868 144180
rect 224920 144208 224926 144220
rect 238110 144208 238116 144220
rect 224920 144180 238116 144208
rect 224920 144168 224926 144180
rect 238110 144168 238116 144180
rect 238168 144168 238174 144220
rect 249058 144168 249064 144220
rect 249116 144208 249122 144220
rect 262214 144208 262220 144220
rect 249116 144180 262220 144208
rect 249116 144168 249122 144180
rect 262214 144168 262220 144180
rect 262272 144168 262278 144220
rect 223666 144032 223672 144084
rect 223724 144072 223730 144084
rect 224494 144072 224500 144084
rect 223724 144044 224500 144072
rect 223724 144032 223730 144044
rect 224494 144032 224500 144044
rect 224552 144032 224558 144084
rect 200114 143964 200120 144016
rect 200172 144004 200178 144016
rect 200390 144004 200396 144016
rect 200172 143976 200396 144004
rect 200172 143964 200178 143976
rect 200390 143964 200396 143976
rect 200448 143964 200454 144016
rect 204254 143964 204260 144016
rect 204312 144004 204318 144016
rect 204622 144004 204628 144016
rect 204312 143976 204628 144004
rect 204312 143964 204318 143976
rect 204622 143964 204628 143976
rect 204680 143964 204686 144016
rect 59262 143556 59268 143608
rect 59320 143596 59326 143608
rect 167730 143596 167736 143608
rect 59320 143568 167736 143596
rect 59320 143556 59326 143568
rect 167730 143556 167736 143568
rect 167788 143556 167794 143608
rect 245010 143596 245016 143608
rect 198660 143568 245016 143596
rect 195422 143488 195428 143540
rect 195480 143528 195486 143540
rect 197906 143528 197912 143540
rect 195480 143500 197912 143528
rect 195480 143488 195486 143500
rect 197906 143488 197912 143500
rect 197964 143528 197970 143540
rect 198660 143528 198688 143568
rect 245010 143556 245016 143568
rect 245068 143556 245074 143608
rect 197964 143500 198688 143528
rect 197964 143488 197970 143500
rect 219526 143488 219532 143540
rect 219584 143528 219590 143540
rect 220170 143528 220176 143540
rect 219584 143500 220176 143528
rect 219584 143488 219590 143500
rect 220170 143488 220176 143500
rect 220228 143488 220234 143540
rect 259362 143488 259368 143540
rect 259420 143528 259426 143540
rect 260098 143528 260104 143540
rect 259420 143500 260104 143528
rect 259420 143488 259426 143500
rect 260098 143488 260104 143500
rect 260156 143488 260162 143540
rect 199010 142916 199016 142928
rect 195946 142888 199016 142916
rect 60642 142808 60648 142860
rect 60700 142848 60706 142860
rect 77938 142848 77944 142860
rect 60700 142820 77944 142848
rect 60700 142808 60706 142820
rect 77938 142808 77944 142820
rect 77996 142808 78002 142860
rect 120718 142808 120724 142860
rect 120776 142848 120782 142860
rect 195946 142848 195974 142888
rect 199010 142876 199016 142888
rect 199068 142916 199074 142928
rect 218238 142916 218244 142928
rect 199068 142888 218244 142916
rect 199068 142876 199074 142888
rect 218238 142876 218244 142888
rect 218296 142876 218302 142928
rect 120776 142820 195974 142848
rect 120776 142808 120782 142820
rect 212902 142808 212908 142860
rect 212960 142848 212966 142860
rect 259362 142848 259368 142860
rect 212960 142820 259368 142848
rect 212960 142808 212966 142820
rect 259362 142808 259368 142820
rect 259420 142808 259426 142860
rect 63126 142128 63132 142180
rect 63184 142168 63190 142180
rect 88518 142168 88524 142180
rect 63184 142140 88524 142168
rect 63184 142128 63190 142140
rect 88518 142128 88524 142140
rect 88576 142128 88582 142180
rect 220078 142128 220084 142180
rect 220136 142168 220142 142180
rect 225690 142168 225696 142180
rect 220136 142140 225696 142168
rect 220136 142128 220142 142140
rect 225690 142128 225696 142140
rect 225748 142128 225754 142180
rect 69842 142060 69848 142112
rect 69900 142100 69906 142112
rect 76006 142100 76012 142112
rect 69900 142072 76012 142100
rect 69900 142060 69906 142072
rect 76006 142060 76012 142072
rect 76064 142060 76070 142112
rect 76006 141380 76012 141432
rect 76064 141420 76070 141432
rect 159450 141420 159456 141432
rect 76064 141392 159456 141420
rect 76064 141380 76070 141392
rect 159450 141380 159456 141392
rect 159508 141420 159514 141432
rect 203150 141420 203156 141432
rect 159508 141392 203156 141420
rect 159508 141380 159514 141392
rect 203150 141380 203156 141392
rect 203208 141380 203214 141432
rect 69106 140836 69112 140888
rect 69164 140876 69170 140888
rect 69842 140876 69848 140888
rect 69164 140848 69848 140876
rect 69164 140836 69170 140848
rect 69842 140836 69848 140848
rect 69900 140836 69906 140888
rect 205634 140836 205640 140888
rect 205692 140876 205698 140888
rect 266354 140876 266360 140888
rect 205692 140848 266360 140876
rect 205692 140836 205698 140848
rect 266354 140836 266360 140848
rect 266412 140876 266418 140888
rect 266998 140876 267004 140888
rect 266412 140848 267004 140876
rect 266412 140836 266418 140848
rect 266998 140836 267004 140848
rect 267056 140836 267062 140888
rect 57790 140768 57796 140820
rect 57848 140808 57854 140820
rect 91094 140808 91100 140820
rect 57848 140780 91100 140808
rect 57848 140768 57854 140780
rect 91094 140768 91100 140780
rect 91152 140768 91158 140820
rect 203426 140768 203432 140820
rect 203484 140808 203490 140820
rect 289078 140808 289084 140820
rect 203484 140780 289084 140808
rect 203484 140768 203490 140780
rect 289078 140768 289084 140780
rect 289136 140768 289142 140820
rect 210142 140604 210148 140616
rect 195946 140576 210148 140604
rect 193030 140496 193036 140548
rect 193088 140536 193094 140548
rect 194870 140536 194876 140548
rect 193088 140508 194876 140536
rect 193088 140496 193094 140508
rect 194870 140496 194876 140508
rect 194928 140496 194934 140548
rect 89070 140088 89076 140140
rect 89128 140128 89134 140140
rect 120718 140128 120724 140140
rect 89128 140100 120724 140128
rect 89128 140088 89134 140100
rect 120718 140088 120724 140100
rect 120776 140088 120782 140140
rect 193398 140088 193404 140140
rect 193456 140128 193462 140140
rect 195946 140128 195974 140576
rect 210142 140564 210148 140576
rect 210200 140564 210206 140616
rect 193456 140100 195974 140128
rect 200776 140508 209774 140536
rect 193456 140088 193462 140100
rect 68646 140020 68652 140072
rect 68704 140060 68710 140072
rect 80698 140060 80704 140072
rect 68704 140032 80704 140060
rect 68704 140020 68710 140032
rect 80698 140020 80704 140032
rect 80756 140020 80762 140072
rect 84470 140020 84476 140072
rect 84528 140060 84534 140072
rect 118878 140060 118884 140072
rect 84528 140032 118884 140060
rect 84528 140020 84534 140032
rect 118878 140020 118884 140032
rect 118936 140020 118942 140072
rect 173250 140020 173256 140072
rect 173308 140060 173314 140072
rect 184474 140060 184480 140072
rect 173308 140032 184480 140060
rect 173308 140020 173314 140032
rect 184474 140020 184480 140032
rect 184532 140020 184538 140072
rect 71314 139408 71320 139460
rect 71372 139448 71378 139460
rect 73798 139448 73804 139460
rect 71372 139420 73804 139448
rect 71372 139408 71378 139420
rect 73798 139408 73804 139420
rect 73856 139408 73862 139460
rect 118878 139408 118884 139460
rect 118936 139448 118942 139460
rect 200776 139448 200804 140508
rect 205174 140428 205180 140480
rect 205232 140428 205238 140480
rect 209746 140468 209774 140508
rect 210050 140496 210056 140548
rect 210108 140536 210114 140548
rect 210108 140508 213040 140536
rect 210108 140496 210114 140508
rect 212534 140468 212540 140480
rect 209746 140440 212540 140468
rect 212534 140428 212540 140440
rect 212592 140428 212598 140480
rect 118936 139420 200804 139448
rect 118936 139408 118942 139420
rect 79410 139340 79416 139392
rect 79468 139380 79474 139392
rect 205192 139380 205220 140428
rect 213012 140400 213040 140508
rect 215386 140428 215392 140480
rect 215444 140468 215450 140480
rect 225138 140468 225144 140480
rect 215444 140440 225144 140468
rect 215444 140428 215450 140440
rect 225138 140428 225144 140440
rect 225196 140428 225202 140480
rect 213012 140372 219434 140400
rect 219406 140060 219434 140372
rect 287698 140060 287704 140072
rect 219406 140032 287704 140060
rect 287698 140020 287704 140032
rect 287756 140020 287762 140072
rect 225138 139408 225144 139460
rect 225196 139448 225202 139460
rect 249702 139448 249708 139460
rect 225196 139420 249708 139448
rect 225196 139408 225202 139420
rect 249702 139408 249708 139420
rect 249760 139448 249766 139460
rect 251174 139448 251180 139460
rect 249760 139420 251180 139448
rect 249760 139408 249766 139420
rect 251174 139408 251180 139420
rect 251232 139408 251238 139460
rect 79468 139352 205220 139380
rect 79468 139340 79474 139352
rect 226702 139204 226708 139256
rect 226760 139244 226766 139256
rect 229186 139244 229192 139256
rect 226760 139216 229192 139244
rect 226760 139204 226766 139216
rect 229186 139204 229192 139216
rect 229244 139204 229250 139256
rect 66162 138660 66168 138712
rect 66220 138700 66226 138712
rect 178678 138700 178684 138712
rect 66220 138672 178684 138700
rect 66220 138660 66226 138672
rect 178678 138660 178684 138672
rect 178736 138660 178742 138712
rect 235994 138660 236000 138712
rect 236052 138700 236058 138712
rect 582650 138700 582656 138712
rect 236052 138672 582656 138700
rect 236052 138660 236058 138672
rect 582650 138660 582656 138672
rect 582708 138660 582714 138712
rect 93854 138048 93860 138100
rect 93912 138088 93918 138100
rect 94314 138088 94320 138100
rect 93912 138060 94320 138088
rect 93912 138048 93918 138060
rect 94314 138048 94320 138060
rect 94372 138048 94378 138100
rect 65886 137980 65892 138032
rect 65944 138020 65950 138032
rect 66162 138020 66168 138032
rect 65944 137992 66168 138020
rect 65944 137980 65950 137992
rect 66162 137980 66168 137992
rect 66220 137980 66226 138032
rect 2866 137912 2872 137964
rect 2924 137952 2930 137964
rect 72970 137952 72976 137964
rect 2924 137924 72976 137952
rect 2924 137912 2930 137924
rect 72970 137912 72976 137924
rect 73028 137952 73034 137964
rect 73154 137952 73160 137964
rect 73028 137924 73160 137952
rect 73028 137912 73034 137924
rect 73154 137912 73160 137924
rect 73212 137912 73218 137964
rect 78490 137912 78496 137964
rect 78548 137952 78554 137964
rect 79410 137952 79416 137964
rect 78548 137924 79416 137952
rect 78548 137912 78554 137924
rect 79410 137912 79416 137924
rect 79468 137912 79474 137964
rect 87046 137912 87052 137964
rect 87104 137952 87110 137964
rect 193214 137952 193220 137964
rect 87104 137924 193220 137952
rect 87104 137912 87110 137924
rect 193214 137912 193220 137924
rect 193272 137912 193278 137964
rect 226702 137912 226708 137964
rect 226760 137952 226766 137964
rect 234614 137952 234620 137964
rect 226760 137924 234620 137952
rect 226760 137912 226766 137924
rect 234614 137912 234620 137924
rect 234672 137952 234678 137964
rect 240870 137952 240876 137964
rect 234672 137924 240876 137952
rect 234672 137912 234678 137924
rect 240870 137912 240876 137924
rect 240928 137912 240934 137964
rect 58894 137232 58900 137284
rect 58952 137272 58958 137284
rect 69198 137272 69204 137284
rect 58952 137244 69204 137272
rect 58952 137232 58958 137244
rect 69198 137232 69204 137244
rect 69256 137232 69262 137284
rect 91094 137232 91100 137284
rect 91152 137272 91158 137284
rect 151354 137272 151360 137284
rect 91152 137244 151360 137272
rect 91152 137232 91158 137244
rect 151354 137232 151360 137244
rect 151412 137232 151418 137284
rect 247678 137232 247684 137284
rect 247736 137272 247742 137284
rect 255314 137272 255320 137284
rect 247736 137244 255320 137272
rect 247736 137232 247742 137244
rect 255314 137232 255320 137244
rect 255372 137232 255378 137284
rect 256142 137232 256148 137284
rect 256200 137272 256206 137284
rect 276014 137272 276020 137284
rect 256200 137244 276020 137272
rect 256200 137232 256206 137244
rect 276014 137232 276020 137244
rect 276072 137232 276078 137284
rect 91002 136824 91008 136876
rect 91060 136864 91066 136876
rect 91830 136864 91836 136876
rect 91060 136836 91836 136864
rect 91060 136824 91066 136836
rect 91830 136824 91836 136836
rect 91888 136824 91894 136876
rect 87046 136728 87052 136740
rect 80026 136700 87052 136728
rect 79594 136620 79600 136672
rect 79652 136660 79658 136672
rect 80026 136660 80054 136700
rect 87046 136688 87052 136700
rect 87104 136688 87110 136740
rect 79652 136632 80054 136660
rect 79652 136620 79658 136632
rect 81342 136620 81348 136672
rect 81400 136660 81406 136672
rect 82170 136660 82176 136672
rect 81400 136632 82176 136660
rect 81400 136620 81406 136632
rect 82170 136620 82176 136632
rect 82228 136620 82234 136672
rect 85482 136620 85488 136672
rect 85540 136660 85546 136672
rect 86218 136660 86224 136672
rect 85540 136632 86224 136660
rect 85540 136620 85546 136632
rect 86218 136620 86224 136632
rect 86276 136620 86282 136672
rect 91186 136552 91192 136604
rect 91244 136592 91250 136604
rect 91738 136592 91744 136604
rect 91244 136564 91744 136592
rect 91244 136552 91250 136564
rect 91738 136552 91744 136564
rect 91796 136552 91802 136604
rect 170398 136552 170404 136604
rect 170456 136592 170462 136604
rect 191558 136592 191564 136604
rect 170456 136564 191564 136592
rect 170456 136552 170462 136564
rect 191558 136552 191564 136564
rect 191616 136552 191622 136604
rect 159450 135940 159456 135992
rect 159508 135980 159514 135992
rect 169018 135980 169024 135992
rect 159508 135952 169024 135980
rect 159508 135940 159514 135952
rect 169018 135940 169024 135952
rect 169076 135940 169082 135992
rect 160186 135872 160192 135924
rect 160244 135912 160250 135924
rect 161382 135912 161388 135924
rect 160244 135884 161388 135912
rect 160244 135872 160250 135884
rect 161382 135872 161388 135884
rect 161440 135912 161446 135924
rect 175918 135912 175924 135924
rect 161440 135884 175924 135912
rect 161440 135872 161446 135884
rect 175918 135872 175924 135884
rect 175976 135872 175982 135924
rect 256050 135872 256056 135924
rect 256108 135912 256114 135924
rect 298738 135912 298744 135924
rect 256108 135884 298744 135912
rect 256108 135872 256114 135884
rect 298738 135872 298744 135884
rect 298796 135872 298802 135924
rect 53098 135328 53104 135380
rect 53156 135368 53162 135380
rect 91278 135368 91284 135380
rect 53156 135340 91284 135368
rect 53156 135328 53162 135340
rect 91278 135328 91284 135340
rect 91336 135328 91342 135380
rect 4798 135260 4804 135312
rect 4856 135300 4862 135312
rect 91186 135300 91192 135312
rect 4856 135272 91192 135300
rect 4856 135260 4862 135272
rect 91186 135260 91192 135272
rect 91244 135260 91250 135312
rect 187694 135260 187700 135312
rect 187752 135300 187758 135312
rect 191558 135300 191564 135312
rect 187752 135272 191564 135300
rect 187752 135260 187758 135272
rect 191558 135260 191564 135272
rect 191616 135260 191622 135312
rect 97902 135192 97908 135244
rect 97960 135232 97966 135244
rect 137462 135232 137468 135244
rect 97960 135204 137468 135232
rect 97960 135192 97966 135204
rect 137462 135192 137468 135204
rect 137520 135192 137526 135244
rect 226702 135192 226708 135244
rect 226760 135232 226766 135244
rect 231946 135232 231952 135244
rect 226760 135204 231952 135232
rect 226760 135192 226766 135204
rect 231946 135192 231952 135204
rect 232004 135192 232010 135244
rect 188430 134852 188436 134904
rect 188488 134892 188494 134904
rect 191190 134892 191196 134904
rect 188488 134864 191196 134892
rect 188488 134852 188494 134864
rect 191190 134852 191196 134864
rect 191248 134852 191254 134904
rect 70302 134784 70308 134836
rect 70360 134824 70366 134836
rect 75362 134824 75368 134836
rect 70360 134796 75368 134824
rect 70360 134784 70366 134796
rect 75362 134784 75368 134796
rect 75420 134784 75426 134836
rect 68554 134580 68560 134632
rect 68612 134620 68618 134632
rect 69750 134620 69756 134632
rect 68612 134592 69756 134620
rect 68612 134580 68618 134592
rect 69750 134580 69756 134592
rect 69808 134580 69814 134632
rect 93762 134580 93768 134632
rect 93820 134620 93826 134632
rect 93820 134580 93854 134620
rect 93826 134552 93854 134580
rect 189166 134552 189172 134564
rect 93826 134524 189172 134552
rect 189166 134512 189172 134524
rect 189224 134512 189230 134564
rect 226610 134512 226616 134564
rect 226668 134552 226674 134564
rect 309778 134552 309784 134564
rect 226668 134524 309784 134552
rect 226668 134512 226674 134524
rect 309778 134512 309784 134524
rect 309836 134512 309842 134564
rect 95142 133832 95148 133884
rect 95200 133872 95206 133884
rect 177574 133872 177580 133884
rect 95200 133844 177580 133872
rect 95200 133832 95206 133844
rect 177574 133832 177580 133844
rect 177632 133832 177638 133884
rect 226610 133832 226616 133884
rect 226668 133872 226674 133884
rect 237374 133872 237380 133884
rect 226668 133844 237380 133872
rect 226668 133832 226674 133844
rect 237374 133832 237380 133844
rect 237432 133832 237438 133884
rect 226702 133628 226708 133680
rect 226760 133668 226766 133680
rect 231118 133668 231124 133680
rect 226760 133640 231124 133668
rect 226760 133628 226766 133640
rect 231118 133628 231124 133640
rect 231176 133628 231182 133680
rect 148502 133220 148508 133272
rect 148560 133260 148566 133272
rect 187694 133260 187700 133272
rect 148560 133232 187700 133260
rect 148560 133220 148566 133232
rect 187694 133220 187700 133232
rect 187752 133220 187758 133272
rect 103698 133152 103704 133204
rect 103756 133192 103762 133204
rect 148594 133192 148600 133204
rect 103756 133164 148600 133192
rect 103756 133152 103762 133164
rect 148594 133152 148600 133164
rect 148652 133152 148658 133204
rect 52178 132404 52184 132456
rect 52236 132444 52242 132456
rect 66898 132444 66904 132456
rect 52236 132416 66904 132444
rect 52236 132404 52242 132416
rect 66898 132404 66904 132416
rect 66956 132404 66962 132456
rect 97902 132404 97908 132456
rect 97960 132444 97966 132456
rect 142982 132444 142988 132456
rect 97960 132416 142988 132444
rect 97960 132404 97966 132416
rect 142982 132404 142988 132416
rect 143040 132404 143046 132456
rect 226702 132404 226708 132456
rect 226760 132444 226766 132456
rect 249886 132444 249892 132456
rect 226760 132416 249892 132444
rect 226760 132404 226766 132416
rect 249886 132404 249892 132416
rect 249944 132404 249950 132456
rect 56318 132336 56324 132388
rect 56376 132376 56382 132388
rect 66806 132376 66812 132388
rect 56376 132348 66812 132376
rect 56376 132336 56382 132348
rect 66806 132336 66812 132348
rect 66864 132336 66870 132388
rect 180150 131792 180156 131844
rect 180208 131832 180214 131844
rect 190454 131832 190460 131844
rect 180208 131804 190460 131832
rect 180208 131792 180214 131804
rect 190454 131792 190460 131804
rect 190512 131792 190518 131844
rect 150434 131724 150440 131776
rect 150492 131764 150498 131776
rect 182910 131764 182916 131776
rect 150492 131736 182916 131764
rect 150492 131724 150498 131736
rect 182910 131724 182916 131736
rect 182968 131724 182974 131776
rect 240778 131724 240784 131776
rect 240836 131764 240842 131776
rect 335446 131764 335452 131776
rect 240836 131736 335452 131764
rect 240836 131724 240842 131736
rect 335446 131724 335452 131736
rect 335504 131724 335510 131776
rect 104894 131112 104900 131164
rect 104952 131152 104958 131164
rect 111058 131152 111064 131164
rect 104952 131124 111064 131152
rect 104952 131112 104958 131124
rect 111058 131112 111064 131124
rect 111116 131112 111122 131164
rect 63126 131044 63132 131096
rect 63184 131084 63190 131096
rect 66806 131084 66812 131096
rect 63184 131056 66812 131084
rect 63184 131044 63190 131056
rect 66806 131044 66812 131056
rect 66864 131044 66870 131096
rect 169202 131044 169208 131096
rect 169260 131084 169266 131096
rect 189810 131084 189816 131096
rect 169260 131056 189816 131084
rect 169260 131044 169266 131056
rect 189810 131044 189816 131056
rect 189868 131044 189874 131096
rect 226702 131044 226708 131096
rect 226760 131084 226766 131096
rect 230658 131084 230664 131096
rect 226760 131056 230664 131084
rect 226760 131044 226766 131056
rect 230658 131044 230664 131056
rect 230716 131084 230722 131096
rect 276106 131084 276112 131096
rect 230716 131056 276112 131084
rect 230716 131044 230722 131056
rect 276106 131044 276112 131056
rect 276164 131044 276170 131096
rect 226794 130976 226800 131028
rect 226852 131016 226858 131028
rect 233234 131016 233240 131028
rect 226852 130988 233240 131016
rect 226852 130976 226858 130988
rect 233234 130976 233240 130988
rect 233292 131016 233298 131028
rect 267734 131016 267740 131028
rect 233292 130988 267740 131016
rect 233292 130976 233298 130988
rect 267734 130976 267740 130988
rect 267792 130976 267798 131028
rect 97534 130568 97540 130620
rect 97592 130608 97598 130620
rect 102870 130608 102876 130620
rect 97592 130580 102876 130608
rect 97592 130568 97598 130580
rect 102870 130568 102876 130580
rect 102928 130568 102934 130620
rect 97718 130364 97724 130416
rect 97776 130404 97782 130416
rect 181530 130404 181536 130416
rect 97776 130376 181536 130404
rect 97776 130364 97782 130376
rect 181530 130364 181536 130376
rect 181588 130364 181594 130416
rect 97902 129684 97908 129736
rect 97960 129724 97966 129736
rect 106366 129724 106372 129736
rect 97960 129696 106372 129724
rect 97960 129684 97966 129696
rect 106366 129684 106372 129696
rect 106424 129684 106430 129736
rect 151354 129684 151360 129736
rect 151412 129724 151418 129736
rect 191742 129724 191748 129736
rect 151412 129696 191748 129724
rect 151412 129684 151418 129696
rect 191742 129684 191748 129696
rect 191800 129684 191806 129736
rect 114554 129072 114560 129124
rect 114612 129112 114618 129124
rect 148410 129112 148416 129124
rect 114612 129084 148416 129112
rect 114612 129072 114618 129084
rect 148410 129072 148416 129084
rect 148468 129072 148474 129124
rect 97442 129004 97448 129056
rect 97500 129044 97506 129056
rect 160830 129044 160836 129056
rect 97500 129016 160836 129044
rect 97500 129004 97506 129016
rect 160830 129004 160836 129016
rect 160888 129004 160894 129056
rect 61746 128324 61752 128376
rect 61804 128364 61810 128376
rect 66806 128364 66812 128376
rect 61804 128336 66812 128364
rect 61804 128324 61810 128336
rect 66806 128324 66812 128336
rect 66864 128324 66870 128376
rect 226426 128324 226432 128376
rect 226484 128364 226490 128376
rect 299474 128364 299480 128376
rect 226484 128336 299480 128364
rect 226484 128324 226490 128336
rect 299474 128324 299480 128336
rect 299532 128324 299538 128376
rect 97626 128256 97632 128308
rect 97684 128296 97690 128308
rect 140130 128296 140136 128308
rect 97684 128268 140136 128296
rect 97684 128256 97690 128268
rect 140130 128256 140136 128268
rect 140188 128256 140194 128308
rect 227898 127644 227904 127696
rect 227956 127684 227962 127696
rect 267826 127684 267832 127696
rect 227956 127656 267832 127684
rect 227956 127644 227962 127656
rect 267826 127644 267832 127656
rect 267884 127644 267890 127696
rect 109126 127576 109132 127628
rect 109184 127616 109190 127628
rect 133230 127616 133236 127628
rect 109184 127588 133236 127616
rect 109184 127576 109190 127588
rect 133230 127576 133236 127588
rect 133288 127576 133294 127628
rect 158070 127576 158076 127628
rect 158128 127616 158134 127628
rect 183462 127616 183468 127628
rect 158128 127588 183468 127616
rect 158128 127576 158134 127588
rect 183462 127576 183468 127588
rect 183520 127576 183526 127628
rect 226702 127576 226708 127628
rect 226760 127616 226766 127628
rect 340874 127616 340880 127628
rect 226760 127588 340880 127616
rect 226760 127576 226766 127588
rect 340874 127576 340880 127588
rect 340932 127576 340938 127628
rect 183462 126964 183468 127016
rect 183520 127004 183526 127016
rect 191742 127004 191748 127016
rect 183520 126976 191748 127004
rect 183520 126964 183526 126976
rect 191742 126964 191748 126976
rect 191800 126964 191806 127016
rect 64506 126896 64512 126948
rect 64564 126936 64570 126948
rect 66806 126936 66812 126948
rect 64564 126908 66812 126936
rect 64564 126896 64570 126908
rect 66806 126896 66812 126908
rect 66864 126896 66870 126948
rect 226702 126896 226708 126948
rect 226760 126936 226766 126948
rect 249794 126936 249800 126948
rect 226760 126908 249800 126936
rect 226760 126896 226766 126908
rect 249794 126896 249800 126908
rect 249852 126936 249858 126948
rect 251082 126936 251088 126948
rect 249852 126908 251088 126936
rect 249852 126896 249858 126908
rect 251082 126896 251088 126908
rect 251140 126896 251146 126948
rect 97902 126828 97908 126880
rect 97960 126868 97966 126880
rect 103698 126868 103704 126880
rect 97960 126840 103704 126868
rect 97960 126828 97966 126840
rect 103698 126828 103704 126840
rect 103756 126828 103762 126880
rect 97166 126216 97172 126268
rect 97224 126256 97230 126268
rect 109126 126256 109132 126268
rect 97224 126228 109132 126256
rect 97224 126216 97230 126228
rect 109126 126216 109132 126228
rect 109184 126216 109190 126268
rect 179230 126216 179236 126268
rect 179288 126256 179294 126268
rect 187510 126256 187516 126268
rect 179288 126228 187516 126256
rect 179288 126216 179294 126228
rect 187510 126216 187516 126228
rect 187568 126256 187574 126268
rect 191558 126256 191564 126268
rect 187568 126228 191564 126256
rect 187568 126216 187574 126228
rect 191558 126216 191564 126228
rect 191616 126216 191622 126268
rect 251082 126216 251088 126268
rect 251140 126256 251146 126268
rect 351914 126256 351920 126268
rect 251140 126228 351920 126256
rect 251140 126216 251146 126228
rect 351914 126216 351920 126228
rect 351972 126216 351978 126268
rect 97902 125536 97908 125588
rect 97960 125576 97966 125588
rect 155402 125576 155408 125588
rect 97960 125548 155408 125576
rect 97960 125536 97966 125548
rect 155402 125536 155408 125548
rect 155460 125536 155466 125588
rect 155862 125536 155868 125588
rect 155920 125576 155926 125588
rect 156690 125576 156696 125588
rect 155920 125548 156696 125576
rect 155920 125536 155926 125548
rect 156690 125536 156696 125548
rect 156748 125536 156754 125588
rect 167730 125536 167736 125588
rect 167788 125576 167794 125588
rect 190362 125576 190368 125588
rect 167788 125548 190368 125576
rect 167788 125536 167794 125548
rect 190362 125536 190368 125548
rect 190420 125536 190426 125588
rect 59262 124924 59268 124976
rect 59320 124964 59326 124976
rect 66806 124964 66812 124976
rect 59320 124936 66812 124964
rect 59320 124924 59326 124936
rect 66806 124924 66812 124936
rect 66864 124924 66870 124976
rect 57790 124856 57796 124908
rect 57848 124896 57854 124908
rect 66990 124896 66996 124908
rect 57848 124868 66996 124896
rect 57848 124856 57854 124868
rect 66990 124856 66996 124868
rect 67048 124856 67054 124908
rect 238110 124856 238116 124908
rect 238168 124896 238174 124908
rect 305638 124896 305644 124908
rect 238168 124868 305644 124896
rect 238168 124856 238174 124868
rect 305638 124856 305644 124868
rect 305696 124856 305702 124908
rect 97810 124788 97816 124840
rect 97868 124828 97874 124840
rect 100754 124828 100760 124840
rect 97868 124800 100760 124828
rect 97868 124788 97874 124800
rect 100754 124788 100760 124800
rect 100812 124788 100818 124840
rect 101582 124176 101588 124228
rect 101640 124216 101646 124228
rect 155862 124216 155868 124228
rect 101640 124188 155868 124216
rect 101640 124176 101646 124188
rect 155862 124176 155868 124188
rect 155920 124176 155926 124228
rect 60458 124108 60464 124160
rect 60516 124148 60522 124160
rect 66898 124148 66904 124160
rect 60516 124120 66904 124148
rect 60516 124108 60522 124120
rect 66898 124108 66904 124120
rect 66956 124108 66962 124160
rect 97902 124108 97908 124160
rect 97960 124148 97966 124160
rect 150434 124148 150440 124160
rect 97960 124120 150440 124148
rect 97960 124108 97966 124120
rect 150434 124108 150440 124120
rect 150492 124108 150498 124160
rect 160738 124108 160744 124160
rect 160796 124148 160802 124160
rect 180150 124148 180156 124160
rect 160796 124120 180156 124148
rect 160796 124108 160802 124120
rect 180150 124108 180156 124120
rect 180208 124108 180214 124160
rect 226702 124108 226708 124160
rect 226760 124148 226766 124160
rect 230566 124148 230572 124160
rect 226760 124120 230572 124148
rect 226760 124108 226766 124120
rect 230566 124108 230572 124120
rect 230624 124148 230630 124160
rect 279418 124148 279424 124160
rect 230624 124120 279424 124148
rect 230624 124108 230630 124120
rect 279418 124108 279424 124120
rect 279476 124148 279482 124160
rect 582834 124148 582840 124160
rect 279476 124120 582840 124148
rect 279476 124108 279482 124120
rect 582834 124108 582840 124120
rect 582892 124108 582898 124160
rect 175918 124040 175924 124092
rect 175976 124080 175982 124092
rect 191742 124080 191748 124092
rect 175976 124052 191748 124080
rect 175976 124040 175982 124052
rect 191742 124040 191748 124052
rect 191800 124040 191806 124092
rect 235258 123428 235264 123480
rect 235316 123468 235322 123480
rect 243538 123468 243544 123480
rect 235316 123440 243544 123468
rect 235316 123428 235322 123440
rect 243538 123428 243544 123440
rect 243596 123428 243602 123480
rect 63310 122748 63316 122800
rect 63368 122788 63374 122800
rect 66346 122788 66352 122800
rect 63368 122760 66352 122788
rect 63368 122748 63374 122760
rect 66346 122748 66352 122760
rect 66404 122748 66410 122800
rect 97902 122748 97908 122800
rect 97960 122788 97966 122800
rect 153930 122788 153936 122800
rect 97960 122760 153936 122788
rect 97960 122748 97966 122760
rect 153930 122748 153936 122760
rect 153988 122748 153994 122800
rect 226518 122748 226524 122800
rect 226576 122788 226582 122800
rect 240226 122788 240232 122800
rect 226576 122760 240232 122788
rect 226576 122748 226582 122760
rect 240226 122748 240232 122760
rect 240284 122748 240290 122800
rect 250530 122068 250536 122120
rect 250588 122108 250594 122120
rect 285674 122108 285680 122120
rect 250588 122080 285680 122108
rect 250588 122068 250594 122080
rect 285674 122068 285680 122080
rect 285732 122068 285738 122120
rect 189074 121592 189080 121644
rect 189132 121632 189138 121644
rect 191742 121632 191748 121644
rect 189132 121604 191748 121632
rect 189132 121592 189138 121604
rect 191742 121592 191748 121604
rect 191800 121592 191806 121644
rect 53742 121388 53748 121440
rect 53800 121428 53806 121440
rect 66898 121428 66904 121440
rect 53800 121400 66904 121428
rect 53800 121388 53806 121400
rect 66898 121388 66904 121400
rect 66956 121388 66962 121440
rect 131850 121388 131856 121440
rect 131908 121428 131914 121440
rect 188982 121428 188988 121440
rect 131908 121400 188988 121428
rect 131908 121388 131914 121400
rect 188982 121388 188988 121400
rect 189040 121428 189046 121440
rect 191006 121428 191012 121440
rect 189040 121400 191012 121428
rect 189040 121388 189046 121400
rect 191006 121388 191012 121400
rect 191064 121388 191070 121440
rect 226702 121388 226708 121440
rect 226760 121428 226766 121440
rect 234706 121428 234712 121440
rect 226760 121400 234712 121428
rect 226760 121388 226766 121400
rect 234706 121388 234712 121400
rect 234764 121388 234770 121440
rect 61930 121320 61936 121372
rect 61988 121360 61994 121372
rect 66806 121360 66812 121372
rect 61988 121332 66812 121360
rect 61988 121320 61994 121332
rect 66806 121320 66812 121332
rect 66864 121320 66870 121372
rect 97074 121320 97080 121372
rect 97132 121360 97138 121372
rect 145650 121360 145656 121372
rect 97132 121332 145656 121360
rect 97132 121320 97138 121332
rect 145650 121320 145656 121332
rect 145708 121320 145714 121372
rect 159542 121320 159548 121372
rect 159600 121360 159606 121372
rect 191190 121360 191196 121372
rect 159600 121332 191196 121360
rect 159600 121320 159606 121332
rect 191190 121320 191196 121332
rect 191248 121320 191254 121372
rect 240778 120776 240784 120828
rect 240836 120816 240842 120828
rect 252554 120816 252560 120828
rect 240836 120788 252560 120816
rect 240836 120776 240842 120788
rect 252554 120776 252560 120788
rect 252612 120776 252618 120828
rect 232498 120708 232504 120760
rect 232556 120748 232562 120760
rect 313274 120748 313280 120760
rect 232556 120720 313280 120748
rect 232556 120708 232562 120720
rect 313274 120708 313280 120720
rect 313332 120708 313338 120760
rect 96062 120300 96068 120352
rect 96120 120340 96126 120352
rect 98822 120340 98828 120352
rect 96120 120312 98828 120340
rect 96120 120300 96126 120312
rect 98822 120300 98828 120312
rect 98880 120300 98886 120352
rect 64690 120028 64696 120080
rect 64748 120068 64754 120080
rect 66806 120068 66812 120080
rect 64748 120040 66812 120068
rect 64748 120028 64754 120040
rect 66806 120028 66812 120040
rect 66864 120028 66870 120080
rect 97902 120028 97908 120080
rect 97960 120068 97966 120080
rect 112438 120068 112444 120080
rect 97960 120040 112444 120068
rect 97960 120028 97966 120040
rect 112438 120028 112444 120040
rect 112496 120028 112502 120080
rect 184290 120028 184296 120080
rect 184348 120068 184354 120080
rect 191742 120068 191748 120080
rect 184348 120040 191748 120068
rect 184348 120028 184354 120040
rect 191742 120028 191748 120040
rect 191800 120028 191806 120080
rect 59078 119960 59084 120012
rect 59136 120000 59142 120012
rect 66898 120000 66904 120012
rect 59136 119972 66904 120000
rect 59136 119960 59142 119972
rect 66898 119960 66904 119972
rect 66956 119960 66962 120012
rect 104158 119348 104164 119400
rect 104216 119388 104222 119400
rect 187694 119388 187700 119400
rect 104216 119360 187700 119388
rect 104216 119348 104222 119360
rect 187694 119348 187700 119360
rect 187752 119348 187758 119400
rect 284294 119348 284300 119400
rect 284352 119388 284358 119400
rect 289814 119388 289820 119400
rect 284352 119360 289820 119388
rect 284352 119348 284358 119360
rect 289814 119348 289820 119360
rect 289872 119348 289878 119400
rect 52270 118600 52276 118652
rect 52328 118640 52334 118652
rect 66622 118640 66628 118652
rect 52328 118612 66628 118640
rect 52328 118600 52334 118612
rect 66622 118600 66628 118612
rect 66680 118600 66686 118652
rect 97902 118600 97908 118652
rect 97960 118640 97966 118652
rect 134702 118640 134708 118652
rect 97960 118612 134708 118640
rect 97960 118600 97966 118612
rect 134702 118600 134708 118612
rect 134760 118600 134766 118652
rect 186130 118600 186136 118652
rect 186188 118640 186194 118652
rect 188982 118640 188988 118652
rect 186188 118612 188988 118640
rect 186188 118600 186194 118612
rect 188982 118600 188988 118612
rect 189040 118600 189046 118652
rect 167638 117920 167644 117972
rect 167696 117960 167702 117972
rect 191742 117960 191748 117972
rect 167696 117932 191748 117960
rect 167696 117920 167702 117932
rect 191742 117920 191748 117932
rect 191800 117920 191806 117972
rect 226518 117376 226524 117428
rect 226576 117416 226582 117428
rect 231118 117416 231124 117428
rect 226576 117388 231124 117416
rect 226576 117376 226582 117388
rect 231118 117376 231124 117388
rect 231176 117376 231182 117428
rect 99466 117308 99472 117360
rect 99524 117348 99530 117360
rect 100662 117348 100668 117360
rect 99524 117320 100668 117348
rect 99524 117308 99530 117320
rect 100662 117308 100668 117320
rect 100720 117348 100726 117360
rect 160738 117348 160744 117360
rect 100720 117320 160744 117348
rect 100720 117308 100726 117320
rect 160738 117308 160744 117320
rect 160796 117308 160802 117360
rect 226610 117308 226616 117360
rect 226668 117348 226674 117360
rect 244274 117348 244280 117360
rect 226668 117320 244280 117348
rect 226668 117308 226674 117320
rect 244274 117308 244280 117320
rect 244332 117308 244338 117360
rect 62022 117240 62028 117292
rect 62080 117280 62086 117292
rect 66622 117280 66628 117292
rect 62080 117252 66628 117280
rect 62080 117240 62086 117252
rect 66622 117240 66628 117252
rect 66680 117240 66686 117292
rect 97350 117240 97356 117292
rect 97408 117280 97414 117292
rect 178862 117280 178868 117292
rect 97408 117252 178868 117280
rect 97408 117240 97414 117252
rect 178862 117240 178868 117252
rect 178920 117240 178926 117292
rect 97902 117172 97908 117224
rect 97960 117212 97966 117224
rect 177482 117212 177488 117224
rect 97960 117184 177488 117212
rect 97960 117172 97966 117184
rect 177482 117172 177488 117184
rect 177540 117172 177546 117224
rect 230382 116628 230388 116680
rect 230440 116668 230446 116680
rect 262398 116668 262404 116680
rect 230440 116640 262404 116668
rect 230440 116628 230446 116640
rect 262398 116628 262404 116640
rect 262456 116628 262462 116680
rect 245010 116560 245016 116612
rect 245068 116600 245074 116612
rect 285674 116600 285680 116612
rect 245068 116572 285680 116600
rect 245068 116560 245074 116572
rect 285674 116560 285680 116572
rect 285732 116560 285738 116612
rect 188430 116084 188436 116136
rect 188488 116124 188494 116136
rect 191558 116124 191564 116136
rect 188488 116096 191564 116124
rect 188488 116084 188494 116096
rect 191558 116084 191564 116096
rect 191616 116084 191622 116136
rect 226702 115948 226708 116000
rect 226760 115988 226766 116000
rect 229186 115988 229192 116000
rect 226760 115960 229192 115988
rect 226760 115948 226766 115960
rect 229186 115948 229192 115960
rect 229244 115988 229250 116000
rect 230382 115988 230388 116000
rect 229244 115960 230388 115988
rect 229244 115948 229250 115960
rect 230382 115948 230388 115960
rect 230440 115948 230446 116000
rect 50890 115880 50896 115932
rect 50948 115920 50954 115932
rect 66806 115920 66812 115932
rect 50948 115892 66812 115920
rect 50948 115880 50954 115892
rect 66806 115880 66812 115892
rect 66864 115880 66870 115932
rect 97810 115880 97816 115932
rect 97868 115920 97874 115932
rect 99466 115920 99472 115932
rect 97868 115892 99472 115920
rect 97868 115880 97874 115892
rect 99466 115880 99472 115892
rect 99524 115880 99530 115932
rect 226150 115880 226156 115932
rect 226208 115920 226214 115932
rect 280154 115920 280160 115932
rect 226208 115892 280160 115920
rect 226208 115880 226214 115892
rect 280154 115880 280160 115892
rect 280212 115880 280218 115932
rect 186222 115608 186228 115660
rect 186280 115648 186286 115660
rect 191742 115648 191748 115660
rect 186280 115620 191748 115648
rect 186280 115608 186286 115620
rect 191742 115608 191748 115620
rect 191800 115608 191806 115660
rect 63402 115540 63408 115592
rect 63460 115580 63466 115592
rect 66898 115580 66904 115592
rect 63460 115552 66904 115580
rect 63460 115540 63466 115552
rect 66898 115540 66904 115552
rect 66956 115540 66962 115592
rect 97902 114520 97908 114572
rect 97960 114560 97966 114572
rect 188338 114560 188344 114572
rect 97960 114532 188344 114560
rect 97960 114520 97966 114532
rect 188338 114520 188344 114532
rect 188396 114520 188402 114572
rect 60550 114452 60556 114504
rect 60608 114492 60614 114504
rect 66806 114492 66812 114504
rect 60608 114464 66812 114492
rect 60608 114452 60614 114464
rect 66806 114452 66812 114464
rect 66864 114452 66870 114504
rect 187694 114452 187700 114504
rect 187752 114492 187758 114504
rect 191742 114492 191748 114504
rect 187752 114464 191748 114492
rect 187752 114452 187758 114464
rect 191742 114452 191748 114464
rect 191800 114452 191806 114504
rect 226426 113840 226432 113892
rect 226484 113880 226490 113892
rect 250530 113880 250536 113892
rect 226484 113852 250536 113880
rect 226484 113840 226490 113852
rect 250530 113840 250536 113852
rect 250588 113840 250594 113892
rect 7558 113772 7564 113824
rect 7616 113812 7622 113824
rect 63402 113812 63408 113824
rect 7616 113784 63408 113812
rect 7616 113772 7622 113784
rect 63402 113772 63408 113784
rect 63460 113812 63466 113824
rect 66898 113812 66904 113824
rect 63460 113784 66904 113812
rect 63460 113772 63466 113784
rect 66898 113772 66904 113784
rect 66956 113772 66962 113824
rect 110506 113772 110512 113824
rect 110564 113812 110570 113824
rect 134610 113812 134616 113824
rect 110564 113784 134616 113812
rect 110564 113772 110570 113784
rect 134610 113772 134616 113784
rect 134668 113772 134674 113824
rect 246390 113772 246396 113824
rect 246448 113812 246454 113824
rect 270494 113812 270500 113824
rect 246448 113784 270500 113812
rect 246448 113772 246454 113784
rect 270494 113772 270500 113784
rect 270552 113772 270558 113824
rect 97534 113160 97540 113212
rect 97592 113200 97598 113212
rect 169018 113200 169024 113212
rect 97592 113172 169024 113200
rect 97592 113160 97598 113172
rect 169018 113160 169024 113172
rect 169076 113160 169082 113212
rect 55122 113092 55128 113144
rect 55180 113132 55186 113144
rect 66806 113132 66812 113144
rect 55180 113104 66812 113132
rect 55180 113092 55186 113104
rect 66806 113092 66812 113104
rect 66864 113092 66870 113144
rect 169662 112412 169668 112464
rect 169720 112452 169726 112464
rect 191742 112452 191748 112464
rect 169720 112424 191748 112452
rect 169720 112412 169726 112424
rect 191742 112412 191748 112424
rect 191800 112412 191806 112464
rect 225690 112412 225696 112464
rect 225748 112452 225754 112464
rect 252554 112452 252560 112464
rect 225748 112424 252560 112452
rect 225748 112412 225754 112424
rect 252554 112412 252560 112424
rect 252612 112452 252618 112464
rect 269114 112452 269120 112464
rect 252612 112424 269120 112452
rect 252612 112412 252618 112424
rect 269114 112412 269120 112424
rect 269172 112412 269178 112464
rect 96706 111868 96712 111920
rect 96764 111908 96770 111920
rect 98638 111908 98644 111920
rect 96764 111880 98644 111908
rect 96764 111868 96770 111880
rect 98638 111868 98644 111880
rect 98696 111868 98702 111920
rect 102042 111868 102048 111920
rect 102100 111908 102106 111920
rect 166258 111908 166264 111920
rect 102100 111880 166264 111908
rect 102100 111868 102106 111880
rect 166258 111868 166264 111880
rect 166316 111868 166322 111920
rect 169110 111868 169116 111920
rect 169168 111908 169174 111920
rect 169662 111908 169668 111920
rect 169168 111880 169668 111908
rect 169168 111868 169174 111880
rect 169662 111868 169668 111880
rect 169720 111868 169726 111920
rect 97902 111800 97908 111852
rect 97960 111840 97966 111852
rect 189718 111840 189724 111852
rect 97960 111812 189724 111840
rect 97960 111800 97966 111812
rect 189718 111800 189724 111812
rect 189776 111800 189782 111852
rect 226334 111800 226340 111852
rect 226392 111840 226398 111852
rect 231946 111840 231952 111852
rect 226392 111812 231952 111840
rect 226392 111800 226398 111812
rect 231946 111800 231952 111812
rect 232004 111840 232010 111852
rect 295334 111840 295340 111852
rect 232004 111812 295340 111840
rect 232004 111800 232010 111812
rect 295334 111800 295340 111812
rect 295392 111800 295398 111852
rect 43990 111732 43996 111784
rect 44048 111772 44054 111784
rect 66806 111772 66812 111784
rect 44048 111744 66812 111772
rect 44048 111732 44054 111744
rect 66806 111732 66812 111744
rect 66864 111732 66870 111784
rect 185578 111732 185584 111784
rect 185636 111772 185642 111784
rect 191742 111772 191748 111784
rect 185636 111744 191748 111772
rect 185636 111732 185642 111744
rect 191742 111732 191748 111744
rect 191800 111732 191806 111784
rect 226702 111528 226708 111580
rect 226760 111568 226766 111580
rect 230474 111568 230480 111580
rect 226760 111540 230480 111568
rect 226760 111528 226766 111540
rect 230474 111528 230480 111540
rect 230532 111528 230538 111580
rect 96798 111120 96804 111172
rect 96856 111160 96862 111172
rect 100018 111160 100024 111172
rect 96856 111132 100024 111160
rect 96856 111120 96862 111132
rect 100018 111120 100024 111132
rect 100076 111120 100082 111172
rect 39942 111052 39948 111104
rect 40000 111092 40006 111104
rect 59262 111092 59268 111104
rect 40000 111064 59268 111092
rect 40000 111052 40006 111064
rect 59262 111052 59268 111064
rect 59320 111092 59326 111104
rect 66898 111092 66904 111104
rect 59320 111064 66904 111092
rect 59320 111052 59326 111064
rect 66898 111052 66904 111064
rect 66956 111052 66962 111104
rect 100110 111052 100116 111104
rect 100168 111092 100174 111104
rect 188430 111092 188436 111104
rect 100168 111064 188436 111092
rect 100168 111052 100174 111064
rect 188430 111052 188436 111064
rect 188488 111052 188494 111104
rect 226334 111052 226340 111104
rect 226392 111092 226398 111104
rect 226392 111064 277394 111092
rect 226392 111052 226398 111064
rect 277366 111024 277394 111064
rect 295334 111052 295340 111104
rect 295392 111092 295398 111104
rect 324314 111092 324320 111104
rect 295392 111064 324320 111092
rect 295392 111052 295398 111064
rect 324314 111052 324320 111064
rect 324372 111052 324378 111104
rect 295426 111024 295432 111036
rect 277366 110996 295432 111024
rect 295426 110984 295432 110996
rect 295484 110984 295490 111036
rect 2866 110780 2872 110832
rect 2924 110820 2930 110832
rect 4798 110820 4804 110832
rect 2924 110792 4804 110820
rect 2924 110780 2930 110792
rect 4798 110780 4804 110792
rect 4856 110780 4862 110832
rect 190362 110440 190368 110492
rect 190420 110480 190426 110492
rect 191834 110480 191840 110492
rect 190420 110452 191840 110480
rect 190420 110440 190426 110452
rect 191834 110440 191840 110452
rect 191892 110440 191898 110492
rect 295426 110440 295432 110492
rect 295484 110480 295490 110492
rect 295978 110480 295984 110492
rect 295484 110452 295984 110480
rect 295484 110440 295490 110452
rect 295978 110440 295984 110452
rect 296036 110440 296042 110492
rect 97810 110372 97816 110424
rect 97868 110412 97874 110424
rect 102042 110412 102048 110424
rect 97868 110384 102048 110412
rect 97868 110372 97874 110384
rect 102042 110372 102048 110384
rect 102100 110372 102106 110424
rect 111150 110372 111156 110424
rect 111208 110412 111214 110424
rect 190638 110412 190644 110424
rect 111208 110384 190644 110412
rect 111208 110372 111214 110384
rect 190638 110372 190644 110384
rect 190696 110372 190702 110424
rect 231118 110372 231124 110424
rect 231176 110412 231182 110424
rect 299658 110412 299664 110424
rect 231176 110384 299664 110412
rect 231176 110372 231182 110384
rect 299658 110372 299664 110384
rect 299716 110412 299722 110424
rect 307018 110412 307024 110424
rect 299716 110384 307024 110412
rect 299716 110372 299722 110384
rect 307018 110372 307024 110384
rect 307076 110372 307082 110424
rect 97902 110304 97908 110356
rect 97960 110344 97966 110356
rect 173250 110344 173256 110356
rect 97960 110316 173256 110344
rect 97960 110304 97966 110316
rect 173250 110304 173256 110316
rect 173308 110304 173314 110356
rect 48222 109012 48228 109064
rect 48280 109052 48286 109064
rect 53834 109052 53840 109064
rect 48280 109024 53840 109052
rect 48280 109012 48286 109024
rect 53834 109012 53840 109024
rect 53892 109052 53898 109064
rect 66898 109052 66904 109064
rect 53892 109024 66904 109052
rect 53892 109012 53898 109024
rect 66898 109012 66904 109024
rect 66956 109012 66962 109064
rect 54938 108944 54944 108996
rect 54996 108984 55002 108996
rect 66806 108984 66812 108996
rect 54996 108956 66812 108984
rect 54996 108944 55002 108956
rect 66806 108944 66812 108956
rect 66864 108944 66870 108996
rect 165522 108944 165528 108996
rect 165580 108984 165586 108996
rect 189074 108984 189080 108996
rect 165580 108956 189080 108984
rect 165580 108944 165586 108956
rect 189074 108944 189080 108956
rect 189132 108944 189138 108996
rect 187602 108876 187608 108928
rect 187660 108916 187666 108928
rect 191742 108916 191748 108928
rect 187660 108888 191748 108916
rect 187660 108876 187666 108888
rect 191742 108876 191748 108888
rect 191800 108876 191806 108928
rect 226518 108876 226524 108928
rect 226576 108916 226582 108928
rect 229094 108916 229100 108928
rect 226576 108888 229100 108916
rect 226576 108876 226582 108888
rect 229094 108876 229100 108888
rect 229152 108876 229158 108928
rect 98822 108332 98828 108384
rect 98880 108372 98886 108384
rect 113266 108372 113272 108384
rect 98880 108344 113272 108372
rect 98880 108332 98886 108344
rect 113266 108332 113272 108344
rect 113324 108332 113330 108384
rect 97902 108264 97908 108316
rect 97960 108304 97966 108316
rect 109034 108304 109040 108316
rect 97960 108276 109040 108304
rect 97960 108264 97966 108276
rect 109034 108264 109040 108276
rect 109092 108304 109098 108316
rect 109678 108304 109684 108316
rect 109092 108276 109684 108304
rect 109092 108264 109098 108276
rect 109678 108264 109684 108276
rect 109736 108264 109742 108316
rect 112438 108264 112444 108316
rect 112496 108304 112502 108316
rect 165522 108304 165528 108316
rect 112496 108276 165528 108304
rect 112496 108264 112502 108276
rect 165522 108264 165528 108276
rect 165580 108264 165586 108316
rect 226978 108264 226984 108316
rect 227036 108304 227042 108316
rect 263686 108304 263692 108316
rect 227036 108276 263692 108304
rect 227036 108264 227042 108276
rect 263686 108264 263692 108276
rect 263744 108264 263750 108316
rect 64598 107584 64604 107636
rect 64656 107624 64662 107636
rect 66622 107624 66628 107636
rect 64656 107596 66628 107624
rect 64656 107584 64662 107596
rect 66622 107584 66628 107596
rect 66680 107584 66686 107636
rect 97902 107584 97908 107636
rect 97960 107624 97966 107636
rect 177390 107624 177396 107636
rect 97960 107596 177396 107624
rect 97960 107584 97966 107596
rect 177390 107584 177396 107596
rect 177448 107584 177454 107636
rect 182818 107584 182824 107636
rect 182876 107624 182882 107636
rect 190822 107624 190828 107636
rect 182876 107596 190828 107624
rect 182876 107584 182882 107596
rect 190822 107584 190828 107596
rect 190880 107584 190886 107636
rect 226702 107584 226708 107636
rect 226760 107624 226766 107636
rect 285766 107624 285772 107636
rect 226760 107596 285772 107624
rect 226760 107584 226766 107596
rect 285766 107584 285772 107596
rect 285824 107624 285830 107636
rect 286226 107624 286232 107636
rect 285824 107596 286232 107624
rect 285824 107584 285830 107596
rect 286226 107584 286232 107596
rect 286284 107584 286290 107636
rect 286226 106904 286232 106956
rect 286284 106944 286290 106956
rect 342898 106944 342904 106956
rect 286284 106916 342904 106944
rect 286284 106904 286290 106916
rect 342898 106904 342904 106916
rect 342956 106904 342962 106956
rect 97902 106496 97908 106548
rect 97960 106536 97966 106548
rect 101674 106536 101680 106548
rect 97960 106508 101680 106536
rect 97960 106496 97966 106508
rect 101674 106496 101680 106508
rect 101732 106496 101738 106548
rect 7558 106292 7564 106344
rect 7616 106332 7622 106344
rect 66806 106332 66812 106344
rect 7616 106304 66812 106332
rect 7616 106292 7622 106304
rect 66806 106292 66812 106304
rect 66864 106292 66870 106344
rect 160830 106224 160836 106276
rect 160888 106264 160894 106276
rect 191190 106264 191196 106276
rect 160888 106236 191196 106264
rect 160888 106224 160894 106236
rect 191190 106224 191196 106236
rect 191248 106224 191254 106276
rect 46842 105544 46848 105596
rect 46900 105584 46906 105596
rect 66162 105584 66168 105596
rect 46900 105556 66168 105584
rect 46900 105544 46906 105556
rect 66162 105544 66168 105556
rect 66220 105584 66226 105596
rect 66622 105584 66628 105596
rect 66220 105556 66628 105584
rect 66220 105544 66226 105556
rect 66622 105544 66628 105556
rect 66680 105544 66686 105596
rect 106182 105544 106188 105596
rect 106240 105584 106246 105596
rect 120166 105584 120172 105596
rect 106240 105556 120172 105584
rect 106240 105544 106246 105556
rect 120166 105544 120172 105556
rect 120224 105584 120230 105596
rect 177390 105584 177396 105596
rect 120224 105556 177396 105584
rect 120224 105544 120230 105556
rect 177390 105544 177396 105556
rect 177448 105544 177454 105596
rect 178678 105544 178684 105596
rect 178736 105584 178742 105596
rect 187602 105584 187608 105596
rect 178736 105556 187608 105584
rect 178736 105544 178742 105556
rect 187602 105544 187608 105556
rect 187660 105584 187666 105596
rect 191742 105584 191748 105596
rect 187660 105556 191748 105584
rect 187660 105544 187666 105556
rect 191742 105544 191748 105556
rect 191800 105544 191806 105596
rect 226334 105544 226340 105596
rect 226392 105584 226398 105596
rect 240778 105584 240784 105596
rect 226392 105556 240784 105584
rect 226392 105544 226398 105556
rect 240778 105544 240784 105556
rect 240836 105544 240842 105596
rect 245010 105544 245016 105596
rect 245068 105584 245074 105596
rect 273254 105584 273260 105596
rect 245068 105556 273260 105584
rect 245068 105544 245074 105556
rect 273254 105544 273260 105556
rect 273312 105544 273318 105596
rect 226702 105000 226708 105052
rect 226760 105040 226766 105052
rect 230566 105040 230572 105052
rect 226760 105012 230572 105040
rect 226760 105000 226766 105012
rect 230566 105000 230572 105012
rect 230624 105000 230630 105052
rect 56502 104796 56508 104848
rect 56560 104836 56566 104848
rect 66806 104836 66812 104848
rect 56560 104808 66812 104836
rect 56560 104796 56566 104808
rect 66806 104796 66812 104808
rect 66864 104796 66870 104848
rect 101306 104796 101312 104848
rect 101364 104836 101370 104848
rect 101490 104836 101496 104848
rect 101364 104808 101496 104836
rect 101364 104796 101370 104808
rect 101490 104796 101496 104808
rect 101548 104796 101554 104848
rect 270402 104796 270408 104848
rect 270460 104836 270466 104848
rect 274634 104836 274640 104848
rect 270460 104808 274640 104836
rect 270460 104796 270466 104808
rect 274634 104796 274640 104808
rect 274692 104796 274698 104848
rect 97902 104184 97908 104236
rect 97960 104224 97966 104236
rect 106182 104224 106188 104236
rect 97960 104196 106188 104224
rect 97960 104184 97966 104196
rect 106182 104184 106188 104196
rect 106240 104184 106246 104236
rect 225690 104116 225696 104168
rect 225748 104156 225754 104168
rect 255958 104156 255964 104168
rect 225748 104128 255964 104156
rect 225748 104116 225754 104128
rect 255958 104116 255964 104128
rect 256016 104116 256022 104168
rect 185578 103544 185584 103556
rect 101416 103516 185584 103544
rect 97902 103436 97908 103488
rect 97960 103476 97966 103488
rect 101306 103476 101312 103488
rect 97960 103448 101312 103476
rect 97960 103436 97966 103448
rect 101306 103436 101312 103448
rect 101364 103476 101370 103488
rect 101416 103476 101444 103516
rect 185578 103504 185584 103516
rect 185636 103504 185642 103556
rect 226702 103504 226708 103556
rect 226760 103544 226766 103556
rect 229094 103544 229100 103556
rect 226760 103516 229100 103544
rect 226760 103504 226766 103516
rect 229094 103504 229100 103516
rect 229152 103544 229158 103556
rect 270402 103544 270408 103556
rect 229152 103516 270408 103544
rect 229152 103504 229158 103516
rect 270402 103504 270408 103516
rect 270460 103504 270466 103556
rect 101364 103448 101444 103476
rect 101364 103436 101370 103448
rect 55030 103368 55036 103420
rect 55088 103408 55094 103420
rect 66438 103408 66444 103420
rect 55088 103380 66444 103408
rect 55088 103368 55094 103380
rect 66438 103368 66444 103380
rect 66496 103368 66502 103420
rect 97902 103028 97908 103080
rect 97960 103068 97966 103080
rect 99374 103068 99380 103080
rect 97960 103040 99380 103068
rect 97960 103028 97966 103040
rect 99374 103028 99380 103040
rect 99432 103028 99438 103080
rect 99374 102756 99380 102808
rect 99432 102796 99438 102808
rect 182818 102796 182824 102808
rect 99432 102768 182824 102796
rect 99432 102756 99438 102768
rect 182818 102756 182824 102768
rect 182876 102756 182882 102808
rect 226702 102756 226708 102808
rect 226760 102796 226766 102808
rect 230474 102796 230480 102808
rect 226760 102768 230480 102796
rect 226760 102756 226766 102768
rect 230474 102756 230480 102768
rect 230532 102796 230538 102808
rect 282914 102796 282920 102808
rect 230532 102768 282920 102796
rect 230532 102756 230538 102768
rect 282914 102756 282920 102768
rect 282972 102796 282978 102808
rect 321646 102796 321652 102808
rect 282972 102768 321652 102796
rect 282972 102756 282978 102768
rect 321646 102756 321652 102768
rect 321704 102756 321710 102808
rect 188522 102144 188528 102196
rect 188580 102184 188586 102196
rect 191006 102184 191012 102196
rect 188580 102156 191012 102184
rect 188580 102144 188586 102156
rect 191006 102144 191012 102156
rect 191064 102144 191070 102196
rect 226702 102144 226708 102196
rect 226760 102184 226766 102196
rect 237374 102184 237380 102196
rect 226760 102156 237380 102184
rect 226760 102144 226766 102156
rect 237374 102144 237380 102156
rect 237432 102144 237438 102196
rect 97902 102076 97908 102128
rect 97960 102116 97966 102128
rect 129182 102116 129188 102128
rect 97960 102088 129188 102116
rect 97960 102076 97966 102088
rect 129182 102076 129188 102088
rect 129240 102076 129246 102128
rect 226334 102076 226340 102128
rect 226392 102116 226398 102128
rect 266446 102116 266452 102128
rect 226392 102088 266452 102116
rect 226392 102076 226398 102088
rect 266446 102076 266452 102088
rect 266504 102076 266510 102128
rect 166902 101464 166908 101516
rect 166960 101504 166966 101516
rect 180794 101504 180800 101516
rect 166960 101476 180800 101504
rect 166960 101464 166966 101476
rect 180794 101464 180800 101476
rect 180852 101504 180858 101516
rect 181898 101504 181904 101516
rect 180852 101476 181904 101504
rect 180852 101464 180858 101476
rect 181898 101464 181904 101476
rect 181956 101464 181962 101516
rect 55122 101396 55128 101448
rect 55180 101436 55186 101448
rect 59170 101436 59176 101448
rect 55180 101408 59176 101436
rect 55180 101396 55186 101408
rect 59170 101396 59176 101408
rect 59228 101436 59234 101448
rect 66714 101436 66720 101448
rect 59228 101408 66720 101436
rect 59228 101396 59234 101408
rect 66714 101396 66720 101408
rect 66772 101396 66778 101448
rect 104158 101396 104164 101448
rect 104216 101436 104222 101448
rect 117406 101436 117412 101448
rect 104216 101408 117412 101436
rect 104216 101396 104222 101408
rect 117406 101396 117412 101408
rect 117464 101396 117470 101448
rect 129182 101396 129188 101448
rect 129240 101436 129246 101448
rect 153930 101436 153936 101448
rect 129240 101408 153936 101436
rect 129240 101396 129246 101408
rect 153930 101396 153936 101408
rect 153988 101396 153994 101448
rect 155862 101396 155868 101448
rect 155920 101436 155926 101448
rect 186958 101436 186964 101448
rect 155920 101408 186964 101436
rect 155920 101396 155926 101408
rect 186958 101396 186964 101408
rect 187016 101396 187022 101448
rect 226702 101396 226708 101448
rect 226760 101436 226766 101448
rect 277394 101436 277400 101448
rect 226760 101408 277400 101436
rect 226760 101396 226766 101408
rect 277394 101396 277400 101408
rect 277452 101396 277458 101448
rect 64690 100716 64696 100768
rect 64748 100756 64754 100768
rect 66806 100756 66812 100768
rect 64748 100728 66812 100756
rect 64748 100716 64754 100728
rect 66806 100716 66812 100728
rect 66864 100716 66870 100768
rect 120718 100716 120724 100768
rect 120776 100756 120782 100768
rect 163498 100756 163504 100768
rect 120776 100728 163504 100756
rect 120776 100716 120782 100728
rect 163498 100716 163504 100728
rect 163556 100756 163562 100768
rect 164142 100756 164148 100768
rect 163556 100728 164148 100756
rect 163556 100716 163562 100728
rect 164142 100716 164148 100728
rect 164200 100716 164206 100768
rect 181898 100716 181904 100768
rect 181956 100756 181962 100768
rect 191742 100756 191748 100768
rect 181956 100728 191748 100756
rect 181956 100716 181962 100728
rect 191742 100716 191748 100728
rect 191800 100716 191806 100768
rect 97902 99968 97908 100020
rect 97960 100008 97966 100020
rect 101398 100008 101404 100020
rect 97960 99980 101404 100008
rect 97960 99968 97966 99980
rect 101398 99968 101404 99980
rect 101456 100008 101462 100020
rect 185670 100008 185676 100020
rect 101456 99980 185676 100008
rect 101456 99968 101462 99980
rect 185670 99968 185676 99980
rect 185728 99968 185734 100020
rect 64782 99628 64788 99680
rect 64840 99668 64846 99680
rect 66806 99668 66812 99680
rect 64840 99640 66812 99668
rect 64840 99628 64846 99640
rect 66806 99628 66812 99640
rect 66864 99628 66870 99680
rect 97534 99356 97540 99408
rect 97592 99396 97598 99408
rect 129642 99396 129648 99408
rect 97592 99368 129648 99396
rect 97592 99356 97598 99368
rect 129642 99356 129648 99368
rect 129700 99356 129706 99408
rect 226334 99356 226340 99408
rect 226392 99396 226398 99408
rect 327718 99396 327724 99408
rect 226392 99368 327724 99396
rect 226392 99356 226398 99368
rect 327718 99356 327724 99368
rect 327776 99356 327782 99408
rect 53650 99288 53656 99340
rect 53708 99328 53714 99340
rect 66806 99328 66812 99340
rect 53708 99300 66812 99328
rect 53708 99288 53714 99300
rect 66806 99288 66812 99300
rect 66864 99288 66870 99340
rect 271874 99288 271880 99340
rect 271932 99328 271938 99340
rect 580166 99328 580172 99340
rect 271932 99300 580172 99328
rect 271932 99288 271938 99300
rect 580166 99288 580172 99300
rect 580224 99288 580230 99340
rect 246482 98744 246488 98796
rect 246540 98784 246546 98796
rect 269298 98784 269304 98796
rect 246540 98756 269304 98784
rect 246540 98744 246546 98756
rect 269298 98744 269304 98756
rect 269356 98744 269362 98796
rect 262858 98676 262864 98728
rect 262916 98716 262922 98728
rect 271874 98716 271880 98728
rect 262916 98688 271880 98716
rect 262916 98676 262922 98688
rect 271874 98676 271880 98688
rect 271932 98676 271938 98728
rect 97534 98608 97540 98660
rect 97592 98648 97598 98660
rect 107746 98648 107752 98660
rect 97592 98620 107752 98648
rect 97592 98608 97598 98620
rect 107746 98608 107752 98620
rect 107804 98608 107810 98660
rect 226610 98608 226616 98660
rect 226668 98648 226674 98660
rect 237282 98648 237288 98660
rect 226668 98620 237288 98648
rect 226668 98608 226674 98620
rect 237282 98608 237288 98620
rect 237340 98648 237346 98660
rect 247678 98648 247684 98660
rect 237340 98620 247684 98648
rect 237340 98608 237346 98620
rect 247678 98608 247684 98620
rect 247736 98608 247742 98660
rect 184290 98064 184296 98116
rect 184348 98104 184354 98116
rect 191742 98104 191748 98116
rect 184348 98076 191748 98104
rect 184348 98064 184354 98076
rect 191742 98064 191748 98076
rect 191800 98064 191806 98116
rect 97902 97996 97908 98048
rect 97960 98036 97966 98048
rect 188798 98036 188804 98048
rect 97960 98008 188804 98036
rect 97960 97996 97966 98008
rect 188798 97996 188804 98008
rect 188856 97996 188862 98048
rect 180242 97928 180248 97980
rect 180300 97968 180306 97980
rect 191650 97968 191656 97980
rect 180300 97940 191656 97968
rect 180300 97928 180306 97940
rect 191650 97928 191656 97940
rect 191708 97928 191714 97980
rect 101398 97248 101404 97300
rect 101456 97288 101462 97300
rect 169110 97288 169116 97300
rect 101456 97260 169116 97288
rect 101456 97248 101462 97260
rect 169110 97248 169116 97260
rect 169168 97248 169174 97300
rect 227162 97248 227168 97300
rect 227220 97288 227226 97300
rect 263594 97288 263600 97300
rect 227220 97260 263600 97288
rect 227220 97248 227226 97260
rect 263594 97248 263600 97260
rect 263652 97248 263658 97300
rect 96706 96976 96712 97028
rect 96764 97016 96770 97028
rect 98730 97016 98736 97028
rect 96764 96988 98736 97016
rect 96764 96976 96770 96988
rect 98730 96976 98736 96988
rect 98788 96976 98794 97028
rect 3050 96636 3056 96688
rect 3108 96676 3114 96688
rect 65518 96676 65524 96688
rect 3108 96648 65524 96676
rect 3108 96636 3114 96648
rect 65518 96636 65524 96648
rect 65576 96636 65582 96688
rect 99006 96636 99012 96688
rect 99064 96676 99070 96688
rect 114646 96676 114652 96688
rect 99064 96648 114652 96676
rect 99064 96636 99070 96648
rect 114646 96636 114652 96648
rect 114704 96676 114710 96688
rect 115842 96676 115848 96688
rect 114704 96648 115848 96676
rect 114704 96636 114710 96648
rect 115842 96636 115848 96648
rect 115900 96636 115906 96688
rect 226702 96568 226708 96620
rect 226760 96608 226766 96620
rect 264974 96608 264980 96620
rect 226760 96580 264980 96608
rect 226760 96568 226766 96580
rect 264974 96568 264980 96580
rect 265032 96568 265038 96620
rect 115842 95888 115848 95940
rect 115900 95928 115906 95940
rect 191926 95928 191932 95940
rect 115900 95900 191932 95928
rect 115900 95888 115906 95900
rect 191926 95888 191932 95900
rect 191984 95888 191990 95940
rect 227990 95888 227996 95940
rect 228048 95928 228054 95940
rect 244918 95928 244924 95940
rect 228048 95900 244924 95928
rect 228048 95888 228054 95900
rect 244918 95888 244924 95900
rect 244976 95888 244982 95940
rect 97902 95208 97908 95260
rect 97960 95248 97966 95260
rect 177482 95248 177488 95260
rect 97960 95220 177488 95248
rect 97960 95208 97966 95220
rect 177482 95208 177488 95220
rect 177540 95208 177546 95260
rect 57698 95140 57704 95192
rect 57756 95180 57762 95192
rect 66806 95180 66812 95192
rect 57756 95152 66812 95180
rect 57756 95140 57762 95152
rect 66806 95140 66812 95152
rect 66864 95140 66870 95192
rect 95970 94528 95976 94580
rect 96028 94568 96034 94580
rect 110598 94568 110604 94580
rect 96028 94540 110604 94568
rect 96028 94528 96034 94540
rect 110598 94528 110604 94540
rect 110656 94528 110662 94580
rect 94866 94460 94872 94512
rect 94924 94500 94930 94512
rect 124306 94500 124312 94512
rect 94924 94472 124312 94500
rect 94924 94460 94930 94472
rect 124306 94460 124312 94472
rect 124364 94500 124370 94512
rect 191834 94500 191840 94512
rect 124364 94472 191840 94500
rect 124364 94460 124370 94472
rect 191834 94460 191840 94472
rect 191892 94460 191898 94512
rect 158622 93848 158628 93900
rect 158680 93888 158686 93900
rect 192018 93888 192024 93900
rect 158680 93860 192024 93888
rect 158680 93848 158686 93860
rect 192018 93848 192024 93860
rect 192076 93848 192082 93900
rect 57882 93780 57888 93832
rect 57940 93820 57946 93832
rect 67174 93820 67180 93832
rect 57940 93792 67180 93820
rect 57940 93780 57946 93792
rect 67174 93780 67180 93792
rect 67232 93780 67238 93832
rect 67450 93780 67456 93832
rect 67508 93820 67514 93832
rect 67726 93820 67732 93832
rect 67508 93792 67732 93820
rect 67508 93780 67514 93792
rect 67726 93780 67732 93792
rect 67784 93780 67790 93832
rect 97902 93780 97908 93832
rect 97960 93820 97966 93832
rect 109218 93820 109224 93832
rect 97960 93792 109224 93820
rect 97960 93780 97966 93792
rect 109218 93780 109224 93792
rect 109276 93780 109282 93832
rect 224034 93372 224040 93424
rect 224092 93412 224098 93424
rect 225138 93412 225144 93424
rect 224092 93384 225144 93412
rect 224092 93372 224098 93384
rect 225138 93372 225144 93384
rect 225196 93372 225202 93424
rect 222102 93304 222108 93356
rect 222160 93344 222166 93356
rect 225690 93344 225696 93356
rect 222160 93316 225696 93344
rect 222160 93304 222166 93316
rect 225690 93304 225696 93316
rect 225748 93304 225754 93356
rect 247678 93100 247684 93152
rect 247736 93140 247742 93152
rect 331214 93140 331220 93152
rect 247736 93112 331220 93140
rect 247736 93100 247742 93112
rect 331214 93100 331220 93112
rect 331272 93100 331278 93152
rect 88656 92692 88662 92744
rect 88714 92732 88720 92744
rect 88714 92704 93854 92732
rect 88714 92692 88720 92704
rect 90128 92624 90134 92676
rect 90186 92664 90192 92676
rect 91002 92664 91008 92676
rect 90186 92636 91008 92664
rect 90186 92624 90192 92636
rect 91002 92624 91008 92636
rect 91060 92624 91066 92676
rect 93826 92664 93854 92704
rect 94866 92664 94872 92676
rect 93826 92636 94872 92664
rect 94866 92624 94872 92636
rect 94924 92624 94930 92676
rect 93808 92556 93814 92608
rect 93866 92596 93872 92608
rect 94498 92596 94504 92608
rect 93866 92568 94504 92596
rect 93866 92556 93872 92568
rect 94498 92556 94504 92568
rect 94556 92596 94562 92608
rect 95878 92596 95884 92608
rect 94556 92568 95884 92596
rect 94556 92556 94562 92568
rect 95878 92556 95884 92568
rect 95936 92556 95942 92608
rect 94682 92488 94688 92540
rect 94740 92528 94746 92540
rect 104158 92528 104164 92540
rect 94740 92500 104164 92528
rect 94740 92488 94746 92500
rect 104158 92488 104164 92500
rect 104216 92488 104222 92540
rect 191926 92488 191932 92540
rect 191984 92528 191990 92540
rect 207382 92528 207388 92540
rect 191984 92500 207388 92528
rect 191984 92488 191990 92500
rect 207382 92488 207388 92500
rect 207440 92488 207446 92540
rect 212902 92488 212908 92540
rect 212960 92528 212966 92540
rect 242250 92528 242256 92540
rect 212960 92500 242256 92528
rect 212960 92488 212966 92500
rect 242250 92488 242256 92500
rect 242308 92488 242314 92540
rect 67358 92420 67364 92472
rect 67416 92460 67422 92472
rect 184290 92460 184296 92472
rect 67416 92432 184296 92460
rect 67416 92420 67422 92432
rect 184290 92420 184296 92432
rect 184348 92420 184354 92472
rect 191834 92420 191840 92472
rect 191892 92460 191898 92472
rect 217134 92460 217140 92472
rect 191892 92432 217140 92460
rect 191892 92420 191898 92432
rect 217134 92420 217140 92432
rect 217192 92420 217198 92472
rect 224862 92420 224868 92472
rect 224920 92460 224926 92472
rect 227806 92460 227812 92472
rect 224920 92432 227812 92460
rect 224920 92420 224926 92432
rect 227806 92420 227812 92432
rect 227864 92420 227870 92472
rect 60642 92352 60648 92404
rect 60700 92392 60706 92404
rect 79410 92392 79416 92404
rect 60700 92364 79416 92392
rect 60700 92352 60706 92364
rect 79410 92352 79416 92364
rect 79468 92352 79474 92404
rect 80606 92352 80612 92404
rect 80664 92392 80670 92404
rect 99006 92392 99012 92404
rect 80664 92364 99012 92392
rect 80664 92352 80670 92364
rect 99006 92352 99012 92364
rect 99064 92352 99070 92404
rect 182082 92352 182088 92404
rect 182140 92392 182146 92404
rect 202598 92392 202604 92404
rect 182140 92364 202604 92392
rect 182140 92352 182146 92364
rect 202598 92352 202604 92364
rect 202656 92352 202662 92404
rect 213270 92352 213276 92404
rect 213328 92392 213334 92404
rect 226610 92392 226616 92404
rect 213328 92364 226616 92392
rect 213328 92352 213334 92364
rect 226610 92352 226616 92364
rect 226668 92352 226674 92404
rect 61838 90992 61844 91044
rect 61896 91032 61902 91044
rect 70302 91032 70308 91044
rect 61896 91004 70308 91032
rect 61896 90992 61902 91004
rect 70302 90992 70308 91004
rect 70360 90992 70366 91044
rect 78950 90992 78956 91044
rect 79008 91032 79014 91044
rect 111886 91032 111892 91044
rect 79008 91004 111892 91032
rect 79008 90992 79014 91004
rect 111886 90992 111892 91004
rect 111944 90992 111950 91044
rect 176562 90992 176568 91044
rect 176620 91032 176626 91044
rect 195974 91032 195980 91044
rect 176620 91004 195980 91032
rect 176620 90992 176626 91004
rect 195974 90992 195980 91004
rect 196032 90992 196038 91044
rect 217134 90992 217140 91044
rect 217192 91032 217198 91044
rect 246390 91032 246396 91044
rect 217192 91004 246396 91032
rect 217192 90992 217198 91004
rect 246390 90992 246396 91004
rect 246448 90992 246454 91044
rect 181990 90924 181996 90976
rect 182048 90964 182054 90976
rect 194686 90964 194692 90976
rect 182048 90936 194692 90964
rect 182048 90924 182054 90936
rect 194686 90924 194692 90936
rect 194744 90924 194750 90976
rect 221366 90924 221372 90976
rect 221424 90964 221430 90976
rect 225598 90964 225604 90976
rect 221424 90936 225604 90964
rect 221424 90924 221430 90936
rect 225598 90924 225604 90936
rect 225656 90924 225662 90976
rect 194686 90516 194692 90568
rect 194744 90556 194750 90568
rect 195238 90556 195244 90568
rect 194744 90528 195244 90556
rect 194744 90516 194750 90528
rect 195238 90516 195244 90528
rect 195296 90516 195302 90568
rect 223758 90516 223764 90568
rect 223816 90556 223822 90568
rect 224862 90556 224868 90568
rect 223816 90528 224868 90556
rect 223816 90516 223822 90528
rect 224862 90516 224868 90528
rect 224920 90516 224926 90568
rect 258718 90312 258724 90364
rect 258776 90352 258782 90364
rect 291194 90352 291200 90364
rect 258776 90324 291200 90352
rect 258776 90312 258782 90324
rect 291194 90312 291200 90324
rect 291252 90312 291258 90364
rect 70302 89700 70308 89752
rect 70360 89740 70366 89752
rect 73798 89740 73804 89752
rect 70360 89712 73804 89740
rect 70360 89700 70366 89712
rect 73798 89700 73804 89712
rect 73856 89700 73862 89752
rect 85206 89700 85212 89752
rect 85264 89740 85270 89752
rect 93118 89740 93124 89752
rect 85264 89712 93124 89740
rect 85264 89700 85270 89712
rect 93118 89700 93124 89712
rect 93176 89700 93182 89752
rect 63402 89632 63408 89684
rect 63460 89672 63466 89684
rect 100110 89672 100116 89684
rect 63460 89644 100116 89672
rect 63460 89632 63466 89644
rect 100110 89632 100116 89644
rect 100168 89632 100174 89684
rect 122190 89632 122196 89684
rect 122248 89672 122254 89684
rect 217686 89672 217692 89684
rect 122248 89644 217692 89672
rect 122248 89632 122254 89644
rect 217686 89632 217692 89644
rect 217744 89632 217750 89684
rect 220630 89632 220636 89684
rect 220688 89672 220694 89684
rect 245010 89672 245016 89684
rect 220688 89644 245016 89672
rect 220688 89632 220694 89644
rect 245010 89632 245016 89644
rect 245068 89632 245074 89684
rect 67266 89564 67272 89616
rect 67324 89604 67330 89616
rect 94682 89604 94688 89616
rect 67324 89576 94688 89604
rect 67324 89564 67330 89576
rect 94682 89564 94688 89576
rect 94740 89564 94746 89616
rect 192018 89564 192024 89616
rect 192076 89604 192082 89616
rect 199378 89604 199384 89616
rect 192076 89576 199384 89604
rect 192076 89564 192082 89576
rect 199378 89564 199384 89576
rect 199436 89564 199442 89616
rect 204438 89564 204444 89616
rect 204496 89604 204502 89616
rect 205726 89604 205732 89616
rect 204496 89576 205732 89604
rect 204496 89564 204502 89576
rect 205726 89564 205732 89576
rect 205784 89564 205790 89616
rect 213362 88952 213368 89004
rect 213420 88992 213426 89004
rect 235258 88992 235264 89004
rect 213420 88964 235264 88992
rect 213420 88952 213426 88964
rect 235258 88952 235264 88964
rect 235316 88952 235322 89004
rect 254578 88952 254584 89004
rect 254636 88992 254642 89004
rect 583018 88992 583024 89004
rect 254636 88964 583024 88992
rect 254636 88952 254642 88964
rect 583018 88952 583024 88964
rect 583076 88952 583082 89004
rect 67450 88272 67456 88324
rect 67508 88312 67514 88324
rect 100018 88312 100024 88324
rect 67508 88284 100024 88312
rect 67508 88272 67514 88284
rect 100018 88272 100024 88284
rect 100076 88272 100082 88324
rect 103514 88312 103520 88324
rect 103486 88272 103520 88312
rect 103572 88312 103578 88324
rect 214006 88312 214012 88324
rect 103572 88284 214012 88312
rect 103572 88272 103578 88284
rect 214006 88272 214012 88284
rect 214064 88272 214070 88324
rect 68922 88204 68928 88256
rect 68980 88244 68986 88256
rect 80698 88244 80704 88256
rect 68980 88216 80704 88244
rect 68980 88204 68986 88216
rect 80698 88204 80704 88216
rect 80756 88204 80762 88256
rect 86126 88204 86132 88256
rect 86184 88244 86190 88256
rect 103486 88244 103514 88272
rect 86184 88216 103514 88244
rect 86184 88204 86190 88216
rect 111886 88204 111892 88256
rect 111944 88244 111950 88256
rect 205542 88244 205548 88256
rect 111944 88216 205548 88244
rect 111944 88204 111950 88216
rect 205542 88204 205548 88216
rect 205600 88204 205606 88256
rect 207382 87592 207388 87644
rect 207440 87632 207446 87644
rect 246298 87632 246304 87644
rect 207440 87604 246304 87632
rect 207440 87592 207446 87604
rect 246298 87592 246304 87604
rect 246356 87592 246362 87644
rect 89806 86912 89812 86964
rect 89864 86952 89870 86964
rect 116670 86952 116676 86964
rect 89864 86924 116676 86952
rect 89864 86912 89870 86924
rect 116670 86912 116676 86924
rect 116728 86952 116734 86964
rect 218238 86952 218244 86964
rect 116728 86924 218244 86952
rect 116728 86912 116734 86924
rect 218238 86912 218244 86924
rect 218296 86912 218302 86964
rect 280246 86952 280252 86964
rect 277366 86924 280252 86952
rect 93302 86844 93308 86896
rect 93360 86884 93366 86896
rect 124858 86884 124864 86896
rect 93360 86856 124864 86884
rect 93360 86844 93366 86856
rect 124858 86844 124864 86856
rect 124916 86884 124922 86896
rect 125502 86884 125508 86896
rect 124916 86856 125508 86884
rect 124916 86844 124922 86856
rect 125502 86844 125508 86856
rect 125560 86844 125566 86896
rect 205726 86844 205732 86896
rect 205784 86884 205790 86896
rect 277366 86884 277394 86924
rect 280246 86912 280252 86924
rect 280304 86952 280310 86964
rect 580166 86952 580172 86964
rect 280304 86924 580172 86952
rect 280304 86912 280310 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 205784 86856 277394 86884
rect 205784 86844 205790 86856
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 53834 85524 53840 85536
rect 3568 85496 53840 85524
rect 3568 85484 3574 85496
rect 53834 85484 53840 85496
rect 53892 85484 53898 85536
rect 78398 85484 78404 85536
rect 78456 85524 78462 85536
rect 106918 85524 106924 85536
rect 78456 85496 106924 85524
rect 78456 85484 78462 85496
rect 106918 85484 106924 85496
rect 106976 85524 106982 85536
rect 204990 85524 204996 85536
rect 106976 85496 204996 85524
rect 106976 85484 106982 85496
rect 204990 85484 204996 85496
rect 205048 85484 205054 85536
rect 214558 85484 214564 85536
rect 214616 85524 214622 85536
rect 246482 85524 246488 85536
rect 214616 85496 246488 85524
rect 214616 85484 214622 85496
rect 246482 85484 246488 85496
rect 246540 85484 246546 85536
rect 198366 85416 198372 85468
rect 198424 85456 198430 85468
rect 262858 85456 262864 85468
rect 198424 85428 262864 85456
rect 198424 85416 198430 85428
rect 262858 85416 262864 85428
rect 262916 85416 262922 85468
rect 88334 84124 88340 84176
rect 88392 84164 88398 84176
rect 122190 84164 122196 84176
rect 88392 84136 122196 84164
rect 88392 84124 88398 84136
rect 122190 84124 122196 84136
rect 122248 84124 122254 84176
rect 169846 84124 169852 84176
rect 169904 84164 169910 84176
rect 171042 84164 171048 84176
rect 169904 84136 171048 84164
rect 169904 84124 169910 84136
rect 171042 84124 171048 84136
rect 171100 84164 171106 84176
rect 193398 84164 193404 84176
rect 171100 84136 193404 84164
rect 171100 84124 171106 84136
rect 193398 84124 193404 84136
rect 193456 84124 193462 84176
rect 74534 84056 74540 84108
rect 74592 84096 74598 84108
rect 101582 84096 101588 84108
rect 74592 84068 101588 84096
rect 74592 84056 74598 84068
rect 101582 84056 101588 84068
rect 101640 84056 101646 84108
rect 193398 83512 193404 83564
rect 193456 83552 193462 83564
rect 226978 83552 226984 83564
rect 193456 83524 226984 83552
rect 193456 83512 193462 83524
rect 226978 83512 226984 83524
rect 227036 83512 227042 83564
rect 193030 83444 193036 83496
rect 193088 83484 193094 83496
rect 259454 83484 259460 83496
rect 193088 83456 259460 83484
rect 193088 83444 193094 83456
rect 259454 83444 259460 83456
rect 259512 83444 259518 83496
rect 227070 82832 227076 82884
rect 227128 82872 227134 82884
rect 241514 82872 241520 82884
rect 227128 82844 241520 82872
rect 227128 82832 227134 82844
rect 241514 82832 241520 82844
rect 241572 82832 241578 82884
rect 77294 82764 77300 82816
rect 77352 82804 77358 82816
rect 108390 82804 108396 82816
rect 77352 82776 108396 82804
rect 77352 82764 77358 82776
rect 108390 82764 108396 82776
rect 108448 82764 108454 82816
rect 185578 82764 185584 82816
rect 185636 82804 185642 82816
rect 229094 82804 229100 82816
rect 185636 82776 229100 82804
rect 185636 82764 185642 82776
rect 229094 82764 229100 82776
rect 229152 82764 229158 82816
rect 75914 82696 75920 82748
rect 75972 82736 75978 82748
rect 94774 82736 94780 82748
rect 75972 82708 94780 82736
rect 75972 82696 75978 82708
rect 94774 82696 94780 82708
rect 94832 82736 94838 82748
rect 95142 82736 95148 82748
rect 94832 82708 95148 82736
rect 94832 82696 94838 82708
rect 95142 82696 95148 82708
rect 95200 82696 95206 82748
rect 186958 82696 186964 82748
rect 187016 82736 187022 82748
rect 200114 82736 200120 82748
rect 187016 82708 200120 82736
rect 187016 82696 187022 82708
rect 200114 82696 200120 82708
rect 200172 82736 200178 82748
rect 201402 82736 201408 82748
rect 200172 82708 201408 82736
rect 200172 82696 200178 82708
rect 201402 82696 201408 82708
rect 201460 82696 201466 82748
rect 201402 82084 201408 82136
rect 201460 82124 201466 82136
rect 214558 82124 214564 82136
rect 201460 82096 214564 82124
rect 201460 82084 201466 82096
rect 214558 82084 214564 82096
rect 214616 82084 214622 82136
rect 242158 82124 242164 82136
rect 219406 82096 242164 82124
rect 215386 81948 215392 82000
rect 215444 81988 215450 82000
rect 216030 81988 216036 82000
rect 215444 81960 216036 81988
rect 215444 81948 215450 81960
rect 216030 81948 216036 81960
rect 216088 81988 216094 82000
rect 219406 81988 219434 82096
rect 242158 82084 242164 82096
rect 242216 82084 242222 82136
rect 216088 81960 219434 81988
rect 216088 81948 216094 81960
rect 85758 81336 85764 81388
rect 85816 81376 85822 81388
rect 103606 81376 103612 81388
rect 85816 81348 103612 81376
rect 85816 81336 85822 81348
rect 103606 81336 103612 81348
rect 103664 81336 103670 81388
rect 109678 81336 109684 81388
rect 109736 81376 109742 81388
rect 224954 81376 224960 81388
rect 109736 81348 224960 81376
rect 109736 81336 109742 81348
rect 224954 81336 224960 81348
rect 225012 81336 225018 81388
rect 69198 81268 69204 81320
rect 69256 81308 69262 81320
rect 169846 81308 169852 81320
rect 69256 81280 169852 81308
rect 69256 81268 69262 81280
rect 169846 81268 169852 81280
rect 169904 81268 169910 81320
rect 201586 80656 201592 80708
rect 201644 80696 201650 80708
rect 253198 80696 253204 80708
rect 201644 80668 253204 80696
rect 201644 80656 201650 80668
rect 253198 80656 253204 80668
rect 253256 80656 253262 80708
rect 201586 80044 201592 80096
rect 201644 80084 201650 80096
rect 202138 80084 202144 80096
rect 201644 80056 202144 80084
rect 201644 80044 201650 80056
rect 202138 80044 202144 80056
rect 202196 80044 202202 80096
rect 54478 79976 54484 80028
rect 54536 80016 54542 80028
rect 55122 80016 55128 80028
rect 54536 79988 55128 80016
rect 54536 79976 54542 79988
rect 55122 79976 55128 79988
rect 55180 80016 55186 80028
rect 188522 80016 188528 80028
rect 55180 79988 188528 80016
rect 55180 79976 55186 79988
rect 188522 79976 188528 79988
rect 188580 79976 188586 80028
rect 66070 79908 66076 79960
rect 66128 79948 66134 79960
rect 112438 79948 112444 79960
rect 66128 79920 112444 79948
rect 66128 79908 66134 79920
rect 112438 79908 112444 79920
rect 112496 79908 112502 79960
rect 177482 79908 177488 79960
rect 177540 79948 177546 79960
rect 227070 79948 227076 79960
rect 177540 79920 227076 79948
rect 177540 79908 177546 79920
rect 227070 79908 227076 79920
rect 227128 79908 227134 79960
rect 191558 79296 191564 79348
rect 191616 79336 191622 79348
rect 280154 79336 280160 79348
rect 191616 79308 280160 79336
rect 191616 79296 191622 79308
rect 280154 79296 280160 79308
rect 280212 79296 280218 79348
rect 82814 78616 82820 78668
rect 82872 78656 82878 78668
rect 178034 78656 178040 78668
rect 82872 78628 178040 78656
rect 82872 78616 82878 78628
rect 178034 78616 178040 78628
rect 178092 78616 178098 78668
rect 186958 78616 186964 78668
rect 187016 78656 187022 78668
rect 190362 78656 190368 78668
rect 187016 78628 190368 78656
rect 187016 78616 187022 78628
rect 190362 78616 190368 78628
rect 190420 78656 190426 78668
rect 263594 78656 263600 78668
rect 190420 78628 263600 78656
rect 190420 78616 190426 78628
rect 263594 78616 263600 78628
rect 263652 78656 263658 78668
rect 264238 78656 264244 78668
rect 263652 78628 264244 78656
rect 263652 78616 263658 78628
rect 264238 78616 264244 78628
rect 264296 78616 264302 78668
rect 177390 78548 177396 78600
rect 177448 78588 177454 78600
rect 230566 78588 230572 78600
rect 177448 78560 230572 78588
rect 177448 78548 177454 78560
rect 230566 78548 230572 78560
rect 230624 78548 230630 78600
rect 85574 77936 85580 77988
rect 85632 77976 85638 77988
rect 105538 77976 105544 77988
rect 85632 77948 105544 77976
rect 85632 77936 85638 77948
rect 105538 77936 105544 77948
rect 105596 77936 105602 77988
rect 260098 77936 260104 77988
rect 260156 77976 260162 77988
rect 295334 77976 295340 77988
rect 260156 77948 295340 77976
rect 260156 77936 260162 77948
rect 295334 77936 295340 77948
rect 295392 77936 295398 77988
rect 65518 77188 65524 77240
rect 65576 77228 65582 77240
rect 102226 77228 102232 77240
rect 65576 77200 102232 77228
rect 65576 77188 65582 77200
rect 102226 77188 102232 77200
rect 102284 77188 102290 77240
rect 169018 77188 169024 77240
rect 169076 77228 169082 77240
rect 229186 77228 229192 77240
rect 169076 77200 229192 77228
rect 169076 77188 169082 77200
rect 229186 77188 229192 77200
rect 229244 77188 229250 77240
rect 80698 76508 80704 76560
rect 80756 76548 80762 76560
rect 100018 76548 100024 76560
rect 80756 76520 100024 76548
rect 80756 76508 80762 76520
rect 100018 76508 100024 76520
rect 100076 76508 100082 76560
rect 109034 76508 109040 76560
rect 109092 76548 109098 76560
rect 135990 76548 135996 76560
rect 109092 76520 135996 76548
rect 109092 76508 109098 76520
rect 135990 76508 135996 76520
rect 136048 76508 136054 76560
rect 193122 76508 193128 76560
rect 193180 76548 193186 76560
rect 338114 76548 338120 76560
rect 193180 76520 338120 76548
rect 193180 76508 193186 76520
rect 338114 76508 338120 76520
rect 338172 76508 338178 76560
rect 182818 75828 182824 75880
rect 182876 75868 182882 75880
rect 230474 75868 230480 75880
rect 182876 75840 230480 75868
rect 182876 75828 182882 75840
rect 230474 75828 230480 75840
rect 230532 75828 230538 75880
rect 67634 75148 67640 75200
rect 67692 75188 67698 75200
rect 171778 75188 171784 75200
rect 67692 75160 171784 75188
rect 67692 75148 67698 75160
rect 171778 75148 171784 75160
rect 171836 75148 171842 75200
rect 190178 75148 190184 75200
rect 190236 75188 190242 75200
rect 248414 75188 248420 75200
rect 190236 75160 248420 75188
rect 190236 75148 190242 75160
rect 248414 75148 248420 75160
rect 248472 75188 248478 75200
rect 249058 75188 249064 75200
rect 248472 75160 249064 75188
rect 248472 75148 248478 75160
rect 249058 75148 249064 75160
rect 249116 75148 249122 75200
rect 85666 74468 85672 74520
rect 85724 74508 85730 74520
rect 120074 74508 120080 74520
rect 85724 74480 120080 74508
rect 85724 74468 85730 74480
rect 120074 74468 120080 74480
rect 120132 74508 120138 74520
rect 213178 74508 213184 74520
rect 120132 74480 213184 74508
rect 120132 74468 120138 74480
rect 213178 74468 213184 74480
rect 213236 74468 213242 74520
rect 153930 74400 153936 74452
rect 153988 74440 153994 74452
rect 237374 74440 237380 74452
rect 153988 74412 237380 74440
rect 153988 74400 153994 74412
rect 237374 74400 237380 74412
rect 237432 74400 237438 74452
rect 237374 73176 237380 73228
rect 237432 73216 237438 73228
rect 238110 73216 238116 73228
rect 237432 73188 238116 73216
rect 237432 73176 237438 73188
rect 238110 73176 238116 73188
rect 238168 73176 238174 73228
rect 258718 73216 258724 73228
rect 258046 73188 258724 73216
rect 64782 73108 64788 73160
rect 64840 73148 64846 73160
rect 190178 73148 190184 73160
rect 64840 73120 190184 73148
rect 64840 73108 64846 73120
rect 190178 73108 190184 73120
rect 190236 73108 190242 73160
rect 207014 73108 207020 73160
rect 207072 73148 207078 73160
rect 258046 73148 258074 73188
rect 258718 73176 258724 73188
rect 258776 73176 258782 73228
rect 207072 73120 258074 73148
rect 207072 73108 207078 73120
rect 129642 73040 129648 73092
rect 129700 73080 129706 73092
rect 227898 73080 227904 73092
rect 129700 73052 227904 73080
rect 129700 73040 129706 73052
rect 227898 73040 227904 73052
rect 227956 73040 227962 73092
rect 227898 71748 227904 71800
rect 227956 71788 227962 71800
rect 228358 71788 228364 71800
rect 227956 71760 228364 71788
rect 227956 71748 227962 71760
rect 228358 71748 228364 71760
rect 228416 71748 228422 71800
rect 93118 71680 93124 71732
rect 93176 71720 93182 71732
rect 106274 71720 106280 71732
rect 93176 71692 106280 71720
rect 93176 71680 93182 71692
rect 106274 71680 106280 71692
rect 106332 71680 106338 71732
rect 166258 71680 166264 71732
rect 166316 71720 166322 71732
rect 231946 71720 231952 71732
rect 166316 71692 231952 71720
rect 166316 71680 166322 71692
rect 231946 71680 231952 71692
rect 232004 71680 232010 71732
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 95326 71652 95332 71664
rect 3568 71624 95332 71652
rect 3568 71612 3574 71624
rect 95326 71612 95332 71624
rect 95384 71612 95390 71664
rect 187602 71000 187608 71052
rect 187660 71040 187666 71052
rect 288434 71040 288440 71052
rect 187660 71012 288440 71040
rect 187660 71000 187666 71012
rect 288434 71000 288440 71012
rect 288492 71000 288498 71052
rect 67542 70320 67548 70372
rect 67600 70360 67606 70372
rect 180794 70360 180800 70372
rect 67600 70332 180800 70360
rect 67600 70320 67606 70332
rect 180794 70320 180800 70332
rect 180852 70360 180858 70372
rect 181438 70360 181444 70372
rect 180852 70332 181444 70360
rect 180852 70320 180858 70332
rect 181438 70320 181444 70332
rect 181496 70320 181502 70372
rect 160738 70252 160744 70304
rect 160796 70292 160802 70304
rect 244274 70292 244280 70304
rect 160796 70264 244280 70292
rect 160796 70252 160802 70264
rect 244274 70252 244280 70264
rect 244332 70252 244338 70304
rect 244274 69844 244280 69896
rect 244332 69884 244338 69896
rect 244918 69884 244924 69896
rect 244332 69856 244924 69884
rect 244332 69844 244338 69856
rect 244918 69844 244924 69856
rect 244976 69844 244982 69896
rect 222286 69028 222292 69080
rect 222344 69068 222350 69080
rect 339494 69068 339500 69080
rect 222344 69040 339500 69068
rect 222344 69028 222350 69040
rect 339494 69028 339500 69040
rect 339552 69028 339558 69080
rect 124858 68960 124864 69012
rect 124916 69000 124922 69012
rect 222194 69000 222200 69012
rect 124916 68972 222200 69000
rect 124916 68960 124922 68972
rect 222194 68960 222200 68972
rect 222252 69000 222258 69012
rect 222838 69000 222844 69012
rect 222252 68972 222844 69000
rect 222252 68960 222258 68972
rect 222838 68960 222844 68972
rect 222896 68960 222902 69012
rect 193306 68892 193312 68944
rect 193364 68932 193370 68944
rect 193858 68932 193864 68944
rect 193364 68904 193864 68932
rect 193364 68892 193370 68904
rect 193858 68892 193864 68904
rect 193916 68932 193922 68944
rect 281534 68932 281540 68944
rect 193916 68904 281540 68932
rect 193916 68892 193922 68904
rect 281534 68892 281540 68904
rect 281592 68892 281598 68944
rect 88334 68280 88340 68332
rect 88392 68320 88398 68332
rect 169754 68320 169760 68332
rect 88392 68292 169760 68320
rect 88392 68280 88398 68292
rect 169754 68280 169760 68292
rect 169812 68280 169818 68332
rect 97258 67532 97264 67584
rect 97316 67572 97322 67584
rect 227714 67572 227720 67584
rect 97316 67544 227720 67572
rect 97316 67532 97322 67544
rect 227714 67532 227720 67544
rect 227772 67532 227778 67584
rect 65518 66852 65524 66904
rect 65576 66892 65582 66904
rect 123478 66892 123484 66904
rect 65576 66864 123484 66892
rect 65576 66852 65582 66864
rect 123478 66852 123484 66864
rect 123536 66852 123542 66904
rect 190270 66852 190276 66904
rect 190328 66892 190334 66904
rect 320266 66892 320272 66904
rect 190328 66864 320272 66892
rect 190328 66852 190334 66864
rect 320266 66852 320272 66864
rect 320324 66852 320330 66904
rect 71866 66172 71872 66224
rect 71924 66212 71930 66224
rect 197998 66212 198004 66224
rect 71924 66184 198004 66212
rect 71924 66172 71930 66184
rect 197998 66172 198004 66184
rect 198056 66172 198062 66224
rect 200758 66172 200764 66224
rect 200816 66212 200822 66224
rect 201402 66212 201408 66224
rect 200816 66184 201408 66212
rect 200816 66172 200822 66184
rect 201402 66172 201408 66184
rect 201460 66212 201466 66224
rect 250438 66212 250444 66224
rect 201460 66184 250444 66212
rect 201460 66172 201466 66184
rect 250438 66172 250444 66184
rect 250496 66172 250502 66224
rect 100018 66104 100024 66156
rect 100076 66144 100082 66156
rect 207014 66144 207020 66156
rect 100076 66116 207020 66144
rect 100076 66104 100082 66116
rect 207014 66104 207020 66116
rect 207072 66104 207078 66156
rect 87046 64812 87052 64864
rect 87104 64852 87110 64864
rect 215294 64852 215300 64864
rect 87104 64824 215300 64852
rect 87104 64812 87110 64824
rect 215294 64812 215300 64824
rect 215352 64812 215358 64864
rect 80054 64744 80060 64796
rect 80112 64784 80118 64796
rect 205634 64784 205640 64796
rect 80112 64756 205640 64784
rect 80112 64744 80118 64756
rect 205634 64744 205640 64756
rect 205692 64744 205698 64796
rect 213178 64132 213184 64184
rect 213236 64172 213242 64184
rect 333974 64172 333980 64184
rect 213236 64144 333980 64172
rect 213236 64132 213242 64144
rect 333974 64132 333980 64144
rect 334032 64132 334038 64184
rect 205634 63520 205640 63572
rect 205692 63560 205698 63572
rect 206278 63560 206284 63572
rect 205692 63532 206284 63560
rect 205692 63520 205698 63532
rect 206278 63520 206284 63532
rect 206336 63520 206342 63572
rect 215294 63520 215300 63572
rect 215352 63560 215358 63572
rect 215938 63560 215944 63572
rect 215352 63532 215944 63560
rect 215352 63520 215358 63532
rect 215938 63520 215944 63532
rect 215996 63520 216002 63572
rect 67726 63452 67732 63504
rect 67784 63492 67790 63504
rect 193858 63492 193864 63504
rect 67784 63464 193864 63492
rect 67784 63452 67790 63464
rect 193858 63452 193864 63464
rect 193916 63452 193922 63504
rect 194778 62024 194784 62076
rect 194836 62064 194842 62076
rect 287146 62064 287152 62076
rect 194836 62036 287152 62064
rect 194836 62024 194842 62036
rect 287146 62024 287152 62036
rect 287204 62064 287210 62076
rect 288342 62064 288348 62076
rect 287204 62036 288348 62064
rect 287204 62024 287210 62036
rect 288342 62024 288348 62036
rect 288400 62024 288406 62076
rect 86954 61956 86960 62008
rect 87012 61996 87018 62008
rect 116026 61996 116032 62008
rect 87012 61968 116032 61996
rect 87012 61956 87018 61968
rect 116026 61956 116032 61968
rect 116084 61996 116090 62008
rect 216030 61996 216036 62008
rect 116084 61968 216036 61996
rect 116084 61956 116090 61968
rect 216030 61956 216036 61968
rect 216088 61956 216094 62008
rect 73798 61888 73804 61940
rect 73856 61928 73862 61940
rect 194686 61928 194692 61940
rect 73856 61900 194692 61928
rect 73856 61888 73862 61900
rect 194686 61888 194692 61900
rect 194744 61888 194750 61940
rect 288342 61344 288348 61396
rect 288400 61384 288406 61396
rect 345014 61384 345020 61396
rect 288400 61356 345020 61384
rect 288400 61344 288406 61356
rect 345014 61344 345020 61356
rect 345072 61344 345078 61396
rect 194686 60732 194692 60784
rect 194744 60772 194750 60784
rect 195238 60772 195244 60784
rect 194744 60744 195244 60772
rect 194744 60732 194750 60744
rect 195238 60732 195244 60744
rect 195296 60732 195302 60784
rect 69106 60664 69112 60716
rect 69164 60704 69170 60716
rect 194778 60704 194784 60716
rect 69164 60676 194784 60704
rect 69164 60664 69170 60676
rect 194778 60664 194784 60676
rect 194836 60664 194842 60716
rect 83458 60596 83464 60648
rect 83516 60636 83522 60648
rect 107654 60636 107660 60648
rect 83516 60608 107660 60636
rect 83516 60596 83522 60608
rect 107654 60596 107660 60608
rect 107712 60636 107718 60648
rect 209774 60636 209780 60648
rect 107712 60608 209780 60636
rect 107712 60596 107718 60608
rect 209774 60596 209780 60608
rect 209832 60636 209838 60648
rect 211062 60636 211068 60648
rect 209832 60608 211068 60636
rect 209832 60596 209838 60608
rect 211062 60596 211068 60608
rect 211120 60596 211126 60648
rect 240870 60052 240876 60104
rect 240928 60092 240934 60104
rect 278038 60092 278044 60104
rect 240928 60064 278044 60092
rect 240928 60052 240934 60064
rect 278038 60052 278044 60064
rect 278096 60052 278102 60104
rect 199378 59984 199384 60036
rect 199436 60024 199442 60036
rect 244274 60024 244280 60036
rect 199436 59996 244280 60024
rect 199436 59984 199442 59996
rect 244274 59984 244280 59996
rect 244332 59984 244338 60036
rect 84838 59304 84844 59356
rect 84896 59344 84902 59356
rect 211154 59344 211160 59356
rect 84896 59316 211160 59344
rect 84896 59304 84902 59316
rect 211154 59304 211160 59316
rect 211212 59344 211218 59356
rect 212442 59344 212448 59356
rect 211212 59316 212448 59344
rect 211212 59304 211218 59316
rect 212442 59304 212448 59316
rect 212500 59304 212506 59356
rect 70486 59236 70492 59288
rect 70544 59276 70550 59288
rect 195974 59276 195980 59288
rect 70544 59248 195980 59276
rect 70544 59236 70550 59248
rect 195974 59236 195980 59248
rect 196032 59276 196038 59288
rect 196618 59276 196624 59288
rect 196032 59248 196624 59276
rect 196032 59236 196038 59248
rect 196618 59236 196624 59248
rect 196676 59236 196682 59288
rect 198734 58624 198740 58676
rect 198792 58664 198798 58676
rect 240134 58664 240140 58676
rect 198792 58636 240140 58664
rect 198792 58624 198798 58636
rect 240134 58624 240140 58636
rect 240192 58624 240198 58676
rect 91002 57876 91008 57928
rect 91060 57916 91066 57928
rect 219526 57916 219532 57928
rect 91060 57888 219532 57916
rect 91060 57876 91066 57888
rect 219526 57876 219532 57888
rect 219584 57916 219590 57928
rect 220078 57916 220084 57928
rect 219584 57888 220084 57916
rect 219584 57876 219590 57888
rect 220078 57876 220084 57888
rect 220136 57876 220142 57928
rect 212442 57808 212448 57860
rect 212500 57848 212506 57860
rect 278682 57848 278688 57860
rect 212500 57820 278688 57848
rect 212500 57808 212506 57820
rect 278682 57808 278688 57820
rect 278740 57808 278746 57860
rect 278682 57196 278688 57248
rect 278740 57236 278746 57248
rect 353294 57236 353300 57248
rect 278740 57208 353300 57236
rect 278740 57196 278746 57208
rect 353294 57196 353300 57208
rect 353352 57196 353358 57248
rect 74626 56516 74632 56568
rect 74684 56556 74690 56568
rect 202138 56556 202144 56568
rect 74684 56528 202144 56556
rect 74684 56516 74690 56528
rect 202138 56516 202144 56528
rect 202196 56516 202202 56568
rect 211062 56516 211068 56568
rect 211120 56556 211126 56568
rect 296714 56556 296720 56568
rect 211120 56528 296720 56556
rect 211120 56516 211126 56528
rect 296714 56516 296720 56528
rect 296772 56556 296778 56568
rect 298002 56556 298008 56568
rect 296772 56528 298008 56556
rect 296772 56516 296778 56528
rect 298002 56516 298008 56528
rect 298060 56516 298066 56568
rect 298002 55836 298008 55888
rect 298060 55876 298066 55888
rect 322934 55876 322940 55888
rect 298060 55848 322940 55876
rect 298060 55836 298066 55848
rect 322934 55836 322940 55848
rect 322992 55836 322998 55888
rect 71774 54476 71780 54528
rect 71832 54516 71838 54528
rect 151170 54516 151176 54528
rect 71832 54488 151176 54516
rect 71832 54476 71838 54488
rect 151170 54476 151176 54488
rect 151228 54476 151234 54528
rect 206278 54476 206284 54528
rect 206336 54516 206342 54528
rect 232498 54516 232504 54528
rect 206336 54488 232504 54516
rect 206336 54476 206342 54488
rect 232498 54476 232504 54488
rect 232556 54476 232562 54528
rect 232590 54476 232596 54528
rect 232648 54516 232654 54528
rect 324406 54516 324412 54528
rect 232648 54488 324412 54516
rect 232648 54476 232654 54488
rect 324406 54476 324412 54488
rect 324464 54476 324470 54528
rect 86954 53048 86960 53100
rect 87012 53088 87018 53100
rect 153838 53088 153844 53100
rect 87012 53060 153844 53088
rect 87012 53048 87018 53060
rect 153838 53048 153844 53060
rect 153896 53048 153902 53100
rect 97258 51688 97264 51740
rect 97316 51728 97322 51740
rect 131758 51728 131764 51740
rect 97316 51700 131764 51728
rect 97316 51688 97322 51700
rect 131758 51688 131764 51700
rect 131816 51688 131822 51740
rect 183462 51688 183468 51740
rect 183520 51728 183526 51740
rect 281534 51728 281540 51740
rect 183520 51700 281540 51728
rect 183520 51688 183526 51700
rect 281534 51688 281540 51700
rect 281592 51688 281598 51740
rect 14 50328 20 50380
rect 72 50368 78 50380
rect 97350 50368 97356 50380
rect 72 50340 97356 50368
rect 72 50328 78 50340
rect 97350 50328 97356 50340
rect 97408 50328 97414 50380
rect 100754 50328 100760 50380
rect 100812 50368 100818 50380
rect 146938 50368 146944 50380
rect 100812 50340 146944 50368
rect 100812 50328 100818 50340
rect 146938 50328 146944 50340
rect 146996 50328 147002 50380
rect 169570 50328 169576 50380
rect 169628 50368 169634 50380
rect 335354 50368 335360 50380
rect 169628 50340 335360 50368
rect 169628 50328 169634 50340
rect 335354 50328 335360 50340
rect 335412 50328 335418 50380
rect 295978 49648 295984 49700
rect 296036 49688 296042 49700
rect 296714 49688 296720 49700
rect 296036 49660 296720 49688
rect 296036 49648 296042 49660
rect 296714 49648 296720 49660
rect 296772 49648 296778 49700
rect 107654 49036 107660 49088
rect 107712 49076 107718 49088
rect 126238 49076 126244 49088
rect 107712 49048 126244 49076
rect 107712 49036 107718 49048
rect 126238 49036 126244 49048
rect 126296 49036 126302 49088
rect 250530 49036 250536 49088
rect 250588 49076 250594 49088
rect 260834 49076 260840 49088
rect 250588 49048 260840 49076
rect 250588 49036 250594 49048
rect 260834 49036 260840 49048
rect 260892 49036 260898 49088
rect 52454 48968 52460 49020
rect 52512 49008 52518 49020
rect 133138 49008 133144 49020
rect 52512 48980 133144 49008
rect 52512 48968 52518 48980
rect 133138 48968 133144 48980
rect 133196 48968 133202 49020
rect 181438 48968 181444 49020
rect 181496 49008 181502 49020
rect 251266 49008 251272 49020
rect 181496 48980 251272 49008
rect 181496 48968 181502 48980
rect 251266 48968 251272 48980
rect 251324 48968 251330 49020
rect 2866 47540 2872 47592
rect 2924 47580 2930 47592
rect 147030 47580 147036 47592
rect 2924 47552 147036 47580
rect 2924 47540 2930 47552
rect 147030 47540 147036 47552
rect 147088 47540 147094 47592
rect 188430 46860 188436 46912
rect 188488 46900 188494 46912
rect 580166 46900 580172 46912
rect 188488 46872 580172 46900
rect 188488 46860 188494 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 46180 3516 46232
rect 3568 46220 3574 46232
rect 54478 46220 54484 46232
rect 3568 46192 54484 46220
rect 3568 46180 3574 46192
rect 54478 46180 54484 46192
rect 54536 46180 54542 46232
rect 78674 46180 78680 46232
rect 78732 46220 78738 46232
rect 142890 46220 142896 46232
rect 78732 46192 142896 46220
rect 78732 46180 78738 46192
rect 142890 46180 142896 46192
rect 142948 46180 142954 46232
rect 186130 43392 186136 43444
rect 186188 43432 186194 43444
rect 249794 43432 249800 43444
rect 186188 43404 249800 43432
rect 186188 43392 186194 43404
rect 249794 43392 249800 43404
rect 249852 43392 249858 43444
rect 75914 42032 75920 42084
rect 75972 42072 75978 42084
rect 137278 42072 137284 42084
rect 75972 42044 137284 42072
rect 75972 42032 75978 42044
rect 137278 42032 137284 42044
rect 137336 42032 137342 42084
rect 184750 42032 184756 42084
rect 184808 42072 184814 42084
rect 298094 42072 298100 42084
rect 184808 42044 298100 42072
rect 184808 42032 184814 42044
rect 298094 42032 298100 42044
rect 298152 42032 298158 42084
rect 45554 40672 45560 40724
rect 45612 40712 45618 40724
rect 156598 40712 156604 40724
rect 45612 40684 156604 40712
rect 45612 40672 45618 40684
rect 156598 40672 156604 40684
rect 156656 40672 156662 40724
rect 27706 39312 27712 39364
rect 27764 39352 27770 39364
rect 159358 39352 159364 39364
rect 27764 39324 159364 39352
rect 27764 39312 27770 39324
rect 159358 39312 159364 39324
rect 159416 39312 159422 39364
rect 179230 39312 179236 39364
rect 179288 39352 179294 39364
rect 309134 39352 309140 39364
rect 179288 39324 309140 39352
rect 179288 39312 179294 39324
rect 309134 39312 309140 39324
rect 309192 39312 309198 39364
rect 84194 37952 84200 38004
rect 84252 37992 84258 38004
rect 122098 37992 122104 38004
rect 84252 37964 122104 37992
rect 84252 37952 84258 37964
rect 122098 37952 122104 37964
rect 122156 37952 122162 38004
rect 113174 37884 113180 37936
rect 113232 37924 113238 37936
rect 160094 37924 160100 37936
rect 113232 37896 160100 37924
rect 113232 37884 113238 37896
rect 160094 37884 160100 37896
rect 160152 37884 160158 37936
rect 208394 37884 208400 37936
rect 208452 37924 208458 37936
rect 278774 37924 278780 37936
rect 208452 37896 278780 37924
rect 208452 37884 208458 37896
rect 278774 37884 278780 37896
rect 278832 37884 278838 37936
rect 73154 36524 73160 36576
rect 73212 36564 73218 36576
rect 155310 36564 155316 36576
rect 73212 36536 155316 36564
rect 73212 36524 73218 36536
rect 155310 36524 155316 36536
rect 155368 36524 155374 36576
rect 82814 35164 82820 35216
rect 82872 35204 82878 35216
rect 145558 35204 145564 35216
rect 82872 35176 145564 35204
rect 82872 35164 82878 35176
rect 145558 35164 145564 35176
rect 145616 35164 145622 35216
rect 60734 33736 60740 33788
rect 60792 33776 60798 33788
rect 174538 33776 174544 33788
rect 60792 33748 174544 33776
rect 60792 33736 60798 33748
rect 174538 33736 174544 33748
rect 174596 33736 174602 33788
rect 195238 33736 195244 33788
rect 195296 33776 195302 33788
rect 311894 33776 311900 33788
rect 195296 33748 311900 33776
rect 195296 33736 195302 33748
rect 311894 33736 311900 33748
rect 311952 33736 311958 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 53098 33096 53104 33108
rect 3568 33068 53104 33096
rect 3568 33056 3574 33068
rect 53098 33056 53104 33068
rect 53156 33056 53162 33108
rect 61746 32376 61752 32428
rect 61804 32416 61810 32428
rect 125594 32416 125600 32428
rect 61804 32388 125600 32416
rect 61804 32376 61810 32388
rect 125594 32376 125600 32388
rect 125652 32376 125658 32428
rect 233878 32376 233884 32428
rect 233936 32416 233942 32428
rect 316034 32416 316040 32428
rect 233936 32388 316040 32416
rect 233936 32376 233942 32388
rect 316034 32376 316040 32388
rect 316092 32376 316098 32428
rect 120074 29656 120080 29708
rect 120132 29696 120138 29708
rect 157978 29696 157984 29708
rect 120132 29668 157984 29696
rect 120132 29656 120138 29668
rect 157978 29656 157984 29668
rect 158036 29656 158042 29708
rect 59354 29588 59360 29640
rect 59412 29628 59418 29640
rect 130470 29628 130476 29640
rect 59412 29600 130476 29628
rect 59412 29588 59418 29600
rect 130470 29588 130476 29600
rect 130528 29588 130534 29640
rect 215938 29588 215944 29640
rect 215996 29628 216002 29640
rect 266354 29628 266360 29640
rect 215996 29600 266360 29628
rect 215996 29588 216002 29600
rect 266354 29588 266360 29600
rect 266412 29588 266418 29640
rect 106274 28228 106280 28280
rect 106332 28268 106338 28280
rect 162118 28268 162124 28280
rect 106332 28240 162124 28268
rect 106332 28228 106338 28240
rect 162118 28228 162124 28240
rect 162176 28228 162182 28280
rect 193858 28228 193864 28280
rect 193916 28268 193922 28280
rect 291194 28268 291200 28280
rect 193916 28240 291200 28268
rect 193916 28228 193922 28240
rect 291194 28228 291200 28240
rect 291252 28228 291258 28280
rect 191650 26868 191656 26920
rect 191708 26908 191714 26920
rect 322198 26908 322204 26920
rect 191708 26880 322204 26908
rect 191708 26868 191714 26880
rect 322198 26868 322204 26880
rect 322256 26868 322262 26920
rect 69106 25508 69112 25560
rect 69164 25548 69170 25560
rect 152550 25548 152556 25560
rect 69164 25520 152556 25548
rect 69164 25508 69170 25520
rect 152550 25508 152556 25520
rect 152608 25508 152614 25560
rect 81434 24080 81440 24132
rect 81492 24120 81498 24132
rect 164234 24120 164240 24132
rect 81492 24092 164240 24120
rect 81492 24080 81498 24092
rect 164234 24080 164240 24092
rect 164292 24080 164298 24132
rect 235258 24080 235264 24132
rect 235316 24120 235322 24132
rect 287054 24120 287060 24132
rect 235316 24092 287060 24120
rect 235316 24080 235322 24092
rect 287054 24080 287060 24092
rect 287112 24080 287118 24132
rect 52546 22720 52552 22772
rect 52604 22760 52610 22772
rect 161474 22760 161480 22772
rect 52604 22732 161480 22760
rect 52604 22720 52610 22732
rect 161474 22720 161480 22732
rect 161532 22720 161538 22772
rect 89714 21360 89720 21412
rect 89772 21400 89778 21412
rect 148318 21400 148324 21412
rect 89772 21372 148324 21400
rect 89772 21360 89778 21372
rect 148318 21360 148324 21372
rect 148376 21360 148382 21412
rect 242158 21360 242164 21412
rect 242216 21400 242222 21412
rect 284386 21400 284392 21412
rect 242216 21372 284392 21400
rect 242216 21360 242222 21372
rect 284386 21360 284392 21372
rect 284444 21360 284450 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 90358 20652 90364 20664
rect 3476 20624 90364 20652
rect 3476 20612 3482 20624
rect 90358 20612 90364 20624
rect 90416 20612 90422 20664
rect 95234 19932 95240 19984
rect 95292 19972 95298 19984
rect 151078 19972 151084 19984
rect 95292 19944 151084 19972
rect 95292 19932 95298 19944
rect 151078 19932 151084 19944
rect 151136 19932 151142 19984
rect 222838 19932 222844 19984
rect 222896 19972 222902 19984
rect 302326 19972 302332 19984
rect 222896 19944 302332 19972
rect 222896 19932 222902 19944
rect 302326 19932 302332 19944
rect 302384 19932 302390 19984
rect 240778 18640 240784 18692
rect 240836 18680 240842 18692
rect 276106 18680 276112 18692
rect 240836 18652 276112 18680
rect 240836 18640 240842 18652
rect 276106 18640 276112 18652
rect 276164 18640 276170 18692
rect 77294 18572 77300 18624
rect 77352 18612 77358 18624
rect 155218 18612 155224 18624
rect 77352 18584 155224 18612
rect 77352 18572 77358 18584
rect 155218 18572 155224 18584
rect 155276 18572 155282 18624
rect 180150 18572 180156 18624
rect 180208 18612 180214 18624
rect 242986 18612 242992 18624
rect 180208 18584 242992 18612
rect 180208 18572 180214 18584
rect 242986 18572 242992 18584
rect 243044 18572 243050 18624
rect 63494 17212 63500 17264
rect 63552 17252 63558 17264
rect 177298 17252 177304 17264
rect 63552 17224 177304 17252
rect 63552 17212 63558 17224
rect 177298 17212 177304 17224
rect 177356 17212 177362 17264
rect 238018 17212 238024 17264
rect 238076 17252 238082 17264
rect 269758 17252 269764 17264
rect 238076 17224 269764 17252
rect 238076 17212 238082 17224
rect 269758 17212 269764 17224
rect 269816 17212 269822 17264
rect 244918 15852 244924 15904
rect 244976 15892 244982 15904
rect 256694 15892 256700 15904
rect 244976 15864 256700 15892
rect 244976 15852 244982 15864
rect 256694 15852 256700 15864
rect 256752 15852 256758 15904
rect 270402 15852 270408 15904
rect 270460 15892 270466 15904
rect 330386 15892 330392 15904
rect 270460 15864 330392 15892
rect 270460 15852 270466 15864
rect 330386 15852 330392 15864
rect 330444 15852 330450 15904
rect 93118 14424 93124 14476
rect 93176 14464 93182 14476
rect 137370 14464 137376 14476
rect 93176 14436 137376 14464
rect 93176 14424 93182 14436
rect 137370 14424 137376 14436
rect 137428 14424 137434 14476
rect 253198 14424 253204 14476
rect 253256 14464 253262 14476
rect 321554 14464 321560 14476
rect 253256 14436 321560 14464
rect 253256 14424 253262 14436
rect 321554 14424 321560 14436
rect 321612 14424 321618 14476
rect 102226 13132 102232 13184
rect 102284 13172 102290 13184
rect 159450 13172 159456 13184
rect 102284 13144 159456 13172
rect 102284 13132 102290 13144
rect 159450 13132 159456 13144
rect 159508 13132 159514 13184
rect 61562 13064 61568 13116
rect 61620 13104 61626 13116
rect 140038 13104 140044 13116
rect 61620 13076 140044 13104
rect 61620 13064 61626 13076
rect 140038 13064 140044 13076
rect 140096 13064 140102 13116
rect 201402 13064 201408 13116
rect 201460 13104 201466 13116
rect 340966 13104 340972 13116
rect 201460 13076 340972 13104
rect 201460 13064 201466 13076
rect 340966 13064 340972 13076
rect 341024 13064 341030 13116
rect 75178 11704 75184 11756
rect 75236 11744 75242 11756
rect 135898 11744 135904 11756
rect 75236 11716 135904 11744
rect 75236 11704 75242 11716
rect 135898 11704 135904 11716
rect 135956 11704 135962 11756
rect 246390 11704 246396 11756
rect 246448 11744 246454 11756
rect 291930 11744 291936 11756
rect 246448 11716 291936 11744
rect 246448 11704 246454 11716
rect 291930 11704 291936 11716
rect 291988 11704 291994 11756
rect 58434 10276 58440 10328
rect 58492 10316 58498 10328
rect 138658 10316 138664 10328
rect 58492 10288 138664 10316
rect 58492 10276 58498 10288
rect 138658 10276 138664 10288
rect 138716 10276 138722 10328
rect 197998 10276 198004 10328
rect 198056 10316 198062 10328
rect 342898 10316 342904 10328
rect 198056 10288 342904 10316
rect 198056 10276 198062 10288
rect 342898 10276 342904 10288
rect 342956 10276 342962 10328
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 184198 8956 184204 8968
rect 10008 8928 184204 8956
rect 10008 8916 10014 8928
rect 184198 8916 184204 8928
rect 184256 8916 184262 8968
rect 196618 8916 196624 8968
rect 196676 8956 196682 8968
rect 258258 8956 258264 8968
rect 196676 8928 258264 8956
rect 196676 8916 196682 8928
rect 258258 8916 258264 8928
rect 258316 8916 258322 8968
rect 258718 8916 258724 8968
rect 258776 8956 258782 8968
rect 274818 8956 274824 8968
rect 258776 8928 274824 8956
rect 258776 8916 258782 8928
rect 274818 8916 274824 8928
rect 274876 8916 274882 8968
rect 97442 7624 97448 7676
rect 97500 7664 97506 7676
rect 141418 7664 141424 7676
rect 97500 7636 141424 7664
rect 97500 7624 97506 7636
rect 141418 7624 141424 7636
rect 141476 7624 141482 7676
rect 44266 7556 44272 7608
rect 44324 7596 44330 7608
rect 97258 7596 97264 7608
rect 44324 7568 97264 7596
rect 44324 7556 44330 7568
rect 97258 7556 97264 7568
rect 97316 7556 97322 7608
rect 220078 7556 220084 7608
rect 220136 7596 220142 7608
rect 346394 7596 346400 7608
rect 220136 7568 346400 7596
rect 220136 7556 220142 7568
rect 346394 7556 346400 7568
rect 346452 7556 346458 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 7558 6848 7564 6860
rect 3476 6820 7564 6848
rect 3476 6808 3482 6820
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 191742 6128 191748 6180
rect 191800 6168 191806 6180
rect 293678 6168 293684 6180
rect 191800 6140 293684 6168
rect 191800 6128 191806 6140
rect 293678 6128 293684 6140
rect 293736 6128 293742 6180
rect 305638 5516 305644 5568
rect 305696 5556 305702 5568
rect 309042 5556 309048 5568
rect 305696 5528 309048 5556
rect 305696 5516 305702 5528
rect 309042 5516 309048 5528
rect 309100 5516 309106 5568
rect 349798 5516 349804 5568
rect 349856 5556 349862 5568
rect 350534 5556 350540 5568
rect 349856 5528 350540 5556
rect 349856 5516 349862 5528
rect 350534 5516 350540 5528
rect 350592 5516 350598 5568
rect 323578 4904 323584 4956
rect 323636 4944 323642 4956
rect 326798 4944 326804 4956
rect 323636 4916 326804 4944
rect 323636 4904 323642 4916
rect 326798 4904 326804 4916
rect 326856 4904 326862 4956
rect 238110 4836 238116 4888
rect 238168 4876 238174 4888
rect 239306 4876 239312 4888
rect 238168 4848 239312 4876
rect 238168 4836 238174 4848
rect 239306 4836 239312 4848
rect 239364 4836 239370 4888
rect 65518 4768 65524 4820
rect 65576 4808 65582 4820
rect 149698 4808 149704 4820
rect 65576 4780 149704 4808
rect 65576 4768 65582 4780
rect 149698 4768 149704 4780
rect 149756 4768 149762 4820
rect 228358 4768 228364 4820
rect 228416 4808 228422 4820
rect 278314 4808 278320 4820
rect 228416 4780 278320 4808
rect 228416 4768 228422 4780
rect 278314 4768 278320 4780
rect 278372 4768 278378 4820
rect 342990 4768 342996 4820
rect 343048 4808 343054 4820
rect 346946 4808 346952 4820
rect 343048 4780 346952 4808
rect 343048 4768 343054 4780
rect 346946 4768 346952 4780
rect 347004 4768 347010 4820
rect 134518 4156 134524 4208
rect 134576 4196 134582 4208
rect 136450 4196 136456 4208
rect 134576 4168 136456 4196
rect 134576 4156 134582 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 309778 4156 309784 4208
rect 309836 4196 309842 4208
rect 315022 4196 315028 4208
rect 309836 4168 315028 4196
rect 309836 4156 309842 4168
rect 315022 4156 315028 4168
rect 315080 4156 315086 4208
rect 317322 4156 317328 4208
rect 317380 4196 317386 4208
rect 321646 4196 321652 4208
rect 317380 4168 321652 4196
rect 317380 4156 317386 4168
rect 321646 4156 321652 4168
rect 321704 4156 321710 4208
rect 337470 4156 337476 4208
rect 337528 4196 337534 4208
rect 340874 4196 340880 4208
rect 337528 4168 340880 4196
rect 337528 4156 337534 4168
rect 340874 4156 340880 4168
rect 340932 4156 340938 4208
rect 63218 4088 63224 4140
rect 63276 4128 63282 4140
rect 65426 4128 65432 4140
rect 63276 4100 65432 4128
rect 63276 4088 63282 4100
rect 65426 4088 65432 4100
rect 65484 4088 65490 4140
rect 266998 4088 267004 4140
rect 267056 4128 267062 4140
rect 267734 4128 267740 4140
rect 267056 4100 267740 4128
rect 267056 4088 267062 4100
rect 267734 4088 267740 4100
rect 267792 4088 267798 4140
rect 333882 4088 333888 4140
rect 333940 4128 333946 4140
rect 335446 4128 335452 4140
rect 333940 4100 335452 4128
rect 333940 4088 333946 4100
rect 335446 4088 335452 4100
rect 335504 4088 335510 4140
rect 150618 3612 150624 3664
rect 150676 3652 150682 3664
rect 152458 3652 152464 3664
rect 150676 3624 152464 3652
rect 150676 3612 150682 3624
rect 152458 3612 152464 3624
rect 152516 3612 152522 3664
rect 148502 3584 148508 3596
rect 142126 3556 148508 3584
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 4062 3516 4068 3528
rect 2832 3488 4068 3516
rect 2832 3476 2838 3488
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 12342 3516 12348 3528
rect 11112 3488 12348 3516
rect 11112 3476 11118 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 37182 3476 37188 3528
rect 37240 3516 37246 3528
rect 47578 3516 47584 3528
rect 37240 3488 47584 3516
rect 37240 3476 37246 3488
rect 47578 3476 47584 3488
rect 47636 3476 47642 3528
rect 69014 3476 69020 3528
rect 69072 3516 69078 3528
rect 70302 3516 70308 3528
rect 69072 3488 70308 3516
rect 69072 3476 69078 3488
rect 70302 3476 70308 3488
rect 70360 3476 70366 3528
rect 77386 3476 77392 3528
rect 77444 3516 77450 3528
rect 79318 3516 79324 3528
rect 77444 3488 79324 3516
rect 77444 3476 77450 3488
rect 79318 3476 79324 3488
rect 79376 3476 79382 3528
rect 85574 3476 85580 3528
rect 85632 3516 85638 3528
rect 86862 3516 86868 3528
rect 85632 3488 86868 3516
rect 85632 3476 85638 3488
rect 86862 3476 86868 3488
rect 86920 3476 86926 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 98638 3516 98644 3528
rect 91612 3488 98644 3516
rect 91612 3476 91618 3488
rect 98638 3476 98644 3488
rect 98696 3476 98702 3528
rect 102134 3476 102140 3528
rect 102192 3516 102198 3528
rect 103330 3516 103336 3528
rect 102192 3488 103336 3516
rect 102192 3476 102198 3488
rect 103330 3476 103336 3488
rect 103388 3476 103394 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 142126 3516 142154 3556
rect 148502 3544 148508 3556
rect 148560 3544 148566 3596
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 252370 3584 252376 3596
rect 251232 3556 252376 3584
rect 251232 3544 251238 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277118 3584 277124 3596
rect 276072 3556 277124 3584
rect 276072 3544 276078 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 140096 3488 142154 3516
rect 140096 3476 140102 3488
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 232498 3476 232504 3528
rect 232556 3516 232562 3528
rect 242894 3516 242900 3528
rect 232556 3488 242900 3516
rect 232556 3476 232562 3488
rect 242894 3476 242900 3488
rect 242952 3476 242958 3528
rect 287698 3476 287704 3528
rect 287756 3516 287762 3528
rect 290182 3516 290188 3528
rect 287756 3488 290188 3516
rect 287756 3476 287762 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 291930 3476 291936 3528
rect 291988 3516 291994 3528
rect 294874 3516 294880 3528
rect 291988 3488 294880 3516
rect 291988 3476 291994 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 300762 3516 300768 3528
rect 299532 3488 300768 3516
rect 299532 3476 299538 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 309134 3476 309140 3528
rect 309192 3516 309198 3528
rect 310238 3516 310244 3528
rect 309192 3488 310244 3516
rect 309192 3476 309198 3488
rect 310238 3476 310244 3488
rect 310296 3476 310302 3528
rect 319714 3476 319720 3528
rect 319772 3516 319778 3528
rect 320174 3516 320180 3528
rect 319772 3488 320180 3516
rect 319772 3476 319778 3488
rect 320174 3476 320180 3488
rect 320232 3476 320238 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 36538 3448 36544 3460
rect 20680 3420 36544 3448
rect 20680 3408 20686 3420
rect 36538 3408 36544 3420
rect 36596 3408 36602 3460
rect 51350 3408 51356 3460
rect 51408 3448 51414 3460
rect 75178 3448 75184 3460
rect 51408 3420 75184 3448
rect 51408 3408 51414 3420
rect 75178 3408 75184 3420
rect 75236 3408 75242 3460
rect 80882 3408 80888 3460
rect 80940 3448 80946 3460
rect 93118 3448 93124 3460
rect 80940 3420 93124 3448
rect 80940 3408 80946 3420
rect 93118 3408 93124 3420
rect 93176 3408 93182 3460
rect 99834 3408 99840 3460
rect 99892 3448 99898 3460
rect 108298 3448 108304 3460
rect 99892 3420 108304 3448
rect 99892 3408 99898 3420
rect 108298 3408 108304 3420
rect 108356 3408 108362 3460
rect 142798 3448 142804 3460
rect 113146 3420 142804 3448
rect 104526 3340 104532 3392
rect 104584 3380 104590 3392
rect 113146 3380 113174 3420
rect 142798 3408 142804 3420
rect 142856 3408 142862 3460
rect 214558 3408 214564 3460
rect 214616 3448 214622 3460
rect 246390 3448 246396 3460
rect 214616 3420 246396 3448
rect 214616 3408 214622 3420
rect 246390 3408 246396 3420
rect 246448 3408 246454 3460
rect 298738 3408 298744 3460
rect 298796 3448 298802 3460
rect 305546 3448 305552 3460
rect 298796 3420 305552 3448
rect 298796 3408 298802 3420
rect 305546 3408 305552 3420
rect 305604 3408 305610 3460
rect 322198 3408 322204 3460
rect 322256 3448 322262 3460
rect 329190 3448 329196 3460
rect 322256 3420 329196 3448
rect 322256 3408 322262 3420
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 334710 3408 334716 3460
rect 334768 3448 334774 3460
rect 344554 3448 344560 3460
rect 334768 3420 344560 3448
rect 334768 3408 334774 3420
rect 344554 3408 344560 3420
rect 344612 3408 344618 3460
rect 104584 3352 113174 3380
rect 104584 3340 104590 3352
rect 278038 3340 278044 3392
rect 278096 3380 278102 3392
rect 283098 3380 283104 3392
rect 278096 3352 283104 3380
rect 278096 3340 278102 3352
rect 283098 3340 283104 3352
rect 283156 3340 283162 3392
rect 346394 3340 346400 3392
rect 346452 3380 346458 3392
rect 349246 3380 349252 3392
rect 346452 3352 349252 3380
rect 346452 3340 346458 3352
rect 349246 3340 349252 3352
rect 349304 3340 349310 3392
rect 260650 3272 260656 3324
rect 260708 3312 260714 3324
rect 262306 3312 262312 3324
rect 260708 3284 262312 3312
rect 260708 3272 260714 3284
rect 262306 3272 262312 3284
rect 262364 3272 262370 3324
rect 327718 3272 327724 3324
rect 327776 3312 327782 3324
rect 332686 3312 332692 3324
rect 327776 3284 332692 3312
rect 327776 3272 327782 3284
rect 332686 3272 332692 3284
rect 332744 3272 332750 3324
rect 338758 3272 338764 3324
rect 338816 3312 338822 3324
rect 342162 3312 342168 3324
rect 338816 3284 342168 3312
rect 338816 3272 338822 3284
rect 342162 3272 342168 3284
rect 342220 3272 342226 3324
rect 348050 3272 348056 3324
rect 348108 3312 348114 3324
rect 351914 3312 351920 3324
rect 348108 3284 351920 3312
rect 348108 3272 348114 3284
rect 351914 3272 351920 3284
rect 351972 3272 351978 3324
rect 580994 3272 581000 3324
rect 581052 3312 581058 3324
rect 582558 3312 582564 3324
rect 581052 3284 582564 3312
rect 581052 3272 581058 3284
rect 582558 3272 582564 3284
rect 582616 3272 582622 3324
rect 269758 3068 269764 3120
rect 269816 3108 269822 3120
rect 272426 3108 272432 3120
rect 269816 3080 272432 3108
rect 269816 3068 269822 3080
rect 272426 3068 272432 3080
rect 272484 3068 272490 3120
rect 299658 3068 299664 3120
rect 299716 3108 299722 3120
rect 302234 3108 302240 3120
rect 299716 3080 302240 3108
rect 299716 3068 299722 3080
rect 302234 3068 302240 3080
rect 302292 3068 302298 3120
rect 246298 2932 246304 2984
rect 246356 2972 246362 2984
rect 247586 2972 247592 2984
rect 246356 2944 247592 2972
rect 246356 2932 246362 2944
rect 247586 2932 247592 2944
rect 247644 2932 247650 2984
rect 289078 2932 289084 2984
rect 289136 2972 289142 2984
rect 292574 2972 292580 2984
rect 289136 2944 292580 2972
rect 289136 2932 289142 2944
rect 292574 2932 292580 2944
rect 292632 2932 292638 2984
rect 307018 2932 307024 2984
rect 307076 2972 307082 2984
rect 307938 2972 307944 2984
rect 307076 2944 307944 2972
rect 307076 2932 307082 2944
rect 307938 2932 307944 2944
rect 307996 2932 308002 2984
rect 351638 2864 351644 2916
rect 351696 2904 351702 2916
rect 353294 2904 353300 2916
rect 351696 2876 353300 2904
rect 351696 2864 351702 2876
rect 353294 2864 353300 2876
rect 353352 2864 353358 2916
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 22738 2088 22744 2100
rect 7708 2060 22744 2088
rect 7708 2048 7714 2060
rect 22738 2048 22744 2060
rect 22796 2048 22802 2100
rect 93946 2048 93952 2100
rect 94004 2088 94010 2100
rect 130378 2088 130384 2100
rect 94004 2060 130384 2088
rect 94004 2048 94010 2060
rect 130378 2048 130384 2060
rect 130436 2048 130442 2100
<< via1 >>
rect 242808 703128 242860 703180
rect 348792 703128 348844 703180
rect 268384 703060 268436 703112
rect 413652 703060 413704 703112
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 218980 702992 219032 703044
rect 269120 702992 269172 703044
rect 280804 702992 280856 703044
rect 429844 702992 429896 703044
rect 179328 702924 179380 702976
rect 332508 702924 332560 702976
rect 188344 702856 188396 702908
rect 235172 702856 235224 702908
rect 249708 702856 249760 702908
rect 494796 702856 494848 702908
rect 154120 702788 154172 702840
rect 233240 702788 233292 702840
rect 285588 702788 285640 702840
rect 462320 702788 462372 702840
rect 187608 702720 187660 702772
rect 364984 702720 365036 702772
rect 205640 702652 205692 702704
rect 397368 702652 397420 702704
rect 24308 702584 24360 702636
rect 85580 702584 85632 702636
rect 137836 702584 137888 702636
rect 215300 702584 215352 702636
rect 222844 702584 222896 702636
rect 478512 702584 478564 702636
rect 67640 702516 67692 702568
rect 170312 702516 170364 702568
rect 224224 702516 224276 702568
rect 255964 702516 256016 702568
rect 543464 702516 543516 702568
rect 8116 702448 8168 702500
rect 96620 702448 96672 702500
rect 166356 702448 166408 702500
rect 527180 702448 527232 702500
rect 71044 700272 71096 700324
rect 105452 700272 105504 700324
rect 251824 700272 251876 700324
rect 283840 700272 283892 700324
rect 559656 700272 559708 700324
rect 582840 700272 582892 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 3424 683136 3476 683188
rect 33784 683136 33836 683188
rect 3516 670692 3568 670744
rect 15844 670692 15896 670744
rect 3424 656888 3476 656940
rect 74540 656888 74592 656940
rect 81440 620984 81492 621036
rect 201500 620984 201552 621036
rect 202144 620984 202196 621036
rect 3516 618264 3568 618316
rect 57244 618264 57296 618316
rect 164148 618264 164200 618316
rect 226340 618264 226392 618316
rect 161388 616836 161440 616888
rect 242900 616836 242952 616888
rect 233240 615952 233292 616004
rect 233884 615952 233936 616004
rect 167644 615544 167696 615596
rect 233240 615544 233292 615596
rect 155592 615476 155644 615528
rect 231860 615476 231912 615528
rect 147588 614184 147640 614236
rect 215944 614184 215996 614236
rect 173808 614116 173860 614168
rect 251916 614116 251968 614168
rect 166264 612824 166316 612876
rect 237472 612824 237524 612876
rect 184296 612756 184348 612808
rect 259460 612756 259512 612808
rect 152556 611396 152608 611448
rect 213184 611396 213236 611448
rect 66168 611328 66220 611380
rect 254124 611328 254176 611380
rect 137928 610036 137980 610088
rect 213092 610036 213144 610088
rect 160744 609968 160796 610020
rect 255320 609968 255372 610020
rect 202144 609288 202196 609340
rect 223028 609288 223080 609340
rect 219348 609220 219400 609272
rect 582840 609220 582892 609272
rect 140688 608608 140740 608660
rect 205732 608608 205784 608660
rect 182824 607248 182876 607300
rect 217692 607248 217744 607300
rect 177304 607180 177356 607232
rect 216956 607180 217008 607232
rect 218796 607180 218848 607232
rect 278044 607180 278096 607232
rect 215944 607112 215996 607164
rect 582380 607112 582432 607164
rect 176568 605888 176620 605940
rect 212540 605888 212592 605940
rect 3516 605820 3568 605872
rect 94688 605820 94740 605872
rect 98644 605820 98696 605872
rect 142804 605820 142856 605872
rect 245476 605820 245528 605872
rect 172428 604528 172480 604580
rect 205548 604528 205600 604580
rect 115204 604460 115256 604512
rect 238484 604460 238536 604512
rect 241796 604460 241848 604512
rect 242808 604460 242860 604512
rect 271880 604460 271932 604512
rect 289728 604460 289780 604512
rect 582840 604460 582892 604512
rect 169024 603168 169076 603220
rect 199108 603168 199160 603220
rect 244924 603168 244976 603220
rect 254676 603168 254728 603220
rect 181812 603100 181864 603152
rect 214380 603100 214432 603152
rect 249708 603100 249760 603152
rect 263600 603100 263652 603152
rect 180064 601740 180116 601792
rect 229100 601740 229152 601792
rect 241060 601740 241112 601792
rect 285680 601740 285732 601792
rect 104164 601672 104216 601724
rect 211252 601672 211304 601724
rect 582748 601672 582800 601724
rect 211804 601604 211856 601656
rect 213184 601604 213236 601656
rect 224224 601604 224276 601656
rect 225236 601604 225288 601656
rect 221372 600788 221424 600840
rect 226340 600788 226392 600840
rect 233884 600652 233936 600704
rect 235356 600652 235408 600704
rect 141424 600380 141476 600432
rect 200396 600380 200448 600432
rect 192484 600312 192536 600364
rect 195428 600312 195480 600364
rect 212448 600312 212500 600364
rect 219532 600312 219584 600364
rect 226340 600312 226392 600364
rect 231768 600312 231820 600364
rect 232228 600312 232280 600364
rect 248328 600312 248380 600364
rect 86960 599564 87012 599616
rect 147680 599564 147732 599616
rect 222660 599428 222712 599480
rect 223028 599428 223080 599480
rect 193404 599088 193456 599140
rect 184204 599020 184256 599072
rect 197636 599020 197688 599072
rect 191196 598952 191248 599004
rect 195612 598952 195664 599004
rect 228640 599020 228692 599072
rect 251456 599020 251508 599072
rect 253296 599020 253348 599072
rect 271972 599020 272024 599072
rect 214748 598952 214800 599004
rect 222844 598952 222896 599004
rect 276112 598952 276164 599004
rect 150164 597592 150216 597644
rect 191012 597592 191064 597644
rect 84108 597524 84160 597576
rect 133696 597524 133748 597576
rect 190368 597524 190420 597576
rect 203340 598884 203392 598936
rect 247684 598884 247736 598936
rect 249064 598884 249116 598936
rect 253480 598884 253532 598936
rect 295340 598204 295392 598256
rect 253480 597524 253532 597576
rect 273260 597524 273312 597576
rect 253388 596776 253440 596828
rect 293960 596776 294012 596828
rect 146944 596232 146996 596284
rect 191380 596232 191432 596284
rect 97264 596164 97316 596216
rect 188252 596164 188304 596216
rect 166356 595416 166408 595468
rect 192668 595416 192720 595468
rect 256608 595416 256660 595468
rect 287060 595416 287112 595468
rect 92480 594804 92532 594856
rect 166356 594804 166408 594856
rect 166632 594804 166684 594856
rect 69848 593376 69900 593428
rect 142620 593376 142672 593428
rect 164884 593376 164936 593428
rect 191288 593376 191340 593428
rect 255412 593376 255464 593428
rect 261024 593376 261076 593428
rect 582656 593376 582708 593428
rect 89720 592628 89772 592680
rect 192576 592628 192628 592680
rect 255412 592628 255464 592680
rect 291200 592628 291252 592680
rect 299480 592628 299532 592680
rect 162124 592016 162176 592068
rect 191380 592016 191432 592068
rect 71780 591268 71832 591320
rect 184296 591268 184348 591320
rect 253388 591268 253440 591320
rect 296720 591268 296772 591320
rect 157984 590656 158036 590708
rect 191288 590656 191340 590708
rect 125508 589908 125560 589960
rect 188436 589908 188488 589960
rect 91376 589296 91428 589348
rect 124220 589296 124272 589348
rect 125508 589296 125560 589348
rect 179236 589296 179288 589348
rect 191380 589296 191432 589348
rect 255412 589296 255464 589348
rect 262404 589296 262456 589348
rect 78128 588616 78180 588668
rect 88248 588616 88300 588668
rect 125600 588616 125652 588668
rect 40040 588548 40092 588600
rect 95332 588548 95384 588600
rect 170404 588548 170456 588600
rect 191656 588548 191708 588600
rect 254676 588548 254728 588600
rect 274732 588548 274784 588600
rect 177948 587120 178000 587172
rect 192484 587120 192536 587172
rect 176016 586508 176068 586560
rect 190460 586508 190512 586560
rect 169668 585828 169720 585880
rect 190552 585828 190604 585880
rect 147496 585760 147548 585812
rect 191748 585760 191800 585812
rect 65984 585148 66036 585200
rect 122196 585148 122248 585200
rect 260748 585148 260800 585200
rect 266360 585148 266412 585200
rect 181444 584400 181496 584452
rect 193404 584400 193456 584452
rect 255412 584400 255464 584452
rect 259460 584400 259512 584452
rect 274824 584400 274876 584452
rect 582380 584400 582432 584452
rect 79968 583788 80020 583840
rect 98552 583788 98604 583840
rect 74264 583720 74316 583772
rect 122104 583720 122156 583772
rect 171784 583720 171836 583772
rect 191748 583720 191800 583772
rect 255504 583720 255556 583772
rect 266360 583720 266412 583772
rect 88248 583176 88300 583228
rect 88984 583176 89036 583228
rect 259368 583040 259420 583092
rect 268384 583040 268436 583092
rect 151728 582972 151780 583024
rect 189724 582972 189776 583024
rect 254584 582972 254636 583024
rect 283104 582972 283156 583024
rect 84108 582632 84160 582684
rect 85028 582632 85080 582684
rect 55128 582428 55180 582480
rect 83004 582428 83056 582480
rect 91008 582428 91060 582480
rect 123484 582428 123536 582480
rect 67364 582360 67416 582412
rect 71044 582360 71096 582412
rect 80704 582360 80756 582412
rect 130476 582360 130528 582412
rect 255412 582360 255464 582412
rect 258172 582360 258224 582412
rect 259368 582360 259420 582412
rect 76288 581068 76340 581120
rect 108304 581068 108356 581120
rect 184848 581068 184900 581120
rect 191196 581068 191248 581120
rect 3332 580932 3384 580984
rect 80244 581000 80296 581052
rect 86592 581000 86644 581052
rect 105544 581000 105596 581052
rect 173164 581000 173216 581052
rect 191748 581000 191800 581052
rect 69020 580660 69072 580712
rect 79048 580660 79100 580712
rect 61936 579708 61988 579760
rect 66904 579708 66956 579760
rect 53748 579640 53800 579692
rect 179052 580388 179104 580440
rect 191012 580388 191064 580440
rect 159364 580252 159416 580304
rect 179328 580252 179380 580304
rect 188436 580252 188488 580304
rect 255504 579708 255556 579760
rect 262220 579708 262272 579760
rect 159364 579640 159416 579692
rect 255412 579640 255464 579692
rect 288716 579640 288768 579692
rect 94964 579572 95016 579624
rect 96712 579572 96764 579624
rect 188988 578280 189040 578332
rect 190920 578280 190972 578332
rect 96896 578212 96948 578264
rect 134524 578212 134576 578264
rect 148968 578212 149020 578264
rect 191656 578212 191708 578264
rect 255320 578212 255372 578264
rect 302240 578212 302292 578264
rect 98552 578144 98604 578196
rect 191748 578144 191800 578196
rect 255412 577056 255464 577108
rect 259552 577056 259604 577108
rect 255412 576852 255464 576904
rect 267740 576852 267792 576904
rect 3424 576784 3476 576836
rect 66168 576784 66220 576836
rect 97908 576784 97960 576836
rect 160744 576784 160796 576836
rect 95884 576104 95936 576156
rect 111064 576104 111116 576156
rect 186136 575560 186188 575612
rect 191656 575560 191708 575612
rect 116584 575492 116636 575544
rect 191748 575492 191800 575544
rect 255412 575492 255464 575544
rect 278780 575492 278832 575544
rect 97908 574744 97960 574796
rect 166448 574744 166500 574796
rect 168288 574744 168340 574796
rect 191288 574744 191340 574796
rect 66076 574064 66128 574116
rect 67364 574064 67416 574116
rect 157248 574064 157300 574116
rect 190828 574064 190880 574116
rect 255412 574064 255464 574116
rect 270500 574064 270552 574116
rect 98000 573316 98052 573368
rect 137100 573316 137152 573368
rect 255964 573316 256016 573368
rect 284300 573316 284352 573368
rect 97540 572976 97592 573028
rect 100760 572976 100812 573028
rect 64788 572704 64840 572756
rect 66812 572704 66864 572756
rect 136640 572704 136692 572756
rect 137100 572704 137152 572756
rect 191748 572704 191800 572756
rect 188436 572636 188488 572688
rect 190828 572636 190880 572688
rect 100760 571956 100812 572008
rect 179420 571956 179472 572008
rect 255412 571412 255464 571464
rect 277492 571412 277544 571464
rect 97724 571344 97776 571396
rect 101404 571344 101456 571396
rect 255504 571344 255556 571396
rect 286324 571344 286376 571396
rect 255412 571276 255464 571328
rect 582564 571276 582616 571328
rect 105544 570596 105596 570648
rect 160100 570596 160152 570648
rect 179420 570596 179472 570648
rect 180524 570596 180576 570648
rect 191748 570596 191800 570648
rect 97908 569916 97960 569968
rect 112536 569916 112588 569968
rect 160100 569916 160152 569968
rect 191748 569916 191800 569968
rect 97908 569168 97960 569220
rect 178684 569168 178736 569220
rect 255504 568624 255556 568676
rect 267924 568624 267976 568676
rect 255412 568556 255464 568608
rect 284392 568556 284444 568608
rect 130384 567808 130436 567860
rect 178776 567808 178828 567860
rect 255688 567808 255740 567860
rect 289820 567808 289872 567860
rect 59268 567196 59320 567248
rect 66904 567196 66956 567248
rect 97908 567196 97960 567248
rect 130384 567196 130436 567248
rect 187056 567196 187108 567248
rect 191380 567196 191432 567248
rect 282000 566448 282052 566500
rect 582472 566448 582524 566500
rect 255504 565904 255556 565956
rect 281540 565904 281592 565956
rect 282000 565904 282052 565956
rect 3424 565836 3476 565888
rect 39304 565836 39356 565888
rect 52368 565836 52420 565888
rect 67640 565836 67692 565888
rect 255596 565836 255648 565888
rect 282920 565836 282972 565888
rect 169576 565156 169628 565208
rect 187608 565156 187660 565208
rect 191748 565156 191800 565208
rect 150256 565088 150308 565140
rect 186964 565088 187016 565140
rect 63408 564408 63460 564460
rect 66444 564408 66496 564460
rect 187700 564408 187752 564460
rect 191288 564408 191340 564460
rect 255504 564408 255556 564460
rect 259460 564408 259512 564460
rect 122196 563660 122248 563712
rect 122748 563660 122800 563712
rect 191748 563660 191800 563712
rect 97908 562300 97960 562352
rect 106188 562300 106240 562352
rect 169024 562300 169076 562352
rect 177856 561688 177908 561740
rect 190920 561688 190972 561740
rect 97908 560940 97960 560992
rect 180064 560940 180116 560992
rect 64696 560328 64748 560380
rect 66812 560328 66864 560380
rect 169484 560260 169536 560312
rect 190828 560260 190880 560312
rect 255504 560260 255556 560312
rect 266452 560260 266504 560312
rect 164056 559512 164108 559564
rect 187700 559512 187752 559564
rect 255504 558968 255556 559020
rect 269212 558968 269264 559020
rect 60648 558900 60700 558952
rect 66812 558900 66864 558952
rect 96896 558900 96948 558952
rect 113824 558900 113876 558952
rect 174544 558900 174596 558952
rect 191748 558900 191800 558952
rect 255596 558900 255648 558952
rect 273352 558900 273404 558952
rect 95148 558832 95200 558884
rect 95332 558832 95384 558884
rect 184204 558832 184256 558884
rect 62028 557540 62080 557592
rect 66812 557540 66864 557592
rect 159916 557540 159968 557592
rect 191748 557540 191800 557592
rect 255596 557540 255648 557592
rect 274640 557540 274692 557592
rect 97908 556792 97960 556844
rect 115204 556792 115256 556844
rect 160836 556792 160888 556844
rect 166356 556792 166408 556844
rect 166356 556180 166408 556232
rect 191748 556180 191800 556232
rect 255596 556180 255648 556232
rect 263692 556180 263744 556232
rect 173716 554820 173768 554872
rect 191472 554820 191524 554872
rect 63316 554752 63368 554804
rect 66536 554752 66588 554804
rect 162216 554752 162268 554804
rect 180064 554752 180116 554804
rect 173256 554004 173308 554056
rect 189724 554004 189776 554056
rect 3424 553664 3476 553716
rect 7564 553664 7616 553716
rect 255596 553460 255648 553512
rect 269488 553460 269540 553512
rect 56416 553392 56468 553444
rect 66904 553392 66956 553444
rect 255688 553392 255740 553444
rect 277584 553392 277636 553444
rect 255596 552644 255648 552696
rect 260748 552644 260800 552696
rect 265072 552644 265124 552696
rect 180616 552100 180668 552152
rect 191104 552100 191156 552152
rect 97908 552032 97960 552084
rect 102048 552032 102100 552084
rect 184204 552032 184256 552084
rect 106188 551284 106240 551336
rect 114744 551284 114796 551336
rect 122104 551284 122156 551336
rect 160192 551284 160244 551336
rect 255596 550672 255648 550724
rect 259644 550672 259696 550724
rect 160192 550604 160244 550656
rect 160744 550604 160796 550656
rect 191748 550604 191800 550656
rect 97816 549856 97868 549908
rect 162308 549856 162360 549908
rect 255596 549856 255648 549908
rect 258080 549856 258132 549908
rect 269120 549856 269172 549908
rect 186044 549312 186096 549364
rect 191748 549312 191800 549364
rect 162308 549244 162360 549296
rect 188528 549244 188580 549296
rect 102048 548496 102100 548548
rect 112444 548496 112496 548548
rect 112536 548496 112588 548548
rect 188436 548496 188488 548548
rect 187516 547884 187568 547936
rect 190644 547884 190696 547936
rect 255596 547884 255648 547936
rect 262312 547884 262364 547936
rect 156604 546524 156656 546576
rect 191656 546524 191708 546576
rect 99380 546456 99432 546508
rect 191564 546456 191616 546508
rect 255504 546456 255556 546508
rect 276204 546456 276256 546508
rect 106924 545708 106976 545760
rect 186964 545708 187016 545760
rect 97080 545232 97132 545284
rect 100024 545232 100076 545284
rect 255504 545232 255556 545284
rect 258356 545232 258408 545284
rect 168196 545096 168248 545148
rect 191656 545096 191708 545148
rect 180064 545028 180116 545080
rect 191564 545028 191616 545080
rect 50988 543736 51040 543788
rect 66812 543736 66864 543788
rect 97540 543736 97592 543788
rect 104256 543736 104308 543788
rect 184756 543736 184808 543788
rect 191012 543736 191064 543788
rect 33784 543668 33836 543720
rect 66260 543668 66312 543720
rect 166448 542988 166500 543040
rect 181536 542988 181588 543040
rect 255596 542444 255648 542496
rect 264980 542444 265032 542496
rect 97540 542376 97592 542428
rect 158812 542376 158864 542428
rect 186320 542376 186372 542428
rect 255504 542376 255556 542428
rect 267832 542376 267884 542428
rect 184664 542308 184716 542360
rect 187056 542308 187108 542360
rect 123484 541696 123536 541748
rect 155776 541696 155828 541748
rect 15844 541628 15896 541680
rect 39948 541628 40000 541680
rect 97908 541628 97960 541680
rect 146944 541628 146996 541680
rect 178408 541628 178460 541680
rect 179144 541628 179196 541680
rect 188344 541628 188396 541680
rect 278044 541628 278096 541680
rect 287152 541628 287204 541680
rect 39948 540948 40000 541000
rect 66260 540948 66312 541000
rect 155776 540948 155828 541000
rect 178408 540948 178460 541000
rect 188528 540540 188580 540592
rect 191656 540540 191708 540592
rect 177396 540200 177448 540252
rect 184756 540200 184808 540252
rect 67824 539792 67876 539844
rect 71780 539792 71832 539844
rect 94136 539656 94188 539708
rect 94780 539656 94832 539708
rect 57796 539588 57848 539640
rect 66260 539588 66312 539640
rect 88156 539588 88208 539640
rect 134616 539588 134668 539640
rect 164332 539588 164384 539640
rect 259552 539656 259604 539708
rect 255504 539588 255556 539640
rect 278872 539588 278924 539640
rect 251456 539316 251508 539368
rect 250444 539248 250496 539300
rect 255780 539248 255832 539300
rect 67640 538840 67692 538892
rect 83464 538840 83516 538892
rect 119344 538840 119396 538892
rect 150440 538840 150492 538892
rect 43444 538296 43496 538348
rect 94596 538296 94648 538348
rect 104164 538296 104216 538348
rect 186320 538296 186372 538348
rect 221372 538296 221424 538348
rect 255504 538296 255556 538348
rect 277400 538296 277452 538348
rect 85580 538228 85632 538280
rect 85764 538228 85816 538280
rect 99380 538228 99432 538280
rect 150440 538228 150492 538280
rect 151636 538228 151688 538280
rect 216404 538228 216456 538280
rect 224684 538228 224736 538280
rect 582932 538228 582984 538280
rect 7564 538160 7616 538212
rect 70676 538160 70728 538212
rect 79968 538160 80020 538212
rect 116584 538160 116636 538212
rect 184204 538160 184256 538212
rect 200396 538160 200448 538212
rect 239220 538160 239272 538212
rect 239404 538160 239456 538212
rect 582380 538160 582432 538212
rect 178684 538092 178736 538144
rect 244372 538092 244424 538144
rect 79232 537684 79284 537736
rect 79968 537684 80020 537736
rect 66076 537480 66128 537532
rect 143632 537480 143684 537532
rect 70676 536800 70728 536852
rect 71044 536800 71096 536852
rect 57244 536732 57296 536784
rect 73252 536732 73304 536784
rect 87696 536732 87748 536784
rect 215300 536732 215352 536784
rect 82176 536664 82228 536716
rect 88156 536664 88208 536716
rect 211988 536664 212040 536716
rect 280804 536664 280856 536716
rect 39304 536052 39356 536104
rect 53656 536052 53708 536104
rect 69388 536052 69440 536104
rect 73252 536052 73304 536104
rect 81440 536052 81492 536104
rect 188344 536052 188396 536104
rect 205548 536052 205600 536104
rect 253204 536052 253256 536104
rect 260840 536052 260892 536104
rect 225236 535984 225288 536036
rect 226984 535984 227036 536036
rect 233424 535780 233476 535832
rect 236644 535780 236696 535832
rect 220084 535508 220136 535560
rect 223396 535508 223448 535560
rect 86224 535440 86276 535492
rect 89812 535440 89864 535492
rect 91008 535440 91060 535492
rect 91836 535440 91888 535492
rect 206376 535440 206428 535492
rect 209964 535440 210016 535492
rect 215944 535440 215996 535492
rect 218980 535440 219032 535492
rect 222844 535440 222896 535492
rect 223948 535440 224000 535492
rect 229652 535440 229704 535492
rect 233884 535440 233936 535492
rect 242992 535440 243044 535492
rect 250628 535440 250680 535492
rect 88248 535372 88300 535424
rect 95424 535372 95476 535424
rect 186964 535372 187016 535424
rect 238208 535372 238260 535424
rect 238668 535372 238720 535424
rect 164332 535304 164384 535356
rect 198004 535304 198056 535356
rect 249064 534760 249116 534812
rect 258172 534760 258224 534812
rect 82728 534692 82780 534744
rect 94688 534692 94740 534744
rect 216036 534692 216088 534744
rect 230388 534692 230440 534744
rect 246396 534692 246448 534744
rect 256884 534692 256936 534744
rect 211988 534420 212040 534472
rect 212724 534420 212776 534472
rect 130476 534012 130528 534064
rect 130936 534012 130988 534064
rect 242992 534012 243044 534064
rect 81440 533400 81492 533452
rect 102784 533400 102836 533452
rect 195980 533400 196032 533452
rect 198832 533400 198884 533452
rect 59176 533332 59228 533384
rect 73160 533332 73212 533384
rect 75828 533332 75880 533384
rect 96804 533332 96856 533384
rect 212540 533332 212592 533384
rect 213460 533332 213512 533384
rect 216680 533332 216732 533384
rect 217324 533332 217376 533384
rect 213184 533196 213236 533248
rect 233424 533400 233476 533452
rect 246948 533400 247000 533452
rect 255872 533400 255924 533452
rect 233240 533332 233292 533384
rect 233700 533332 233752 533384
rect 234620 533332 234672 533384
rect 234988 533332 235040 533384
rect 237380 533332 237432 533384
rect 237564 533332 237616 533384
rect 240140 533332 240192 533384
rect 240692 533332 240744 533384
rect 247040 533332 247092 533384
rect 247684 533332 247736 533384
rect 251916 533332 251968 533384
rect 280344 533332 280396 533384
rect 201500 532720 201552 532772
rect 202052 532720 202104 532772
rect 231860 532720 231912 532772
rect 232412 532720 232464 532772
rect 179144 532652 179196 532704
rect 206836 532652 206888 532704
rect 83096 532040 83148 532092
rect 109684 532040 109736 532092
rect 244372 532040 244424 532092
rect 266544 532040 266596 532092
rect 48228 531972 48280 532024
rect 96896 531972 96948 532024
rect 100024 531972 100076 532024
rect 129004 531972 129056 532024
rect 173164 531972 173216 532024
rect 195428 531972 195480 532024
rect 202972 531972 203024 532024
rect 270592 531972 270644 532024
rect 93124 531292 93176 531344
rect 94044 531292 94096 531344
rect 183376 530612 183428 530664
rect 254216 530612 254268 530664
rect 81992 530544 82044 530596
rect 187608 530544 187660 530596
rect 193036 530544 193088 530596
rect 200212 530544 200264 530596
rect 207664 530544 207716 530596
rect 222292 530544 222344 530596
rect 231216 530544 231268 530596
rect 260932 530544 260984 530596
rect 204628 529184 204680 529236
rect 238024 529184 238076 529236
rect 248512 529184 248564 529236
rect 280252 529184 280304 529236
rect 226248 528572 226300 528624
rect 229100 528572 229152 528624
rect 59268 528504 59320 528556
rect 169760 528504 169812 528556
rect 170496 528504 170548 528556
rect 3424 528436 3476 528488
rect 98000 528436 98052 528488
rect 193128 527892 193180 527944
rect 205640 527892 205692 527944
rect 245660 527892 245712 527944
rect 258264 527892 258316 527944
rect 201592 527824 201644 527876
rect 248512 527824 248564 527876
rect 88340 527076 88392 527128
rect 208492 527076 208544 527128
rect 243544 526464 243596 526516
rect 254032 526464 254084 526516
rect 188988 526396 189040 526448
rect 193312 526396 193364 526448
rect 202144 526396 202196 526448
rect 227812 526396 227864 526448
rect 229836 526396 229888 526448
rect 251272 526396 251324 526448
rect 131028 525104 131080 525156
rect 182916 525104 182968 525156
rect 195980 525104 196032 525156
rect 220084 525104 220136 525156
rect 234712 525104 234764 525156
rect 254676 525104 254728 525156
rect 71872 525036 71924 525088
rect 122840 525036 122892 525088
rect 172336 525036 172388 525088
rect 239404 525036 239456 525088
rect 71044 523676 71096 523728
rect 118700 523676 118752 523728
rect 199384 523676 199436 523728
rect 208400 523676 208452 523728
rect 233332 523676 233384 523728
rect 251272 523676 251324 523728
rect 63316 522928 63368 522980
rect 162216 522928 162268 522980
rect 3424 522248 3476 522300
rect 93124 522248 93176 522300
rect 94504 522248 94556 522300
rect 195244 522248 195296 522300
rect 204444 522248 204496 522300
rect 144828 519528 144880 519580
rect 244924 519528 244976 519580
rect 72424 518168 72476 518220
rect 99380 518168 99432 518220
rect 141976 518168 142028 518220
rect 216772 518168 216824 518220
rect 218704 518168 218756 518220
rect 237472 518168 237524 518220
rect 65984 517216 66036 517268
rect 69664 517216 69716 517268
rect 210424 516808 210476 516860
rect 253940 516808 253992 516860
rect 158444 516740 158496 516792
rect 238760 516740 238812 516792
rect 61936 515380 61988 515432
rect 92572 515380 92624 515432
rect 181996 515380 182048 515432
rect 216036 515380 216088 515432
rect 237564 515380 237616 515432
rect 254584 515380 254636 515432
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 193128 514088 193180 514140
rect 205732 514088 205784 514140
rect 145656 514020 145708 514072
rect 234620 514020 234672 514072
rect 236092 513272 236144 513324
rect 238116 513272 238168 513324
rect 184664 512592 184716 512644
rect 246396 512592 246448 512644
rect 50988 511912 51040 511964
rect 168840 511912 168892 511964
rect 168840 511232 168892 511284
rect 169576 511232 169628 511284
rect 198096 511232 198148 511284
rect 165068 509872 165120 509924
rect 214012 509872 214064 509924
rect 154488 508512 154540 508564
rect 229836 508512 229888 508564
rect 139308 507084 139360 507136
rect 267924 507084 267976 507136
rect 187516 505792 187568 505844
rect 214564 505792 214616 505844
rect 136548 505724 136600 505776
rect 219440 505724 219492 505776
rect 186964 504432 187016 504484
rect 244464 504432 244516 504484
rect 143356 504364 143408 504416
rect 231952 504364 232004 504416
rect 189724 503004 189776 503056
rect 215944 503004 215996 503056
rect 205088 502936 205140 502988
rect 240232 502936 240284 502988
rect 76012 502256 76064 502308
rect 77208 502256 77260 502308
rect 212632 501712 212684 501764
rect 213276 501712 213328 501764
rect 188436 501644 188488 501696
rect 262404 501644 262456 501696
rect 77208 501576 77260 501628
rect 212632 501576 212684 501628
rect 142068 500216 142120 500268
rect 250444 500216 250496 500268
rect 155684 498788 155736 498840
rect 229744 498788 229796 498840
rect 242900 498788 242952 498840
rect 291384 498788 291436 498840
rect 192576 497428 192628 497480
rect 203524 497428 203576 497480
rect 220820 497428 220872 497480
rect 256792 497428 256844 497480
rect 162676 496068 162728 496120
rect 254124 496068 254176 496120
rect 244372 495456 244424 495508
rect 298100 495456 298152 495508
rect 127624 494708 127676 494760
rect 244372 494708 244424 494760
rect 242900 493960 242952 494012
rect 243544 493960 243596 494012
rect 246304 493348 246356 493400
rect 251824 493348 251876 493400
rect 163964 493280 164016 493332
rect 206376 493280 206428 493332
rect 223488 493280 223540 493332
rect 253388 493280 253440 493332
rect 132408 492668 132460 492720
rect 242900 492668 242952 492720
rect 196624 491988 196676 492040
rect 218704 491988 218756 492040
rect 171876 491920 171928 491972
rect 213184 491920 213236 491972
rect 222108 491920 222160 491972
rect 247132 491920 247184 491972
rect 239404 491308 239456 491360
rect 241428 491308 241480 491360
rect 198096 490628 198148 490680
rect 215944 490628 215996 490680
rect 176108 490560 176160 490612
rect 200304 490560 200356 490612
rect 142896 488520 142948 488572
rect 143448 488520 143500 488572
rect 232596 488520 232648 488572
rect 104256 488452 104308 488504
rect 198832 488452 198884 488504
rect 226984 488180 227036 488232
rect 229100 488180 229152 488232
rect 198832 487840 198884 487892
rect 227076 487840 227128 487892
rect 175004 487772 175056 487824
rect 198740 487772 198792 487824
rect 199476 487772 199528 487824
rect 241612 487772 241664 487824
rect 104256 487160 104308 487212
rect 104808 487160 104860 487212
rect 160008 486412 160060 486464
rect 174544 486412 174596 486464
rect 179420 485732 179472 485784
rect 180524 485732 180576 485784
rect 580172 485732 580224 485784
rect 153108 485052 153160 485104
rect 179420 485052 179472 485104
rect 144736 484372 144788 484424
rect 241428 484372 241480 484424
rect 252560 484372 252612 484424
rect 93952 483624 94004 483676
rect 94596 483624 94648 483676
rect 209872 483624 209924 483676
rect 210608 483624 210660 483676
rect 226156 482944 226208 482996
rect 226340 482944 226392 482996
rect 226432 481652 226484 481704
rect 245568 481652 245620 481704
rect 248420 481652 248472 481704
rect 192484 480904 192536 480956
rect 215300 480904 215352 480956
rect 146944 480224 146996 480276
rect 240784 480224 240836 480276
rect 175096 479544 175148 479596
rect 202144 479544 202196 479596
rect 210608 479544 210660 479596
rect 227812 479544 227864 479596
rect 233240 479544 233292 479596
rect 252560 479544 252612 479596
rect 111064 479476 111116 479528
rect 251272 479476 251324 479528
rect 110420 478864 110472 478916
rect 111064 478864 111116 478916
rect 251272 478864 251324 478916
rect 251916 478864 251968 478916
rect 168104 478184 168156 478236
rect 211160 478184 211212 478236
rect 35164 478116 35216 478168
rect 43444 478116 43496 478168
rect 126244 478116 126296 478168
rect 208492 478116 208544 478168
rect 277676 478116 277728 478168
rect 218152 476824 218204 476876
rect 250444 476824 250496 476876
rect 85488 476756 85540 476808
rect 94136 476756 94188 476808
rect 102140 476756 102192 476808
rect 102784 476756 102836 476808
rect 259644 476756 259696 476808
rect 3332 475328 3384 475380
rect 35164 475328 35216 475380
rect 133144 475192 133196 475244
rect 133696 475192 133748 475244
rect 106924 474784 106976 474836
rect 241704 474784 241756 474836
rect 242164 474784 242216 474836
rect 133696 474716 133748 474768
rect 291292 474716 291344 474768
rect 240140 473968 240192 474020
rect 256884 473968 256936 474020
rect 133236 473356 133288 473408
rect 270592 473356 270644 473408
rect 79968 472608 80020 472660
rect 101404 472608 101456 472660
rect 148324 472064 148376 472116
rect 229100 472064 229152 472116
rect 284484 472064 284536 472116
rect 105544 471996 105596 472048
rect 258080 471996 258132 472048
rect 216772 471316 216824 471368
rect 265072 471316 265124 471368
rect 79324 471248 79376 471300
rect 91192 471248 91244 471300
rect 111064 471248 111116 471300
rect 158720 471248 158772 471300
rect 166816 471248 166868 471300
rect 169484 471248 169536 471300
rect 255504 471248 255556 471300
rect 116584 469820 116636 469872
rect 150164 469820 150216 469872
rect 281632 469820 281684 469872
rect 90364 469208 90416 469260
rect 91008 469208 91060 469260
rect 187056 469208 187108 469260
rect 187608 469208 187660 469260
rect 253480 469208 253532 469260
rect 180524 468528 180576 468580
rect 213920 468528 213972 468580
rect 245568 468528 245620 468580
rect 265716 468528 265768 468580
rect 114468 468460 114520 468512
rect 258264 468460 258316 468512
rect 113824 467848 113876 467900
rect 114468 467848 114520 467900
rect 149704 466488 149756 466540
rect 181536 466488 181588 466540
rect 182088 466488 182140 466540
rect 227720 466488 227772 466540
rect 290004 466488 290056 466540
rect 175924 466420 175976 466472
rect 248420 466420 248472 466472
rect 182088 465672 182140 465724
rect 215300 465672 215352 465724
rect 223580 465672 223632 465724
rect 246948 465672 247000 465724
rect 262864 465672 262916 465724
rect 94504 465536 94556 465588
rect 95148 465536 95200 465588
rect 95148 465060 95200 465112
rect 217416 465060 217468 465112
rect 236000 465060 236052 465112
rect 271972 465060 272024 465112
rect 272524 465060 272576 465112
rect 162308 464992 162360 465044
rect 162768 464992 162820 465044
rect 187700 464992 187752 465044
rect 241428 464380 241480 464432
rect 259644 464380 259696 464432
rect 98644 464312 98696 464364
rect 162768 464312 162820 464364
rect 193036 464312 193088 464364
rect 212540 464312 212592 464364
rect 227076 464312 227128 464364
rect 245660 464312 245712 464364
rect 279424 464312 279476 464364
rect 289820 464312 289872 464364
rect 159364 463700 159416 463752
rect 197360 463700 197412 463752
rect 205548 462952 205600 463004
rect 270500 462952 270552 463004
rect 3240 462340 3292 462392
rect 17224 462340 17276 462392
rect 112444 462340 112496 462392
rect 249064 462340 249116 462392
rect 137744 461592 137796 461644
rect 152556 461592 152608 461644
rect 213828 461592 213880 461644
rect 278780 461592 278832 461644
rect 201500 461456 201552 461508
rect 202144 461456 202196 461508
rect 185676 461320 185728 461372
rect 186136 461320 186188 461372
rect 174544 460980 174596 461032
rect 201500 460980 201552 461032
rect 61936 460912 61988 460964
rect 74540 460912 74592 460964
rect 186136 460912 186188 460964
rect 259736 460912 259788 460964
rect 85580 460844 85632 460896
rect 105544 460844 105596 460896
rect 62028 460164 62080 460216
rect 85672 460164 85724 460216
rect 217416 460164 217468 460216
rect 233148 460164 233200 460216
rect 104900 459892 104952 459944
rect 105544 459892 105596 459944
rect 137836 459620 137888 459672
rect 213276 459620 213328 459672
rect 213828 459620 213880 459672
rect 215300 459620 215352 459672
rect 216036 459620 216088 459672
rect 153844 459552 153896 459604
rect 252560 459552 252612 459604
rect 253572 459552 253624 459604
rect 68284 458804 68336 458856
rect 90364 458804 90416 458856
rect 96528 458804 96580 458856
rect 142896 458804 142948 458856
rect 169484 458804 169536 458856
rect 176016 458804 176068 458856
rect 241520 458804 241572 458856
rect 254308 458804 254360 458856
rect 254676 458804 254728 458856
rect 270500 458804 270552 458856
rect 204536 458600 204588 458652
rect 205548 458600 205600 458652
rect 52184 458260 52236 458312
rect 149796 458260 149848 458312
rect 178684 458260 178736 458312
rect 204536 458260 204588 458312
rect 142988 458192 143040 458244
rect 247408 458192 247460 458244
rect 277584 458124 277636 458176
rect 214564 457512 214616 457564
rect 234436 457512 234488 457564
rect 162768 457444 162820 457496
rect 173716 457444 173768 457496
rect 218888 457444 218940 457496
rect 70308 456764 70360 456816
rect 194600 456764 194652 456816
rect 195060 456764 195112 456816
rect 225052 456764 225104 456816
rect 226156 456764 226208 456816
rect 302332 456764 302384 456816
rect 288348 456016 288400 456068
rect 580172 456016 580224 456068
rect 238760 455880 238812 455932
rect 239404 455880 239456 455932
rect 48228 455472 48280 455524
rect 144184 455472 144236 455524
rect 185584 455472 185636 455524
rect 196072 455472 196124 455524
rect 239404 455472 239456 455524
rect 277492 455472 277544 455524
rect 82728 455404 82780 455456
rect 211160 455404 211212 455456
rect 220084 455404 220136 455456
rect 269764 455404 269816 455456
rect 75184 455336 75236 455388
rect 75828 455336 75880 455388
rect 185584 455336 185636 455388
rect 222568 455064 222620 455116
rect 223488 455064 223540 455116
rect 243544 454656 243596 454708
rect 258080 454656 258132 454708
rect 270868 454656 270920 454708
rect 189080 454112 189132 454164
rect 187056 454044 187108 454096
rect 193588 454044 193640 454096
rect 209780 454044 209832 454096
rect 210424 454044 210476 454096
rect 222568 454044 222620 454096
rect 258080 454044 258132 454096
rect 202144 453976 202196 454028
rect 207020 453976 207072 454028
rect 214564 453976 214616 454028
rect 215944 453976 215996 454028
rect 227812 453976 227864 454028
rect 228732 453976 228784 454028
rect 230756 453976 230808 454028
rect 232596 453976 232648 454028
rect 248604 453976 248656 454028
rect 249708 453976 249760 454028
rect 251548 453976 251600 454028
rect 251916 453976 251968 454028
rect 249064 453908 249116 453960
rect 253388 453908 253440 453960
rect 265716 453296 265768 453348
rect 274916 453296 274968 453348
rect 221188 453160 221240 453212
rect 223672 453160 223724 453212
rect 66076 453024 66128 453076
rect 70492 453024 70544 453076
rect 180064 452684 180116 452736
rect 180616 452684 180668 452736
rect 207940 452684 207992 452736
rect 236460 452684 236512 452736
rect 244280 452684 244332 452736
rect 77668 452616 77720 452668
rect 160836 452616 160888 452668
rect 200212 452616 200264 452668
rect 234436 452616 234488 452668
rect 262404 452616 262456 452668
rect 199292 452548 199344 452600
rect 199476 452548 199528 452600
rect 210516 451868 210568 451920
rect 251088 451868 251140 451920
rect 176476 451324 176528 451376
rect 199292 451324 199344 451376
rect 240140 451324 240192 451376
rect 241428 451324 241480 451376
rect 257344 451324 257396 451376
rect 101404 451256 101456 451308
rect 129096 451256 129148 451308
rect 241060 451256 241112 451308
rect 250628 451256 250680 451308
rect 255228 451256 255280 451308
rect 288532 451256 288584 451308
rect 582656 451256 582708 451308
rect 68928 450576 68980 450628
rect 80060 450576 80112 450628
rect 95148 450576 95200 450628
rect 96712 450576 96764 450628
rect 107936 450576 107988 450628
rect 142160 450644 142212 450696
rect 142988 450644 143040 450696
rect 77300 450508 77352 450560
rect 113824 450508 113876 450560
rect 154396 450508 154448 450560
rect 255228 450508 255280 450560
rect 298284 450508 298336 450560
rect 251180 450440 251232 450492
rect 259644 450440 259696 450492
rect 250444 450236 250496 450288
rect 254124 450236 254176 450288
rect 166448 449896 166500 449948
rect 167644 449896 167696 449948
rect 183376 449896 183428 449948
rect 184940 449896 184992 449948
rect 186228 449896 186280 449948
rect 205640 449896 205692 449948
rect 191932 449692 191984 449744
rect 202328 449692 202380 449744
rect 251824 449692 251876 449744
rect 253940 449692 253992 449744
rect 253480 449556 253532 449608
rect 255688 449556 255740 449608
rect 254584 449216 254636 449268
rect 265072 449216 265124 449268
rect 147772 449148 147824 449200
rect 148876 449148 148928 449200
rect 188344 449148 188396 449200
rect 255596 449148 255648 449200
rect 276020 449148 276072 449200
rect 70860 448604 70912 448656
rect 147772 448604 147824 448656
rect 3148 448536 3200 448588
rect 40684 448536 40736 448588
rect 63224 448536 63276 448588
rect 166264 448536 166316 448588
rect 166448 448468 166500 448520
rect 190460 448468 190512 448520
rect 191840 448400 191892 448452
rect 193404 448400 193456 448452
rect 73160 447788 73212 447840
rect 77668 447788 77720 447840
rect 131764 447788 131816 447840
rect 154396 447788 154448 447840
rect 254492 447448 254544 447500
rect 258724 447448 258776 447500
rect 167000 447040 167052 447092
rect 168196 447040 168248 447092
rect 191564 447040 191616 447092
rect 255504 447040 255556 447092
rect 277584 447040 277636 447092
rect 283012 447040 283064 447092
rect 95240 446428 95292 446480
rect 148324 446428 148376 446480
rect 71136 446360 71188 446412
rect 167000 446360 167052 446412
rect 67640 445680 67692 445732
rect 70860 445680 70912 445732
rect 137836 445680 137888 445732
rect 138020 445680 138072 445732
rect 158720 445680 158772 445732
rect 159364 445680 159416 445732
rect 77116 445000 77168 445052
rect 86224 445000 86276 445052
rect 86868 445000 86920 445052
rect 138020 445000 138072 445052
rect 153016 445000 153068 445052
rect 190368 445000 190420 445052
rect 191564 445000 191616 445052
rect 83464 444456 83516 444508
rect 86868 444456 86920 444508
rect 101404 444456 101456 444508
rect 104164 444456 104216 444508
rect 70400 444388 70452 444440
rect 158720 444388 158772 444440
rect 173164 444320 173216 444372
rect 180064 444320 180116 444372
rect 255504 443640 255556 443692
rect 260564 443640 260616 443692
rect 78680 443028 78732 443080
rect 173164 443028 173216 443080
rect 66168 442960 66220 443012
rect 193036 442960 193088 443012
rect 270592 442960 270644 443012
rect 77208 442892 77260 442944
rect 83188 442892 83240 442944
rect 184756 442892 184808 442944
rect 184940 442892 184992 442944
rect 269304 442892 269356 442944
rect 262864 442280 262916 442332
rect 272064 442280 272116 442332
rect 260564 442212 260616 442264
rect 269304 442212 269356 442264
rect 88248 441668 88300 441720
rect 184204 441668 184256 441720
rect 67732 441600 67784 441652
rect 184756 441600 184808 441652
rect 191380 441600 191432 441652
rect 64696 440852 64748 440904
rect 186044 440852 186096 440904
rect 190644 440852 190696 440904
rect 78588 440240 78640 440292
rect 174544 440240 174596 440292
rect 155684 440172 155736 440224
rect 191656 440172 191708 440224
rect 4804 439492 4856 439544
rect 103796 439492 103848 439544
rect 177948 439492 178000 439544
rect 185584 439492 185636 439544
rect 255504 439492 255556 439544
rect 288624 439492 288676 439544
rect 104808 438948 104860 439000
rect 107660 438948 107712 439000
rect 67364 438880 67416 438932
rect 154028 438880 154080 438932
rect 103796 438812 103848 438864
rect 104440 438812 104492 438864
rect 106924 438812 106976 438864
rect 178040 438132 178092 438184
rect 179236 438132 179288 438184
rect 190644 438132 190696 438184
rect 255504 438132 255556 438184
rect 281632 438132 281684 438184
rect 67272 437452 67324 437504
rect 67548 437452 67600 437504
rect 147036 437452 147088 437504
rect 255504 437452 255556 437504
rect 296812 437452 296864 437504
rect 102508 436772 102560 436824
rect 111064 436772 111116 436824
rect 177948 436772 178000 436824
rect 184664 436772 184716 436824
rect 191656 436772 191708 436824
rect 110788 436704 110840 436756
rect 186320 436704 186372 436756
rect 255688 436704 255740 436756
rect 285956 436704 286008 436756
rect 94044 436636 94096 436688
rect 98644 436636 98696 436688
rect 78220 436364 78272 436416
rect 79324 436364 79376 436416
rect 59268 436160 59320 436212
rect 69664 436160 69716 436212
rect 70032 436160 70084 436212
rect 81164 436160 81216 436212
rect 88984 436160 89036 436212
rect 15844 436092 15896 436144
rect 70860 436092 70912 436144
rect 75184 436092 75236 436144
rect 87328 436092 87380 436144
rect 88248 436092 88300 436144
rect 148324 435344 148376 435396
rect 185676 435344 185728 435396
rect 255504 435344 255556 435396
rect 259736 435344 259788 435396
rect 276296 435344 276348 435396
rect 65892 434800 65944 434852
rect 158812 434800 158864 434852
rect 3424 434732 3476 434784
rect 112444 434732 112496 434784
rect 272524 434732 272576 434784
rect 295524 434732 295576 434784
rect 67548 434664 67600 434716
rect 71320 434664 71372 434716
rect 115756 434664 115808 434716
rect 146944 434664 146996 434716
rect 187056 434664 187108 434716
rect 189080 434664 189132 434716
rect 255504 434664 255556 434716
rect 68652 434052 68704 434104
rect 71780 434052 71832 434104
rect 72700 434052 72752 434104
rect 53748 433984 53800 434036
rect 61752 433984 61804 434036
rect 66812 433984 66864 434036
rect 72608 433984 72660 434036
rect 132500 433984 132552 434036
rect 73988 433644 74040 433696
rect 52368 432624 52420 432676
rect 115848 433236 115900 433288
rect 150256 433236 150308 433288
rect 150532 433236 150584 433288
rect 151084 433168 151136 433220
rect 255964 432624 256016 432676
rect 256884 432624 256936 432676
rect 266636 432624 266688 432676
rect 53656 432556 53708 432608
rect 145656 432556 145708 432608
rect 258724 432556 258776 432608
rect 271972 432556 272024 432608
rect 115572 431876 115624 431928
rect 126244 431876 126296 431928
rect 155776 431876 155828 431928
rect 178040 431876 178092 431928
rect 191656 431944 191708 431996
rect 112904 431196 112956 431248
rect 124864 431196 124916 431248
rect 154028 431196 154080 431248
rect 170496 431196 170548 431248
rect 191748 431196 191800 431248
rect 255412 431196 255464 431248
rect 289912 431196 289964 431248
rect 65800 430652 65852 430704
rect 66076 430652 66128 430704
rect 63316 430584 63368 430636
rect 67548 430584 67600 430636
rect 115756 430516 115808 430568
rect 133236 430516 133288 430568
rect 166356 430516 166408 430568
rect 191012 430516 191064 430568
rect 139308 429836 139360 429888
rect 155316 429836 155368 429888
rect 60556 429224 60608 429276
rect 66076 429224 66128 429276
rect 66628 429224 66680 429276
rect 115848 429088 115900 429140
rect 151268 429088 151320 429140
rect 152924 429088 152976 429140
rect 190828 429088 190880 429140
rect 176660 427728 176712 427780
rect 190828 427728 190880 427780
rect 119344 427048 119396 427100
rect 133144 427048 133196 427100
rect 151636 427048 151688 427100
rect 176660 427048 176712 427100
rect 285772 427048 285824 427100
rect 291292 427048 291344 427100
rect 582564 427048 582616 427100
rect 64696 426436 64748 426488
rect 66812 426436 66864 426488
rect 255412 426436 255464 426488
rect 285772 426436 285824 426488
rect 115848 426368 115900 426420
rect 124220 426368 124272 426420
rect 255504 426368 255556 426420
rect 273536 426368 273588 426420
rect 41328 425688 41380 425740
rect 65800 425688 65852 425740
rect 66628 425688 66680 425740
rect 173808 425688 173860 425740
rect 191748 425688 191800 425740
rect 273536 425688 273588 425740
rect 283196 425688 283248 425740
rect 115848 425008 115900 425060
rect 155224 425008 155276 425060
rect 175188 424328 175240 424380
rect 186136 424328 186188 424380
rect 191748 424328 191800 424380
rect 53748 423648 53800 423700
rect 66812 423648 66864 423700
rect 115848 423580 115900 423632
rect 118700 423580 118752 423632
rect 148324 423580 148376 423632
rect 155868 423580 155920 423632
rect 158812 423580 158864 423632
rect 191012 423580 191064 423632
rect 50988 422288 51040 422340
rect 66260 422288 66312 422340
rect 255504 422288 255556 422340
rect 281816 422288 281868 422340
rect 64604 421064 64656 421116
rect 67180 421064 67232 421116
rect 48136 420928 48188 420980
rect 66904 420928 66956 420980
rect 143448 420928 143500 420980
rect 192484 420928 192536 420980
rect 255504 420928 255556 420980
rect 298376 420928 298428 420980
rect 155592 420860 155644 420912
rect 191748 420860 191800 420912
rect 263784 420180 263836 420232
rect 264888 420180 264940 420232
rect 298100 420180 298152 420232
rect 255504 419500 255556 419552
rect 263784 419500 263836 419552
rect 149796 419432 149848 419484
rect 191748 419432 191800 419484
rect 255412 419432 255464 419484
rect 285680 419432 285732 419484
rect 287428 419432 287480 419484
rect 582380 419432 582432 419484
rect 115848 419364 115900 419416
rect 153844 419364 153896 419416
rect 176568 418752 176620 418804
rect 187700 418752 187752 418804
rect 61660 418208 61712 418260
rect 63224 418208 63276 418260
rect 66628 418208 66680 418260
rect 61936 418072 61988 418124
rect 66996 418072 67048 418124
rect 281448 418072 281500 418124
rect 582472 418072 582524 418124
rect 148876 417392 148928 417444
rect 166356 417392 166408 417444
rect 255412 417392 255464 417444
rect 280436 417392 280488 417444
rect 281448 417392 281500 417444
rect 118700 417188 118752 417240
rect 119344 417188 119396 417240
rect 115848 416780 115900 416832
rect 118700 416780 118752 416832
rect 126244 416780 126296 416832
rect 154396 416780 154448 416832
rect 166356 416780 166408 416832
rect 166724 416780 166776 416832
rect 191748 416780 191800 416832
rect 255412 416780 255464 416832
rect 265164 416780 265216 416832
rect 149060 416100 149112 416152
rect 150256 416100 150308 416152
rect 169760 416100 169812 416152
rect 50896 416032 50948 416084
rect 56416 416032 56468 416084
rect 66812 416032 66864 416084
rect 120080 416032 120132 416084
rect 151176 416032 151228 416084
rect 153108 416032 153160 416084
rect 190644 416032 190696 416084
rect 115848 415420 115900 415472
rect 120080 415420 120132 415472
rect 122196 415420 122248 415472
rect 149060 415420 149112 415472
rect 144184 415352 144236 415404
rect 191472 415352 191524 415404
rect 184848 415284 184900 415336
rect 188344 415284 188396 415336
rect 115848 414672 115900 414724
rect 122748 414672 122800 414724
rect 125692 414672 125744 414724
rect 55036 413992 55088 414044
rect 66812 413992 66864 414044
rect 115756 413924 115808 413976
rect 127624 413924 127676 413976
rect 255412 413788 255464 413840
rect 259644 413788 259696 413840
rect 114744 413584 114796 413636
rect 117320 413584 117372 413636
rect 55128 413244 55180 413296
rect 66628 413244 66680 413296
rect 184848 412632 184900 412684
rect 191748 412632 191800 412684
rect 255412 412428 255464 412480
rect 258264 412428 258316 412480
rect 115020 411884 115072 411936
rect 122840 411884 122892 411936
rect 123484 411884 123536 411936
rect 147036 411884 147088 411936
rect 158812 411884 158864 411936
rect 260104 411884 260156 411936
rect 288716 411884 288768 411936
rect 61936 411272 61988 411324
rect 66904 411272 66956 411324
rect 158812 411272 158864 411324
rect 159364 411272 159416 411324
rect 192852 411272 192904 411324
rect 52184 411204 52236 411256
rect 66812 411204 66864 411256
rect 115572 411204 115624 411256
rect 122196 411204 122248 411256
rect 44088 410524 44140 410576
rect 52184 410524 52236 410576
rect 177856 410524 177908 410576
rect 190460 410524 190512 410576
rect 187516 410388 187568 410440
rect 189080 410388 189132 410440
rect 2780 410184 2832 410236
rect 4804 410184 4856 410236
rect 121460 409844 121512 409896
rect 155776 409844 155828 409896
rect 160100 409844 160152 409896
rect 115848 409776 115900 409828
rect 126244 409776 126296 409828
rect 49608 408484 49660 408536
rect 66812 408484 66864 408536
rect 115848 408484 115900 408536
rect 151176 408484 151228 408536
rect 191748 408484 191800 408536
rect 255412 408484 255464 408536
rect 270776 408484 270828 408536
rect 276112 408484 276164 408536
rect 39856 408416 39908 408468
rect 48228 408416 48280 408468
rect 66904 408416 66956 408468
rect 140688 408416 140740 408468
rect 186320 408416 186372 408468
rect 255412 407804 255464 407856
rect 259644 407804 259696 407856
rect 265072 407804 265124 407856
rect 159916 407736 159968 407788
rect 167000 407736 167052 407788
rect 255504 407736 255556 407788
rect 273536 407736 273588 407788
rect 167000 407124 167052 407176
rect 191656 407124 191708 407176
rect 113088 407056 113140 407108
rect 131764 407056 131816 407108
rect 57888 406376 57940 406428
rect 64788 406376 64840 406428
rect 66812 406376 66864 406428
rect 154488 406376 154540 406428
rect 191748 406376 191800 406428
rect 255504 405696 255556 405748
rect 276112 405696 276164 405748
rect 115848 405628 115900 405680
rect 121460 405628 121512 405680
rect 152924 405628 152976 405680
rect 154488 405628 154540 405680
rect 63224 404336 63276 404388
rect 66812 404336 66864 404388
rect 115848 404336 115900 404388
rect 153844 404404 153896 404456
rect 162216 404336 162268 404388
rect 162584 404336 162636 404388
rect 177488 404336 177540 404388
rect 164056 404268 164108 404320
rect 169760 404268 169812 404320
rect 53656 403588 53708 403640
rect 67640 403588 67692 403640
rect 119988 403588 120040 403640
rect 162584 403588 162636 403640
rect 172428 403588 172480 403640
rect 182916 403588 182968 403640
rect 115848 402976 115900 403028
rect 148324 402976 148376 403028
rect 169760 402976 169812 403028
rect 191748 402976 191800 403028
rect 256884 402976 256936 403028
rect 291292 402976 291344 403028
rect 255320 402908 255372 402960
rect 287152 402908 287204 402960
rect 185584 401820 185636 401872
rect 193128 401820 193180 401872
rect 116584 401616 116636 401668
rect 181444 401616 181496 401668
rect 186044 401004 186096 401056
rect 186964 401004 187016 401056
rect 118884 400868 118936 400920
rect 143540 400868 143592 400920
rect 172060 400868 172112 400920
rect 191564 400868 191616 400920
rect 115572 400664 115624 400716
rect 119988 400664 120040 400716
rect 115756 400528 115808 400580
rect 122196 400528 122248 400580
rect 59084 400188 59136 400240
rect 66812 400188 66864 400240
rect 123668 400188 123720 400240
rect 186044 400188 186096 400240
rect 255412 400188 255464 400240
rect 280436 400188 280488 400240
rect 148968 399440 149020 399492
rect 181536 399440 181588 399492
rect 115848 398896 115900 398948
rect 137284 398896 137336 398948
rect 53656 398828 53708 398880
rect 66812 398828 66864 398880
rect 129004 398828 129056 398880
rect 190276 398828 190328 398880
rect 191748 398828 191800 398880
rect 255412 398828 255464 398880
rect 60648 398760 60700 398812
rect 65892 398760 65944 398812
rect 66536 398760 66588 398812
rect 268384 398760 268436 398812
rect 274824 398760 274876 398812
rect 115848 398284 115900 398336
rect 116032 398284 116084 398336
rect 118884 398284 118936 398336
rect 255412 398216 255464 398268
rect 258908 398216 258960 398268
rect 118884 398148 118936 398200
rect 147496 398148 147548 398200
rect 173256 398148 173308 398200
rect 175004 398148 175056 398200
rect 180156 398148 180208 398200
rect 145656 398080 145708 398132
rect 188896 398080 188948 398132
rect 189724 398080 189776 398132
rect 183560 398012 183612 398064
rect 191748 398080 191800 398132
rect 265624 398080 265676 398132
rect 275008 398080 275060 398132
rect 36544 397468 36596 397520
rect 67088 397468 67140 397520
rect 163504 397400 163556 397452
rect 163964 397400 164016 397452
rect 140044 396720 140096 396772
rect 180524 396720 180576 396772
rect 187148 396720 187200 396772
rect 115112 396516 115164 396568
rect 118884 396516 118936 396568
rect 115572 396040 115624 396092
rect 122104 396040 122156 396092
rect 163504 396040 163556 396092
rect 192484 396040 192536 396092
rect 57704 395292 57756 395344
rect 67272 395292 67324 395344
rect 168288 395292 168340 395344
rect 176108 395292 176160 395344
rect 164056 394952 164108 395004
rect 164976 394952 165028 395004
rect 115848 394748 115900 394800
rect 151084 394748 151136 394800
rect 115848 394612 115900 394664
rect 157984 394680 158036 394732
rect 161480 394680 161532 394732
rect 162676 394680 162728 394732
rect 191840 394680 191892 394732
rect 155316 394612 155368 394664
rect 155960 394612 156012 394664
rect 117228 393932 117280 393984
rect 136640 393932 136692 393984
rect 61844 393388 61896 393440
rect 65984 393388 66036 393440
rect 177396 393320 177448 393372
rect 191012 393320 191064 393372
rect 255504 393320 255556 393372
rect 278964 393320 279016 393372
rect 160100 393252 160152 393304
rect 161388 393252 161440 393304
rect 191932 393252 191984 393304
rect 148416 392640 148468 392692
rect 161480 392640 161532 392692
rect 144184 392572 144236 392624
rect 160100 392572 160152 392624
rect 253664 392572 253716 392624
rect 279424 392572 279476 392624
rect 115940 392300 115992 392352
rect 117228 392300 117280 392352
rect 57704 391960 57756 392012
rect 66812 391960 66864 392012
rect 115848 391960 115900 392012
rect 145656 391960 145708 392012
rect 162216 391960 162268 392012
rect 171876 391960 171928 392012
rect 172428 391960 172480 392012
rect 254308 391960 254360 392012
rect 255320 391960 255372 392012
rect 35164 391280 35216 391332
rect 68560 391280 68612 391332
rect 4804 391212 4856 391264
rect 68560 391076 68612 391128
rect 93952 390940 94004 390992
rect 94964 390940 95016 390992
rect 112720 391280 112772 391332
rect 116584 391280 116636 391332
rect 253572 391280 253624 391332
rect 295340 391280 295392 391332
rect 173624 391212 173676 391264
rect 107292 390940 107344 390992
rect 264244 391212 264296 391264
rect 280344 391212 280396 391264
rect 286324 391212 286376 391264
rect 292580 391212 292632 391264
rect 580264 391212 580316 391264
rect 194140 390940 194192 390992
rect 112720 390872 112772 390924
rect 191840 390872 191892 390924
rect 195980 390872 196032 390924
rect 171968 390600 172020 390652
rect 173624 390600 173676 390652
rect 158444 390532 158496 390584
rect 163596 390532 163648 390584
rect 191748 390532 191800 390584
rect 251824 390532 251876 390584
rect 259644 390532 259696 390584
rect 67640 390124 67692 390176
rect 68790 390124 68842 390176
rect 154488 389852 154540 389904
rect 164884 389852 164936 389904
rect 160100 389784 160152 389836
rect 160744 389784 160796 389836
rect 186412 389784 186464 389836
rect 40684 389240 40736 389292
rect 100760 389240 100812 389292
rect 110788 389240 110840 389292
rect 141424 389240 141476 389292
rect 187148 389240 187200 389292
rect 215300 389240 215352 389292
rect 238760 389240 238812 389292
rect 239036 389240 239088 389292
rect 260104 389240 260156 389292
rect 17224 389172 17276 389224
rect 81716 389172 81768 389224
rect 98920 389172 98972 389224
rect 160100 389172 160152 389224
rect 178868 389172 178920 389224
rect 200212 389172 200264 389224
rect 201592 389172 201644 389224
rect 267832 389172 267884 389224
rect 169024 389104 169076 389156
rect 169484 389104 169536 389156
rect 205916 389104 205968 389156
rect 253388 389104 253440 389156
rect 276204 389104 276256 389156
rect 172428 389036 172480 389088
rect 202972 389036 203024 389088
rect 250720 389036 250772 389088
rect 253664 389036 253716 389088
rect 164884 388560 164936 388612
rect 171784 388560 171836 388612
rect 59176 388424 59228 388476
rect 67364 388424 67416 388476
rect 71044 388424 71096 388476
rect 82728 388424 82780 388476
rect 108396 388424 108448 388476
rect 233332 388424 233384 388476
rect 245844 388424 245896 388476
rect 247684 388424 247736 388476
rect 251364 388424 251416 388476
rect 262864 388424 262916 388476
rect 291384 388424 291436 388476
rect 71688 388356 71740 388408
rect 238116 388356 238168 388408
rect 239404 388356 239456 388408
rect 71688 387948 71740 388000
rect 72516 387948 72568 388000
rect 83188 387880 83240 387932
rect 84108 387880 84160 387932
rect 70860 387812 70912 387864
rect 72516 387812 72568 387864
rect 77208 387812 77260 387864
rect 78036 387812 78088 387864
rect 88248 387744 88300 387796
rect 92020 387744 92072 387796
rect 93400 387744 93452 387796
rect 123576 387812 123628 387864
rect 125600 387812 125652 387864
rect 166632 387812 166684 387864
rect 167644 387812 167696 387864
rect 220176 387812 220228 387864
rect 221924 387812 221976 387864
rect 227628 387812 227680 387864
rect 228364 387812 228416 387864
rect 232504 387812 232556 387864
rect 234252 387812 234304 387864
rect 244924 387812 244976 387864
rect 245660 387812 245712 387864
rect 252008 387812 252060 387864
rect 253388 387812 253440 387864
rect 188344 387744 188396 387796
rect 218704 387744 218756 387796
rect 225788 387744 225840 387796
rect 260932 387744 260984 387796
rect 186780 387676 186832 387728
rect 211620 387676 211672 387728
rect 242900 387676 242952 387728
rect 266544 387676 266596 387728
rect 266728 387676 266780 387728
rect 219992 387268 220044 387320
rect 225788 387268 225840 387320
rect 240968 387200 241020 387252
rect 242900 387200 242952 387252
rect 100392 387064 100444 387116
rect 69020 386996 69072 387048
rect 69756 386996 69808 387048
rect 78680 386996 78732 387048
rect 79508 386996 79560 387048
rect 93860 386996 93912 387048
rect 94136 386996 94188 387048
rect 102140 386996 102192 387048
rect 102508 386996 102560 387048
rect 109040 386996 109092 387048
rect 109500 386996 109552 387048
rect 110696 387064 110748 387116
rect 188620 387064 188672 387116
rect 266728 387064 266780 387116
rect 272248 387064 272300 387116
rect 281448 387064 281500 387116
rect 582380 387064 582432 387116
rect 111064 386996 111116 387048
rect 155224 386452 155276 386504
rect 163504 386452 163556 386504
rect 84936 386316 84988 386368
rect 140044 386316 140096 386368
rect 186412 386316 186464 386368
rect 232504 386316 232556 386368
rect 245844 386316 245896 386368
rect 246948 386316 247000 386368
rect 262864 386316 262916 386368
rect 39948 386248 40000 386300
rect 88432 386248 88484 386300
rect 89260 386248 89312 386300
rect 107752 386248 107804 386300
rect 134616 386248 134668 386300
rect 135168 386248 135220 386300
rect 195428 386248 195480 386300
rect 197360 386248 197412 386300
rect 217324 386248 217376 386300
rect 218244 386248 218296 386300
rect 239496 386248 239548 386300
rect 253572 386248 253624 386300
rect 135168 385704 135220 385756
rect 163504 385704 163556 385756
rect 139400 385636 139452 385688
rect 189724 385636 189776 385688
rect 129740 384956 129792 385008
rect 130936 384956 130988 385008
rect 230572 384956 230624 385008
rect 231492 384956 231544 385008
rect 242164 384956 242216 385008
rect 271880 384956 271932 385008
rect 96896 384276 96948 384328
rect 116584 384276 116636 384328
rect 129740 384276 129792 384328
rect 3516 383664 3568 383716
rect 113456 383664 113508 383716
rect 228364 383664 228416 383716
rect 280344 383664 280396 383716
rect 111064 383596 111116 383648
rect 135904 383596 135956 383648
rect 177488 383596 177540 383648
rect 256884 383596 256936 383648
rect 87052 383324 87104 383376
rect 91284 383324 91336 383376
rect 135904 382984 135956 383036
rect 174268 382984 174320 383036
rect 65984 382916 66036 382968
rect 75184 382916 75236 382968
rect 78772 382916 78824 382968
rect 97264 382916 97316 382968
rect 97448 382916 97500 382968
rect 118700 382916 118752 382968
rect 231860 382916 231912 382968
rect 281724 382916 281776 382968
rect 182088 382168 182140 382220
rect 229100 382168 229152 382220
rect 181444 381692 181496 381744
rect 182088 381692 182140 381744
rect 102048 381556 102100 381608
rect 113364 381556 113416 381608
rect 214564 381556 214616 381608
rect 238760 381556 238812 381608
rect 77484 381488 77536 381540
rect 161388 381488 161440 381540
rect 169024 381488 169076 381540
rect 230572 381488 230624 381540
rect 277676 381488 277728 381540
rect 75276 380808 75328 380860
rect 161480 380808 161532 380860
rect 162216 380808 162268 380860
rect 188620 380808 188672 380860
rect 188988 380808 189040 380860
rect 250720 380808 250772 380860
rect 109132 380128 109184 380180
rect 129004 380128 129056 380180
rect 141424 380128 141476 380180
rect 187700 380128 187752 380180
rect 190276 380128 190328 380180
rect 265072 380128 265124 380180
rect 273352 380128 273404 380180
rect 82820 379448 82872 379500
rect 164884 379448 164936 379500
rect 189172 379448 189224 379500
rect 273536 379448 273588 379500
rect 187700 379380 187752 379432
rect 247684 379380 247736 379432
rect 273352 379244 273404 379296
rect 273536 379244 273588 379296
rect 104900 378768 104952 378820
rect 153936 378768 153988 378820
rect 252468 378768 252520 378820
rect 266544 378768 266596 378820
rect 72516 378088 72568 378140
rect 148416 378088 148468 378140
rect 161296 378088 161348 378140
rect 223580 378088 223632 378140
rect 224224 378088 224276 378140
rect 236644 378088 236696 378140
rect 264244 378088 264296 378140
rect 93952 377408 94004 377460
rect 120724 377408 120776 377460
rect 228364 377408 228416 377460
rect 151176 376660 151228 376712
rect 247132 376660 247184 376712
rect 77208 376592 77260 376644
rect 154488 376592 154540 376644
rect 75920 376048 75972 376100
rect 77208 376048 77260 376100
rect 46756 375980 46808 376032
rect 78680 375980 78732 376032
rect 108856 375980 108908 376032
rect 116032 375980 116084 376032
rect 65892 375300 65944 375352
rect 171876 375300 171928 375352
rect 172060 375300 172112 375352
rect 174268 375300 174320 375352
rect 236000 375300 236052 375352
rect 236644 375300 236696 375352
rect 279424 375300 279476 375352
rect 281540 375300 281592 375352
rect 236644 374688 236696 374740
rect 291384 374688 291436 374740
rect 88340 374620 88392 374672
rect 141516 374620 141568 374672
rect 142252 374620 142304 374672
rect 148324 374620 148376 374672
rect 241520 374620 241572 374672
rect 251824 374620 251876 374672
rect 163504 373940 163556 373992
rect 245752 373940 245804 373992
rect 77208 373328 77260 373380
rect 84292 373328 84344 373380
rect 107568 373328 107620 373380
rect 115940 373328 115992 373380
rect 153936 373328 153988 373380
rect 186412 373328 186464 373380
rect 244924 373328 244976 373380
rect 258724 373328 258776 373380
rect 74540 373260 74592 373312
rect 157340 373260 157392 373312
rect 191104 373260 191156 373312
rect 203524 373260 203576 373312
rect 251916 373260 251968 373312
rect 266636 373260 266688 373312
rect 117964 372580 118016 372632
rect 147496 372580 147548 372632
rect 147680 372580 147732 372632
rect 245752 372580 245804 372632
rect 246304 372580 246356 372632
rect 179052 372512 179104 372564
rect 227720 372512 227772 372564
rect 84108 372444 84160 372496
rect 180064 372444 180116 372496
rect 182916 372444 182968 372496
rect 222200 372444 222252 372496
rect 48228 371832 48280 371884
rect 75920 371832 75972 371884
rect 249708 371832 249760 371884
rect 269396 371832 269448 371884
rect 179420 371764 179472 371816
rect 180064 371764 180116 371816
rect 222200 371220 222252 371272
rect 222844 371220 222896 371272
rect 227720 371220 227772 371272
rect 228456 371220 228508 371272
rect 270408 371220 270460 371272
rect 274916 371220 274968 371272
rect 155684 371152 155736 371204
rect 240140 371152 240192 371204
rect 240876 371152 240928 371204
rect 247040 371152 247092 371204
rect 248328 371152 248380 371204
rect 295432 371152 295484 371204
rect 85580 371084 85632 371136
rect 160744 371084 160796 371136
rect 170404 371084 170456 371136
rect 234620 371084 234672 371136
rect 234620 370472 234672 370524
rect 244924 370472 244976 370524
rect 160100 370268 160152 370320
rect 160744 370268 160796 370320
rect 97264 369792 97316 369844
rect 129740 369792 129792 369844
rect 187700 369792 187752 369844
rect 242164 369792 242216 369844
rect 164884 369724 164936 369776
rect 213920 369724 213972 369776
rect 129740 369180 129792 369232
rect 130384 369180 130436 369232
rect 180064 369180 180116 369232
rect 71688 369112 71740 369164
rect 163964 369112 164016 369164
rect 165068 369112 165120 369164
rect 234528 369112 234580 369164
rect 259460 369112 259512 369164
rect 111064 368432 111116 368484
rect 113272 368432 113324 368484
rect 276112 368432 276164 368484
rect 71044 368364 71096 368416
rect 169760 368364 169812 368416
rect 228364 367752 228416 367804
rect 263692 367752 263744 367804
rect 67732 367004 67784 367056
rect 155960 367004 156012 367056
rect 157340 367004 157392 367056
rect 158444 367004 158496 367056
rect 201500 367004 201552 367056
rect 75184 366936 75236 366988
rect 137468 366936 137520 366988
rect 176108 366936 176160 366988
rect 176752 366936 176804 366988
rect 176752 366324 176804 366376
rect 254124 366324 254176 366376
rect 73252 365644 73304 365696
rect 167000 365644 167052 365696
rect 167644 365644 167696 365696
rect 186412 365644 186464 365696
rect 240968 365644 241020 365696
rect 248972 365644 249024 365696
rect 249800 365644 249852 365696
rect 57704 365576 57756 365628
rect 144184 365576 144236 365628
rect 163964 365576 164016 365628
rect 196072 365576 196124 365628
rect 196072 365168 196124 365220
rect 196624 365168 196676 365220
rect 242256 364964 242308 365016
rect 284484 364964 284536 365016
rect 69112 364284 69164 364336
rect 171140 364284 171192 364336
rect 171968 364284 172020 364336
rect 180064 364284 180116 364336
rect 180616 364284 180668 364336
rect 207020 364284 207072 364336
rect 123576 364216 123628 364268
rect 226340 364216 226392 364268
rect 228456 363672 228508 363724
rect 251824 363672 251876 363724
rect 260104 363672 260156 363724
rect 296720 363672 296772 363724
rect 226340 363604 226392 363656
rect 266636 363604 266688 363656
rect 111800 362856 111852 362908
rect 112536 362856 112588 362908
rect 252008 362856 252060 362908
rect 266636 362856 266688 362908
rect 293960 362856 294012 362908
rect 93860 362176 93912 362228
rect 110512 362176 110564 362228
rect 151084 362176 151136 362228
rect 216680 362176 216732 362228
rect 249616 361564 249668 361616
rect 274732 361564 274784 361616
rect 73160 361496 73212 361548
rect 140780 361496 140832 361548
rect 153844 361496 153896 361548
rect 270776 361496 270828 361548
rect 140780 360816 140832 360868
rect 142068 360816 142120 360868
rect 168380 360816 168432 360868
rect 69020 360136 69072 360188
rect 69664 360136 69716 360188
rect 197360 360136 197412 360188
rect 168380 360068 168432 360120
rect 169484 360068 169536 360120
rect 178868 360068 178920 360120
rect 206284 359456 206336 359508
rect 260840 359456 260892 359508
rect 3332 358708 3384 358760
rect 36544 358708 36596 358760
rect 145656 358708 145708 358760
rect 255320 358708 255372 358760
rect 100760 358028 100812 358080
rect 122840 358028 122892 358080
rect 123760 358028 123812 358080
rect 123760 357416 123812 357468
rect 239404 357416 239456 357468
rect 196624 356736 196676 356788
rect 240140 356736 240192 356788
rect 129004 356668 129056 356720
rect 168380 356668 168432 356720
rect 214656 356668 214708 356720
rect 229008 356668 229060 356720
rect 256792 356668 256844 356720
rect 75184 355988 75236 356040
rect 75828 355988 75880 356040
rect 191104 355988 191156 356040
rect 102232 355920 102284 355972
rect 103336 355920 103388 355972
rect 214564 355920 214616 355972
rect 213184 355376 213236 355428
rect 258172 355376 258224 355428
rect 214564 355308 214616 355360
rect 269212 355308 269264 355360
rect 102140 354628 102192 354680
rect 239496 354628 239548 354680
rect 244188 354016 244240 354068
rect 262404 354016 262456 354068
rect 213828 353948 213880 354000
rect 259552 353948 259604 354000
rect 153844 353268 153896 353320
rect 198740 353268 198792 353320
rect 147496 353200 147548 353252
rect 217324 353200 217376 353252
rect 108856 352520 108908 352572
rect 280436 352520 280488 352572
rect 108396 351908 108448 351960
rect 108856 351908 108908 351960
rect 162584 351160 162636 351212
rect 194600 351160 194652 351212
rect 216588 351160 216640 351212
rect 238116 351160 238168 351212
rect 84200 350548 84252 350600
rect 270684 350548 270736 350600
rect 270960 350548 271012 350600
rect 88248 350480 88300 350532
rect 220084 350480 220136 350532
rect 207664 349800 207716 349852
rect 235264 349800 235316 349852
rect 146944 348440 146996 348492
rect 188896 348440 188948 348492
rect 206376 348440 206428 348492
rect 209136 348440 209188 348492
rect 233884 348440 233936 348492
rect 106924 348304 106976 348356
rect 107568 348304 107620 348356
rect 278964 348372 279016 348424
rect 234436 347012 234488 347064
rect 267740 347012 267792 347064
rect 134616 346468 134668 346520
rect 214564 346468 214616 346520
rect 147128 346400 147180 346452
rect 290004 346400 290056 346452
rect 71964 345584 72016 345636
rect 73068 345584 73120 345636
rect 122104 345108 122156 345160
rect 217416 345108 217468 345160
rect 3332 345040 3384 345092
rect 35164 345040 35216 345092
rect 73068 345040 73120 345092
rect 292672 345040 292724 345092
rect 245016 344360 245068 344412
rect 253940 344360 253992 344412
rect 15200 344292 15252 344344
rect 150348 344292 150400 344344
rect 197360 344292 197412 344344
rect 198004 344292 198056 344344
rect 236644 344292 236696 344344
rect 250444 344292 250496 344344
rect 267740 344292 267792 344344
rect 44180 342864 44232 342916
rect 189172 342864 189224 342916
rect 206468 342864 206520 342916
rect 253940 342864 253992 342916
rect 124864 342524 124916 342576
rect 125508 342524 125560 342576
rect 125508 342252 125560 342304
rect 269396 342252 269448 342304
rect 177304 341504 177356 341556
rect 185032 341504 185084 341556
rect 67456 340892 67508 340944
rect 295616 340892 295668 340944
rect 215944 340144 215996 340196
rect 243084 340144 243136 340196
rect 116768 339532 116820 339584
rect 183560 339532 183612 339584
rect 184296 339532 184348 339584
rect 82728 339464 82780 339516
rect 220084 339464 220136 339516
rect 183284 339396 183336 339448
rect 186320 339396 186372 339448
rect 234344 339396 234396 339448
rect 234804 339396 234856 339448
rect 187608 338784 187660 338836
rect 251916 338784 251968 338836
rect 155224 338716 155276 338768
rect 234804 338716 234856 338768
rect 178040 337424 178092 337476
rect 237380 337424 237432 337476
rect 252008 337424 252060 337476
rect 261024 337424 261076 337476
rect 217324 337356 217376 337408
rect 294144 337356 294196 337408
rect 41420 336812 41472 336864
rect 178040 336812 178092 336864
rect 178132 336744 178184 336796
rect 212632 336744 212684 336796
rect 186136 335996 186188 336048
rect 244464 335996 244516 336048
rect 137376 335316 137428 335368
rect 245016 335316 245068 335368
rect 178592 334024 178644 334076
rect 230572 334024 230624 334076
rect 178868 333956 178920 334008
rect 242256 333956 242308 334008
rect 210424 333208 210476 333260
rect 274640 333208 274692 333260
rect 169024 332664 169076 332716
rect 200212 332664 200264 332716
rect 141608 332596 141660 332648
rect 247132 332596 247184 332648
rect 247684 332596 247736 332648
rect 219348 331916 219400 331968
rect 260104 331916 260156 331968
rect 141700 331848 141752 331900
rect 183376 331848 183428 331900
rect 236000 331848 236052 331900
rect 163504 331236 163556 331288
rect 191840 331236 191892 331288
rect 193036 331236 193088 331288
rect 127624 330488 127676 330540
rect 204168 330488 204220 330540
rect 246304 330488 246356 330540
rect 259460 330488 259512 330540
rect 264888 330488 264940 330540
rect 272156 330488 272208 330540
rect 205732 329876 205784 329928
rect 245660 329876 245712 329928
rect 166356 329808 166408 329860
rect 166724 329808 166776 329860
rect 258172 329808 258224 329860
rect 153016 329740 153068 329792
rect 157340 329740 157392 329792
rect 8300 329060 8352 329112
rect 153200 329060 153252 329112
rect 186228 329060 186280 329112
rect 187516 329060 187568 329112
rect 205732 329060 205784 329112
rect 233884 329060 233936 329112
rect 253204 329060 253256 329112
rect 157340 328448 157392 328500
rect 243176 328448 243228 328500
rect 193036 328176 193088 328228
rect 195980 328176 196032 328228
rect 96712 327700 96764 327752
rect 249892 327700 249944 327752
rect 241520 326408 241572 326460
rect 242348 326408 242400 326460
rect 251824 326408 251876 326460
rect 260840 326408 260892 326460
rect 33140 326340 33192 326392
rect 154028 326340 154080 326392
rect 184296 326340 184348 326392
rect 251916 326340 251968 326392
rect 155316 325660 155368 325712
rect 241520 325660 241572 325712
rect 280528 325660 280580 325712
rect 580908 325660 580960 325712
rect 153936 324980 153988 325032
rect 215300 324980 215352 325032
rect 256884 324980 256936 325032
rect 88984 324912 89036 324964
rect 166356 324912 166408 324964
rect 193128 324912 193180 324964
rect 255504 324912 255556 324964
rect 151084 323620 151136 323672
rect 162124 323620 162176 323672
rect 176016 323620 176068 323672
rect 204260 323620 204312 323672
rect 211804 323620 211856 323672
rect 246396 323620 246448 323672
rect 152556 323552 152608 323604
rect 183468 323552 183520 323604
rect 209780 323552 209832 323604
rect 220084 323552 220136 323604
rect 262220 323552 262272 323604
rect 115204 321648 115256 321700
rect 185676 321648 185728 321700
rect 155868 321580 155920 321632
rect 158812 321580 158864 321632
rect 263784 321580 263836 321632
rect 126888 321512 126940 321564
rect 281540 321512 281592 321564
rect 281540 321308 281592 321360
rect 281816 321308 281868 321360
rect 104256 320832 104308 320884
rect 125692 320832 125744 320884
rect 126888 320832 126940 320884
rect 106188 320152 106240 320204
rect 261024 320152 261076 320204
rect 251824 320084 251876 320136
rect 252008 320084 252060 320136
rect 4068 319404 4120 319456
rect 15844 319404 15896 319456
rect 188344 319404 188396 319456
rect 267924 319404 267976 319456
rect 181904 319064 181956 319116
rect 187056 319064 187108 319116
rect 162124 318792 162176 318844
rect 251824 318792 251876 318844
rect 182824 318044 182876 318096
rect 185032 318044 185084 318096
rect 233884 318044 233936 318096
rect 240876 318044 240928 318096
rect 256792 318044 256844 318096
rect 149980 317500 150032 317552
rect 182180 317500 182232 317552
rect 178684 317432 178736 317484
rect 236644 317432 236696 317484
rect 246304 317432 246356 317484
rect 250996 317432 251048 317484
rect 75276 317364 75328 317416
rect 81440 317364 81492 317416
rect 151636 316752 151688 316804
rect 169668 316752 169720 316804
rect 32404 316684 32456 316736
rect 159364 316684 159416 316736
rect 263600 316684 263652 316736
rect 169668 316004 169720 316056
rect 264980 316004 265032 316056
rect 89536 315256 89588 315308
rect 99472 315256 99524 315308
rect 256700 315256 256752 315308
rect 257436 315256 257488 315308
rect 295524 315256 295576 315308
rect 160744 314712 160796 314764
rect 256700 314712 256752 314764
rect 60648 314644 60700 314696
rect 263692 314644 263744 314696
rect 182180 313964 182232 314016
rect 247776 313964 247828 314016
rect 129096 313896 129148 313948
rect 260932 313896 260984 313948
rect 104440 313284 104492 313336
rect 124864 313284 124916 313336
rect 129096 313284 129148 313336
rect 249616 313284 249668 313336
rect 296720 313284 296772 313336
rect 104348 312604 104400 312656
rect 115204 312604 115256 312656
rect 242164 312604 242216 312656
rect 252744 312604 252796 312656
rect 73804 312536 73856 312588
rect 80244 312536 80296 312588
rect 108212 312536 108264 312588
rect 142160 312536 142212 312588
rect 262496 312536 262548 312588
rect 148416 311856 148468 311908
rect 217416 311856 217468 311908
rect 126336 311176 126388 311228
rect 149796 311312 149848 311364
rect 82912 311108 82964 311160
rect 147128 311108 147180 311160
rect 164976 311108 165028 311160
rect 173164 311108 173216 311160
rect 218060 311108 218112 311160
rect 239404 311108 239456 311160
rect 255412 311108 255464 311160
rect 155408 310496 155460 310548
rect 276296 310496 276348 310548
rect 97264 309816 97316 309868
rect 108212 309816 108264 309868
rect 163780 309816 163832 309868
rect 257344 309816 257396 309868
rect 259552 309816 259604 309868
rect 61752 309748 61804 309800
rect 166448 309748 166500 309800
rect 230480 309748 230532 309800
rect 252652 309748 252704 309800
rect 189080 309136 189132 309188
rect 190368 309136 190420 309188
rect 218704 309136 218756 309188
rect 178592 308456 178644 308508
rect 189080 308456 189132 308508
rect 99196 308388 99248 308440
rect 125508 308388 125560 308440
rect 131120 308388 131172 308440
rect 151176 308388 151228 308440
rect 157248 308388 157300 308440
rect 207572 308388 207624 308440
rect 224868 308388 224920 308440
rect 255596 308388 255648 308440
rect 189724 307776 189776 307828
rect 225972 307776 226024 307828
rect 239496 307776 239548 307828
rect 241428 307776 241480 307828
rect 138020 307708 138072 307760
rect 149980 307708 150032 307760
rect 173716 307708 173768 307760
rect 175280 307708 175332 307760
rect 196256 307708 196308 307760
rect 196716 307708 196768 307760
rect 71136 307096 71188 307148
rect 77392 307096 77444 307148
rect 122196 307096 122248 307148
rect 74632 307028 74684 307080
rect 138020 307028 138072 307080
rect 145564 307028 145616 307080
rect 176752 307164 176804 307216
rect 176016 307096 176068 307148
rect 176476 307096 176528 307148
rect 176752 307028 176804 307080
rect 196256 307028 196308 307080
rect 236644 307028 236696 307080
rect 267832 307028 267884 307080
rect 169484 306552 169536 306604
rect 172520 306552 172572 306604
rect 176016 306348 176068 306400
rect 259736 306348 259788 306400
rect 67364 305600 67416 305652
rect 88984 305600 89036 305652
rect 91192 305600 91244 305652
rect 104440 305600 104492 305652
rect 109040 305600 109092 305652
rect 118792 305600 118844 305652
rect 119344 305600 119396 305652
rect 144276 305600 144328 305652
rect 185676 305600 185728 305652
rect 193864 305600 193916 305652
rect 206376 305600 206428 305652
rect 215392 305600 215444 305652
rect 4068 305124 4120 305176
rect 7564 305124 7616 305176
rect 193588 305056 193640 305108
rect 228364 305056 228416 305108
rect 252468 305056 252520 305108
rect 258080 305056 258132 305108
rect 258724 305056 258776 305108
rect 80060 304988 80112 305040
rect 109040 304988 109092 305040
rect 144828 304988 144880 305040
rect 197452 304988 197504 305040
rect 253388 304988 253440 305040
rect 284484 304988 284536 305040
rect 223396 304920 223448 304972
rect 227628 304920 227680 304972
rect 229836 304920 229888 304972
rect 251916 304784 251968 304836
rect 258264 304784 258316 304836
rect 232228 304580 232280 304632
rect 240784 304580 240836 304632
rect 123576 304308 123628 304360
rect 144184 304308 144236 304360
rect 218428 304308 218480 304360
rect 219348 304308 219400 304360
rect 242440 304308 242492 304360
rect 252468 304308 252520 304360
rect 96620 304240 96672 304292
rect 147220 304240 147272 304292
rect 181444 304240 181496 304292
rect 229008 304240 229060 304292
rect 247776 304240 247828 304292
rect 258356 304240 258408 304292
rect 262680 304240 262732 304292
rect 298192 304240 298244 304292
rect 232504 303696 232556 303748
rect 233976 303696 234028 303748
rect 148324 303628 148376 303680
rect 213184 303628 213236 303680
rect 214564 303628 214616 303680
rect 217232 303628 217284 303680
rect 220912 303628 220964 303680
rect 221740 303628 221792 303680
rect 223580 303628 223632 303680
rect 224132 303628 224184 303680
rect 225052 303628 225104 303680
rect 226248 303628 226300 303680
rect 230572 303628 230624 303680
rect 231308 303628 231360 303680
rect 233884 303628 233936 303680
rect 234620 303628 234672 303680
rect 237380 303628 237432 303680
rect 237932 303628 237984 303680
rect 242256 303628 242308 303680
rect 244188 303628 244240 303680
rect 248696 303628 248748 303680
rect 249340 303628 249392 303680
rect 201592 303560 201644 303612
rect 202880 303560 202932 303612
rect 203708 303560 203760 303612
rect 204260 303560 204312 303612
rect 204812 303560 204864 303612
rect 201592 303356 201644 303408
rect 216588 303356 216640 303408
rect 218980 303356 219032 303408
rect 233424 303152 233476 303204
rect 234436 303152 234488 303204
rect 121460 302880 121512 302932
rect 216588 302880 216640 302932
rect 240600 302268 240652 302320
rect 262312 302268 262364 302320
rect 262680 302268 262732 302320
rect 73068 302200 73120 302252
rect 164976 302200 165028 302252
rect 187056 302200 187108 302252
rect 233424 302200 233476 302252
rect 231124 302132 231176 302184
rect 268108 302200 268160 302252
rect 258724 302132 258776 302184
rect 266360 302132 266412 302184
rect 86224 301520 86276 301572
rect 129188 301520 129240 301572
rect 242348 301520 242400 301572
rect 34520 301452 34572 301504
rect 179328 301452 179380 301504
rect 254124 301452 254176 301504
rect 244372 301384 244424 301436
rect 245108 301384 245160 301436
rect 193680 300908 193732 300960
rect 197636 300908 197688 300960
rect 166264 300840 166316 300892
rect 215668 301044 215720 301096
rect 211068 300976 211120 301028
rect 156604 300772 156656 300824
rect 160836 300772 160888 300824
rect 191104 300772 191156 300824
rect 129188 300160 129240 300212
rect 141700 300160 141752 300212
rect 190920 300160 190972 300212
rect 216864 300908 216916 300960
rect 227720 300908 227772 300960
rect 249248 300908 249300 300960
rect 258724 300908 258776 300960
rect 255320 300160 255372 300212
rect 274640 300160 274692 300212
rect 140228 300092 140280 300144
rect 193588 300092 193640 300144
rect 252468 300092 252520 300144
rect 254032 300092 254084 300144
rect 258724 300092 258776 300144
rect 282920 300092 282972 300144
rect 253020 299412 253072 299464
rect 272064 299412 272116 299464
rect 159548 298800 159600 298852
rect 188988 298800 189040 298852
rect 191748 298800 191800 298852
rect 138756 298732 138808 298784
rect 187700 298732 187752 298784
rect 256608 298120 256660 298172
rect 261484 298120 261536 298172
rect 304264 298120 304316 298172
rect 580172 298120 580224 298172
rect 168472 298052 168524 298104
rect 189724 298052 189776 298104
rect 122932 297372 122984 297424
rect 132408 297372 132460 297424
rect 184848 297372 184900 297424
rect 191748 297372 191800 297424
rect 88432 297168 88484 297220
rect 89536 297168 89588 297220
rect 89536 296692 89588 296744
rect 115388 296692 115440 296744
rect 255320 296692 255372 296744
rect 267924 296692 267976 296744
rect 256608 296012 256660 296064
rect 272064 296012 272116 296064
rect 161940 295944 161992 295996
rect 175188 295944 175240 295996
rect 185676 295944 185728 295996
rect 258540 295944 258592 295996
rect 288716 295944 288768 295996
rect 165528 295332 165580 295384
rect 168380 295332 168432 295384
rect 256608 295264 256660 295316
rect 267740 295264 267792 295316
rect 274824 295264 274876 295316
rect 155960 294652 156012 294704
rect 156604 294652 156656 294704
rect 137468 294584 137520 294636
rect 144736 294584 144788 294636
rect 175188 294584 175240 294636
rect 69664 293972 69716 294024
rect 155960 293972 156012 294024
rect 175188 293972 175240 294024
rect 191748 293972 191800 294024
rect 256332 293972 256384 294024
rect 290004 293972 290056 294024
rect 92572 293904 92624 293956
rect 93768 293904 93820 293956
rect 122932 293904 122984 293956
rect 261576 293904 261628 293956
rect 262220 293904 262272 293956
rect 261484 293836 261536 293888
rect 302332 293904 302384 293956
rect 255964 293224 256016 293276
rect 258816 293224 258868 293276
rect 256148 293088 256200 293140
rect 260748 293088 260800 293140
rect 168380 292612 168432 292664
rect 169116 292612 169168 292664
rect 191564 292612 191616 292664
rect 3516 292544 3568 292596
rect 22836 292544 22888 292596
rect 84568 292544 84620 292596
rect 177856 292544 177908 292596
rect 184756 292544 184808 292596
rect 188712 292544 188764 292596
rect 99288 292476 99340 292528
rect 157156 292476 157208 292528
rect 168380 292476 168432 292528
rect 255964 292136 256016 292188
rect 256884 292136 256936 292188
rect 258632 292136 258684 292188
rect 177856 292068 177908 292120
rect 178868 292068 178920 292120
rect 178960 291864 179012 291916
rect 188344 291864 188396 291916
rect 60464 291796 60516 291848
rect 75184 291796 75236 291848
rect 151360 291796 151412 291848
rect 189816 291796 189868 291848
rect 257344 291796 257396 291848
rect 261024 291796 261076 291848
rect 98368 291252 98420 291304
rect 99288 291252 99340 291304
rect 89536 291184 89588 291236
rect 121552 291184 121604 291236
rect 255504 290980 255556 291032
rect 258172 290980 258224 291032
rect 71872 290436 71924 290488
rect 161940 290436 161992 290488
rect 188712 290028 188764 290080
rect 188988 290028 189040 290080
rect 191196 290028 191248 290080
rect 162216 289824 162268 289876
rect 191656 289824 191708 289876
rect 162768 289756 162820 289808
rect 191748 289756 191800 289808
rect 260748 289756 260800 289808
rect 269212 289756 269264 289808
rect 255504 289688 255556 289740
rect 262496 289688 262548 289740
rect 76196 289416 76248 289468
rect 76564 289416 76616 289468
rect 64788 289076 64840 289128
rect 151084 289076 151136 289128
rect 159456 289076 159508 289128
rect 162768 289076 162820 289128
rect 45468 288396 45520 288448
rect 76196 288396 76248 288448
rect 79232 288396 79284 288448
rect 79968 288396 80020 288448
rect 159456 288396 159508 288448
rect 35164 288328 35216 288380
rect 70584 288328 70636 288380
rect 71044 288328 71096 288380
rect 255504 288328 255556 288380
rect 281540 288328 281592 288380
rect 255320 288260 255372 288312
rect 263784 288260 263836 288312
rect 74632 287784 74684 287836
rect 75368 287784 75420 287836
rect 92480 287784 92532 287836
rect 92940 287784 92992 287836
rect 68284 287716 68336 287768
rect 158812 287716 158864 287768
rect 78588 287648 78640 287700
rect 184204 287648 184256 287700
rect 182916 287512 182968 287564
rect 190184 287512 190236 287564
rect 170496 286968 170548 287020
rect 191748 286968 191800 287020
rect 255412 286628 255464 286680
rect 257344 286628 257396 286680
rect 80428 286424 80480 286476
rect 81256 286424 81308 286476
rect 83464 286424 83516 286476
rect 144184 286288 144236 286340
rect 187056 286288 187108 286340
rect 255504 286288 255556 286340
rect 258356 286288 258408 286340
rect 260840 286288 260892 286340
rect 81992 286084 82044 286136
rect 82728 286084 82780 286136
rect 84660 286084 84712 286136
rect 95332 286084 95384 286136
rect 97264 286084 97316 286136
rect 52184 285744 52236 285796
rect 69020 285812 69072 285864
rect 73804 285812 73856 285864
rect 53564 285676 53616 285728
rect 69020 285676 69072 285728
rect 72424 285676 72476 285728
rect 87512 285676 87564 285728
rect 90364 285676 90416 285728
rect 90824 285676 90876 285728
rect 118056 285676 118108 285728
rect 167644 285676 167696 285728
rect 170496 285676 170548 285728
rect 255412 285608 255464 285660
rect 260932 285608 260984 285660
rect 54300 284928 54352 284980
rect 87604 284928 87656 284980
rect 176568 284928 176620 284980
rect 185584 284928 185636 284980
rect 91100 284384 91152 284436
rect 98460 284384 98512 284436
rect 37924 284316 37976 284368
rect 54300 284316 54352 284368
rect 54852 284316 54904 284368
rect 58900 284316 58952 284368
rect 71872 284316 71924 284368
rect 88156 284316 88208 284368
rect 99380 284316 99432 284368
rect 128268 284316 128320 284368
rect 191748 284316 191800 284368
rect 266544 284316 266596 284368
rect 266728 284316 266780 284368
rect 255412 284248 255464 284300
rect 295616 284248 295668 284300
rect 169668 284112 169720 284164
rect 169944 284112 169996 284164
rect 86086 283704 86138 283756
rect 86868 283704 86920 283756
rect 52368 283568 52420 283620
rect 56416 283568 56468 283620
rect 66260 283568 66312 283620
rect 162768 283568 162820 283620
rect 176016 283568 176068 283620
rect 88616 283364 88668 283416
rect 88984 283364 89036 283416
rect 98092 283364 98144 283416
rect 98368 283364 98420 283416
rect 255504 283364 255556 283416
rect 259736 283364 259788 283416
rect 68652 283228 68704 283280
rect 69388 283228 69440 283280
rect 70308 283228 70360 283280
rect 83556 283228 83608 283280
rect 84016 283228 84068 283280
rect 67548 283024 67600 283076
rect 69020 282684 69072 282736
rect 69664 282956 69716 283008
rect 158720 282956 158772 283008
rect 68928 282616 68980 282668
rect 162768 282888 162820 282940
rect 175924 282888 175976 282940
rect 180156 282888 180208 282940
rect 191748 282888 191800 282940
rect 98460 282820 98512 282872
rect 163780 282820 163832 282872
rect 255504 282820 255556 282872
rect 263600 282820 263652 282872
rect 68560 282140 68612 282192
rect 98920 282140 98972 282192
rect 169024 282140 169076 282192
rect 182824 282140 182876 282192
rect 259276 282140 259328 282192
rect 267832 282140 267884 282192
rect 273444 282140 273496 282192
rect 291384 282140 291436 282192
rect 255412 281936 255464 281988
rect 259368 281936 259420 281988
rect 184296 281596 184348 281648
rect 192024 281596 192076 281648
rect 100760 281528 100812 281580
rect 108488 281528 108540 281580
rect 155500 281528 155552 281580
rect 191748 281528 191800 281580
rect 100852 281460 100904 281512
rect 103428 281460 103480 281512
rect 107568 281460 107620 281512
rect 255504 281460 255556 281512
rect 276112 281460 276164 281512
rect 255412 281392 255464 281444
rect 263692 281392 263744 281444
rect 160836 280780 160888 280832
rect 161388 280780 161440 280832
rect 191748 280780 191800 280832
rect 175924 280644 175976 280696
rect 178776 280644 178828 280696
rect 43444 280168 43496 280220
rect 66720 280168 66772 280220
rect 68928 280168 68980 280220
rect 107016 280168 107068 280220
rect 114468 280168 114520 280220
rect 114652 280168 114704 280220
rect 263600 280168 263652 280220
rect 264244 280168 264296 280220
rect 292580 280168 292632 280220
rect 100760 280100 100812 280152
rect 130476 280100 130528 280152
rect 255504 280100 255556 280152
rect 269396 280100 269448 280152
rect 7564 279420 7616 279472
rect 35808 279420 35860 279472
rect 60648 279420 60700 279472
rect 66812 279420 66864 279472
rect 123484 279420 123536 279472
rect 153936 279420 153988 279472
rect 158720 278740 158772 278792
rect 160192 278740 160244 278792
rect 191748 278740 191800 278792
rect 255412 278672 255464 278724
rect 280344 278672 280396 278724
rect 255504 278604 255556 278656
rect 263600 278604 263652 278656
rect 65892 278264 65944 278316
rect 67548 278264 67600 278316
rect 99380 277992 99432 278044
rect 118884 277992 118936 278044
rect 138664 277992 138716 278044
rect 158444 277992 158496 278044
rect 183376 277992 183428 278044
rect 183376 277380 183428 277432
rect 191564 277380 191616 277432
rect 52276 277312 52328 277364
rect 66904 277312 66956 277364
rect 100208 277312 100260 277364
rect 184664 277312 184716 277364
rect 255596 277312 255648 277364
rect 278964 277312 279016 277364
rect 255412 276632 255464 276684
rect 276296 276632 276348 276684
rect 184664 276088 184716 276140
rect 189816 276088 189868 276140
rect 100760 276020 100812 276072
rect 129096 276020 129148 276072
rect 151268 276020 151320 276072
rect 191748 276020 191800 276072
rect 276112 276020 276164 276072
rect 276296 276020 276348 276072
rect 61844 275952 61896 276004
rect 66904 275952 66956 276004
rect 255504 275952 255556 276004
rect 277676 275952 277728 276004
rect 100944 275272 100996 275324
rect 155408 275272 155460 275324
rect 177948 275272 178000 275324
rect 184204 275272 184256 275324
rect 100760 274660 100812 274712
rect 136088 274660 136140 274712
rect 255412 274660 255464 274712
rect 270684 274660 270736 274712
rect 272248 274660 272300 274712
rect 100852 274592 100904 274644
rect 160744 274592 160796 274644
rect 163596 274592 163648 274644
rect 182916 274592 182968 274644
rect 255504 274592 255556 274644
rect 281724 274592 281776 274644
rect 255412 274252 255464 274304
rect 259552 274252 259604 274304
rect 60648 273232 60700 273284
rect 63316 273232 63368 273284
rect 66904 273232 66956 273284
rect 67272 273232 67324 273284
rect 68284 273232 68336 273284
rect 156696 273232 156748 273284
rect 160836 273232 160888 273284
rect 162768 273232 162820 273284
rect 163596 273232 163648 273284
rect 185584 273232 185636 273284
rect 188896 273232 188948 273284
rect 191748 273232 191800 273284
rect 100852 273164 100904 273216
rect 107016 273164 107068 273216
rect 255412 273164 255464 273216
rect 259460 273164 259512 273216
rect 291292 273164 291344 273216
rect 580172 273164 580224 273216
rect 135996 272552 136048 272604
rect 155224 272552 155276 272604
rect 100760 272484 100812 272536
rect 113180 272484 113232 272536
rect 141700 272484 141752 272536
rect 282000 272484 282052 272536
rect 290096 272484 290148 272536
rect 60556 271940 60608 271992
rect 61752 271940 61804 271992
rect 66904 271940 66956 271992
rect 136548 271804 136600 271856
rect 160100 271804 160152 271856
rect 191288 271872 191340 271924
rect 255412 271872 255464 271924
rect 281724 271872 281776 271924
rect 282000 271872 282052 271924
rect 158628 271736 158680 271788
rect 161480 271736 161532 271788
rect 184296 271804 184348 271856
rect 255504 271804 255556 271856
rect 261576 271804 261628 271856
rect 100760 271192 100812 271244
rect 114560 271192 114612 271244
rect 101220 271124 101272 271176
rect 102048 271124 102100 271176
rect 133696 271124 133748 271176
rect 259368 271124 259420 271176
rect 280436 271124 280488 271176
rect 184388 270648 184440 270700
rect 186228 270648 186280 270700
rect 191748 270648 191800 270700
rect 64696 270580 64748 270632
rect 66904 270580 66956 270632
rect 56508 270444 56560 270496
rect 59084 270444 59136 270496
rect 133696 270444 133748 270496
rect 151360 270444 151412 270496
rect 162124 270444 162176 270496
rect 169576 270444 169628 270496
rect 191196 270444 191248 270496
rect 255412 270240 255464 270292
rect 259368 270240 259420 270292
rect 41328 269764 41380 269816
rect 50804 269764 50856 269816
rect 59084 269764 59136 269816
rect 66904 269764 66956 269816
rect 98828 269764 98880 269816
rect 159640 269764 159692 269816
rect 261024 269764 261076 269816
rect 273260 269764 273312 269816
rect 255412 269152 255464 269204
rect 261024 269152 261076 269204
rect 100760 269084 100812 269136
rect 115480 269084 115532 269136
rect 178776 269084 178828 269136
rect 193404 269084 193456 269136
rect 259368 269084 259420 269136
rect 291292 269084 291344 269136
rect 52276 269016 52328 269068
rect 53748 269016 53800 269068
rect 66720 269016 66772 269068
rect 166264 269016 166316 269068
rect 167736 269016 167788 269068
rect 267832 269016 267884 269068
rect 270776 269016 270828 269068
rect 100024 268336 100076 268388
rect 115296 268336 115348 268388
rect 120816 268336 120868 268388
rect 133144 268336 133196 268388
rect 181904 268336 181956 268388
rect 192576 268336 192628 268388
rect 255412 268336 255464 268388
rect 271144 268336 271196 268388
rect 271788 268336 271840 268388
rect 99012 267996 99064 268048
rect 104256 267996 104308 268048
rect 255412 267724 255464 267776
rect 267832 267724 267884 267776
rect 271788 267724 271840 267776
rect 280436 267724 280488 267776
rect 3516 267656 3568 267708
rect 37924 267656 37976 267708
rect 50988 267656 51040 267708
rect 60740 267656 60792 267708
rect 98736 267656 98788 267708
rect 146208 267656 146260 267708
rect 100760 267044 100812 267096
rect 106096 267044 106148 267096
rect 146208 267044 146260 267096
rect 177396 267044 177448 267096
rect 118056 266976 118108 267028
rect 182916 266976 182968 267028
rect 265624 266976 265676 267028
rect 277492 266976 277544 267028
rect 62028 266364 62080 266416
rect 64604 266364 64656 266416
rect 66904 266364 66956 266416
rect 106188 266364 106240 266416
rect 112536 266364 112588 266416
rect 255412 266364 255464 266416
rect 258356 266364 258408 266416
rect 270408 266364 270460 266416
rect 270776 266364 270828 266416
rect 100760 265616 100812 265668
rect 148600 265616 148652 265668
rect 163596 265616 163648 265668
rect 191564 265616 191616 265668
rect 255320 265616 255372 265668
rect 265072 265616 265124 265668
rect 63408 264936 63460 264988
rect 66260 264936 66312 264988
rect 105636 264936 105688 264988
rect 109684 264936 109736 264988
rect 170312 264936 170364 264988
rect 191748 264936 191800 264988
rect 253848 264936 253900 264988
rect 273260 264936 273312 264988
rect 3424 264868 3476 264920
rect 32404 264868 32456 264920
rect 104440 264188 104492 264240
rect 173348 264188 173400 264240
rect 255412 264188 255464 264240
rect 184756 264120 184808 264172
rect 191748 264120 191800 264172
rect 263784 264052 263836 264104
rect 264336 264052 264388 264104
rect 60556 263848 60608 263900
rect 61660 263848 61712 263900
rect 66260 263848 66312 263900
rect 100760 263576 100812 263628
rect 113824 263576 113876 263628
rect 255504 263576 255556 263628
rect 259736 263576 259788 263628
rect 100668 263508 100720 263560
rect 113088 263508 113140 263560
rect 155500 263508 155552 263560
rect 255412 263508 255464 263560
rect 274732 263508 274784 263560
rect 277400 263508 277452 263560
rect 255504 262828 255556 262880
rect 287244 262828 287296 262880
rect 7564 262216 7616 262268
rect 49516 262216 49568 262268
rect 66260 262216 66312 262268
rect 99288 262148 99340 262200
rect 104348 262148 104400 262200
rect 133788 262080 133840 262132
rect 164240 262080 164292 262132
rect 191748 262216 191800 262268
rect 165528 262012 165580 262064
rect 191564 262148 191616 262200
rect 104808 261944 104860 261996
rect 110604 261944 110656 261996
rect 50896 261536 50948 261588
rect 66260 261536 66312 261588
rect 4068 261468 4120 261520
rect 66168 261468 66220 261520
rect 111800 261468 111852 261520
rect 129188 261468 129240 261520
rect 149888 261468 149940 261520
rect 166264 261468 166316 261520
rect 255504 261468 255556 261520
rect 278320 261468 278372 261520
rect 266452 260788 266504 260840
rect 279424 260788 279476 260840
rect 188988 260176 189040 260228
rect 193220 260176 193272 260228
rect 43996 260108 44048 260160
rect 66260 260108 66312 260160
rect 173256 260108 173308 260160
rect 191748 260108 191800 260160
rect 255412 260108 255464 260160
rect 266452 260108 266504 260160
rect 100760 259496 100812 259548
rect 137560 259496 137612 259548
rect 100852 259428 100904 259480
rect 163780 259428 163832 259480
rect 255412 259428 255464 259480
rect 263600 259428 263652 259480
rect 61936 259360 61988 259412
rect 66628 259360 66680 259412
rect 255596 259360 255648 259412
rect 294144 259360 294196 259412
rect 55128 258680 55180 258732
rect 58992 258680 59044 258732
rect 66352 258680 66404 258732
rect 100760 258680 100812 258732
rect 155316 258680 155368 258732
rect 255504 258680 255556 258732
rect 266452 258680 266504 258732
rect 285956 258068 286008 258120
rect 287336 258068 287388 258120
rect 66352 258000 66404 258052
rect 68192 258000 68244 258052
rect 101680 258000 101732 258052
rect 111064 258000 111116 258052
rect 44088 257320 44140 257372
rect 53840 257320 53892 257372
rect 102048 257320 102100 257372
rect 126428 257320 126480 257372
rect 136088 257320 136140 257372
rect 178868 257320 178920 257372
rect 255412 256776 255464 256828
rect 262588 256776 262640 256828
rect 262772 256776 262824 256828
rect 53840 256708 53892 256760
rect 54944 256708 54996 256760
rect 66260 256708 66312 256760
rect 174544 256640 174596 256692
rect 183468 256640 183520 256692
rect 190644 256640 190696 256692
rect 49608 255960 49660 256012
rect 64604 255960 64656 256012
rect 66904 255960 66956 256012
rect 100852 255960 100904 256012
rect 137376 255960 137428 256012
rect 283104 255960 283156 256012
rect 580724 255960 580776 256012
rect 255412 255348 255464 255400
rect 278964 255348 279016 255400
rect 100760 255280 100812 255332
rect 188528 255280 188580 255332
rect 254584 255280 254636 255332
rect 255596 255280 255648 255332
rect 283104 255280 283156 255332
rect 3424 255212 3476 255264
rect 43444 255212 43496 255264
rect 57888 254668 57940 254720
rect 66904 254668 66956 254720
rect 272340 254600 272392 254652
rect 280252 254600 280304 254652
rect 46848 254532 46900 254584
rect 66720 254532 66772 254584
rect 126888 254532 126940 254584
rect 162216 254532 162268 254584
rect 255412 254532 255464 254584
rect 285956 254532 286008 254584
rect 100760 253988 100812 254040
rect 111064 253988 111116 254040
rect 167828 253988 167880 254040
rect 170772 253988 170824 254040
rect 184296 253988 184348 254040
rect 56600 253920 56652 253972
rect 57888 253920 57940 253972
rect 102968 253920 103020 253972
rect 103336 253920 103388 253972
rect 125600 253920 125652 253972
rect 126888 253920 126940 253972
rect 190644 253920 190696 253972
rect 255504 253920 255556 253972
rect 271880 253920 271932 253972
rect 272340 253920 272392 253972
rect 63224 253852 63276 253904
rect 66628 253852 66680 253904
rect 131028 253852 131080 253904
rect 161480 253852 161532 253904
rect 163688 253240 163740 253292
rect 174636 253240 174688 253292
rect 32404 253172 32456 253224
rect 66904 253172 66956 253224
rect 67272 253172 67324 253224
rect 102876 253172 102928 253224
rect 173808 253172 173860 253224
rect 174728 253172 174780 253224
rect 179328 253172 179380 253224
rect 192668 253172 192720 253224
rect 255412 253172 255464 253224
rect 262496 253172 262548 253224
rect 281632 252764 281684 252816
rect 285864 252764 285916 252816
rect 101588 252492 101640 252544
rect 104808 252492 104860 252544
rect 128268 252492 128320 252544
rect 129740 252492 129792 252544
rect 255504 251880 255556 251932
rect 266452 251880 266504 251932
rect 55036 251812 55088 251864
rect 66076 251812 66128 251864
rect 66628 251812 66680 251864
rect 164148 251812 164200 251864
rect 191748 251812 191800 251864
rect 255412 251812 255464 251864
rect 281632 251812 281684 251864
rect 64880 251132 64932 251184
rect 66260 251132 66312 251184
rect 106096 251132 106148 251184
rect 106924 251132 106976 251184
rect 169576 251132 169628 251184
rect 191564 251132 191616 251184
rect 48136 250452 48188 250504
rect 66996 250452 67048 250504
rect 100760 250452 100812 250504
rect 106096 250452 106148 250504
rect 122196 250452 122248 250504
rect 167828 250452 167880 250504
rect 274916 250452 274968 250504
rect 582656 250452 582708 250504
rect 255504 249772 255556 249824
rect 274916 249772 274968 249824
rect 165528 249568 165580 249620
rect 168380 249568 168432 249620
rect 53656 249024 53708 249076
rect 64788 249024 64840 249076
rect 66904 249024 66956 249076
rect 100852 249024 100904 249076
rect 106188 249024 106240 249076
rect 129188 249024 129240 249076
rect 151268 249092 151320 249144
rect 137468 249024 137520 249076
rect 160284 249024 160336 249076
rect 182824 249024 182876 249076
rect 191656 249024 191708 249076
rect 187516 248820 187568 248872
rect 191288 248820 191340 248872
rect 255412 248480 255464 248532
rect 278044 248480 278096 248532
rect 255504 248412 255556 248464
rect 292672 248412 292724 248464
rect 582472 248412 582524 248464
rect 148600 247664 148652 247716
rect 180340 247664 180392 247716
rect 255504 247664 255556 247716
rect 259552 247664 259604 247716
rect 271972 247664 272024 247716
rect 53656 247052 53708 247104
rect 66628 247052 66680 247104
rect 181536 247052 181588 247104
rect 191748 247052 191800 247104
rect 254124 247052 254176 247104
rect 259644 247052 259696 247104
rect 59176 246984 59228 247036
rect 64880 246984 64932 247036
rect 101036 246304 101088 246356
rect 101404 246304 101456 246356
rect 159548 246304 159600 246356
rect 183376 246304 183428 246356
rect 192484 246304 192536 246356
rect 280068 246304 280120 246356
rect 298376 246304 298428 246356
rect 254676 246168 254728 246220
rect 258356 246168 258408 246220
rect 166356 245624 166408 245676
rect 169852 245624 169904 245676
rect 255688 245624 255740 245676
rect 279424 245624 279476 245676
rect 280068 245624 280120 245676
rect 100944 245556 100996 245608
rect 165620 245556 165672 245608
rect 255504 245556 255556 245608
rect 289820 245556 289872 245608
rect 100852 245148 100904 245200
rect 105636 245148 105688 245200
rect 184204 244944 184256 244996
rect 193680 244944 193732 244996
rect 165620 244876 165672 244928
rect 193128 244876 193180 244928
rect 255596 244876 255648 244928
rect 258540 244876 258592 244928
rect 284300 244876 284352 244928
rect 289820 244264 289872 244316
rect 294052 244264 294104 244316
rect 57704 244196 57756 244248
rect 66904 244196 66956 244248
rect 98552 243516 98604 243568
rect 106280 243516 106332 243568
rect 106924 243516 106976 243568
rect 125048 243516 125100 243568
rect 153844 243516 153896 243568
rect 189080 243516 189132 243568
rect 255504 243516 255556 243568
rect 277492 243516 277544 243568
rect 280252 243516 280304 243568
rect 100852 243448 100904 243500
rect 102784 243448 102836 243500
rect 185676 243448 185728 243500
rect 173808 243176 173860 243228
rect 176660 243176 176712 243228
rect 57704 242904 57756 242956
rect 66536 242904 66588 242956
rect 189080 242904 189132 242956
rect 191748 242904 191800 242956
rect 141700 242836 141752 242888
rect 184848 242836 184900 242888
rect 191104 242836 191156 242888
rect 186320 242768 186372 242820
rect 100852 242224 100904 242276
rect 103612 242224 103664 242276
rect 186320 242224 186372 242276
rect 187608 242224 187660 242276
rect 193588 242224 193640 242276
rect 69020 242156 69072 242208
rect 98184 242156 98236 242208
rect 258172 243448 258224 243500
rect 255688 242836 255740 242888
rect 258356 242836 258408 242888
rect 259276 242836 259328 242888
rect 252376 242292 252428 242344
rect 252928 242292 252980 242344
rect 259276 242224 259328 242276
rect 278780 242224 278832 242276
rect 255504 242156 255556 242208
rect 284392 242156 284444 242208
rect 192668 242020 192720 242072
rect 198004 242020 198056 242072
rect 198096 242020 198148 242072
rect 242992 242020 243044 242072
rect 95424 241748 95476 241800
rect 102968 241748 103020 241800
rect 57888 241476 57940 241528
rect 66904 241476 66956 241528
rect 193680 241476 193732 241528
rect 215300 241476 215352 241528
rect 216312 241476 216364 241528
rect 22836 241408 22888 241460
rect 93446 241408 93498 241460
rect 255596 241408 255648 241460
rect 268108 241408 268160 241460
rect 283012 241408 283064 241460
rect 3424 241068 3476 241120
rect 7564 241068 7616 241120
rect 94044 240796 94096 240848
rect 126980 240796 127032 240848
rect 110604 240728 110656 240780
rect 180708 240728 180760 240780
rect 193128 240728 193180 240780
rect 207296 240728 207348 240780
rect 250444 240728 250496 240780
rect 266636 240728 266688 240780
rect 68652 240592 68704 240644
rect 76656 240592 76708 240644
rect 249064 240592 249116 240644
rect 254124 240592 254176 240644
rect 69020 240116 69072 240168
rect 69940 240116 69992 240168
rect 73160 240116 73212 240168
rect 73804 240116 73856 240168
rect 74540 240116 74592 240168
rect 75460 240116 75512 240168
rect 78680 240116 78732 240168
rect 79324 240116 79376 240168
rect 89720 240116 89772 240168
rect 90364 240116 90416 240168
rect 126980 240116 127032 240168
rect 225604 240116 225656 240168
rect 48228 240048 48280 240100
rect 76012 240048 76064 240100
rect 76564 240048 76616 240100
rect 78220 240048 78272 240100
rect 80980 240048 81032 240100
rect 81808 240048 81860 240100
rect 182088 240048 182140 240100
rect 211528 240048 211580 240100
rect 213184 240048 213236 240100
rect 70492 239980 70544 240032
rect 71320 239980 71372 240032
rect 98552 239980 98604 240032
rect 166908 239980 166960 240032
rect 195336 239980 195388 240032
rect 89628 239912 89680 239964
rect 182088 239912 182140 239964
rect 71780 239776 71832 239828
rect 72700 239776 72752 239828
rect 75184 239640 75236 239692
rect 77300 239640 77352 239692
rect 82636 239504 82688 239556
rect 88432 239504 88484 239556
rect 83648 239436 83700 239488
rect 91008 239436 91060 239488
rect 224224 239368 224276 239420
rect 235540 239368 235592 239420
rect 252468 239368 252520 239420
rect 261484 239368 261536 239420
rect 91284 239300 91336 239352
rect 93952 239300 94004 239352
rect 252100 239164 252152 239216
rect 254032 239164 254084 239216
rect 224868 238960 224920 239012
rect 225972 238960 226024 239012
rect 84936 238756 84988 238808
rect 85488 238756 85540 238808
rect 46756 238688 46808 238740
rect 75000 238688 75052 238740
rect 160008 238688 160060 238740
rect 261024 238688 261076 238740
rect 80796 238620 80848 238672
rect 164884 238620 164936 238672
rect 222108 238620 222160 238672
rect 270776 238620 270828 238672
rect 193772 238484 193824 238536
rect 201500 238348 201552 238400
rect 201960 238348 202012 238400
rect 93860 238008 93912 238060
rect 113180 238008 113232 238060
rect 122840 238008 122892 238060
rect 68560 237940 68612 237992
rect 76748 237940 76800 237992
rect 221096 237668 221148 237720
rect 222108 237668 222160 237720
rect 78588 237396 78640 237448
rect 78772 237396 78824 237448
rect 67824 237328 67876 237380
rect 166356 237328 166408 237380
rect 193680 237328 193732 237380
rect 213920 237328 213972 237380
rect 164884 237260 164936 237312
rect 196624 237260 196676 237312
rect 86960 237124 87012 237176
rect 87604 237124 87656 237176
rect 196624 236716 196676 236768
rect 197176 236716 197228 236768
rect 214656 236716 214708 236768
rect 252376 236716 252428 236768
rect 50988 236648 51040 236700
rect 71872 236648 71924 236700
rect 93952 236648 94004 236700
rect 116676 236648 116728 236700
rect 118700 236648 118752 236700
rect 197360 236648 197412 236700
rect 259736 236648 259788 236700
rect 118976 236240 119028 236292
rect 124956 236240 125008 236292
rect 89536 235968 89588 236020
rect 89812 235968 89864 236020
rect 213920 235968 213972 236020
rect 214564 235968 214616 236020
rect 89352 235900 89404 235952
rect 110512 235900 110564 235952
rect 115480 235900 115532 235952
rect 259552 235900 259604 235952
rect 259828 235900 259880 235952
rect 182916 235832 182968 235884
rect 265256 235832 265308 235884
rect 280160 235220 280212 235272
rect 580264 235220 580316 235272
rect 182916 235016 182968 235068
rect 183468 235016 183520 235068
rect 43444 234608 43496 234660
rect 96896 234608 96948 234660
rect 97356 234608 97408 234660
rect 97908 234608 97960 234660
rect 99472 234608 99524 234660
rect 88340 234540 88392 234592
rect 120724 234540 120776 234592
rect 122932 234540 122984 234592
rect 167736 234540 167788 234592
rect 256792 234540 256844 234592
rect 137836 234472 137888 234524
rect 181536 234472 181588 234524
rect 192576 234472 192628 234524
rect 205640 234472 205692 234524
rect 207664 234472 207716 234524
rect 266544 234472 266596 234524
rect 205640 234064 205692 234116
rect 206744 234064 206796 234116
rect 97264 233860 97316 233912
rect 98092 233860 98144 233912
rect 69112 233180 69164 233232
rect 171048 233180 171100 233232
rect 207296 233180 207348 233232
rect 237380 233180 237432 233232
rect 237932 233180 237984 233232
rect 54852 233112 54904 233164
rect 87052 233112 87104 233164
rect 88248 233112 88300 233164
rect 89720 233112 89772 233164
rect 116584 233112 116636 233164
rect 122196 233112 122248 233164
rect 247684 232568 247736 232620
rect 262312 232568 262364 232620
rect 242164 232500 242216 232552
rect 268016 232500 268068 232552
rect 278044 232500 278096 232552
rect 580172 232500 580224 232552
rect 85488 231752 85540 231804
rect 140872 231752 140924 231804
rect 141516 231752 141568 231804
rect 171048 231752 171100 231804
rect 209136 231752 209188 231804
rect 225604 231752 225656 231804
rect 292580 231752 292632 231804
rect 80060 231072 80112 231124
rect 114652 231072 114704 231124
rect 123484 231072 123536 231124
rect 140872 231072 140924 231124
rect 178868 231072 178920 231124
rect 246304 231072 246356 231124
rect 267924 231072 267976 231124
rect 78680 230392 78732 230444
rect 108948 230392 109000 230444
rect 111892 230392 111944 230444
rect 163780 230392 163832 230444
rect 262404 230392 262456 230444
rect 268384 229984 268436 230036
rect 272064 229984 272116 230036
rect 74540 229712 74592 229764
rect 87604 229712 87656 229764
rect 88248 229712 88300 229764
rect 103520 229712 103572 229764
rect 111064 229712 111116 229764
rect 119344 229712 119396 229764
rect 152648 229712 152700 229764
rect 219440 229712 219492 229764
rect 258356 229712 258408 229764
rect 278688 229576 278740 229628
rect 284484 229576 284536 229628
rect 178868 229032 178920 229084
rect 214656 229032 214708 229084
rect 223488 229032 223540 229084
rect 289912 229032 289964 229084
rect 238024 228352 238076 228404
rect 263784 228352 263836 228404
rect 49516 227740 49568 227792
rect 55128 227740 55180 227792
rect 169944 227740 169996 227792
rect 170496 227740 170548 227792
rect 178868 227740 178920 227792
rect 179328 227740 179380 227792
rect 222936 227740 222988 227792
rect 223488 227740 223540 227792
rect 189724 227060 189776 227112
rect 209044 227060 209096 227112
rect 108488 226992 108540 227044
rect 229100 226992 229152 227044
rect 229928 226992 229980 227044
rect 256056 226788 256108 226840
rect 259644 226788 259696 226840
rect 229928 226312 229980 226364
rect 256056 226312 256108 226364
rect 137560 226244 137612 226296
rect 280436 226244 280488 226296
rect 210516 226176 210568 226228
rect 262496 226176 262548 226228
rect 280160 225020 280212 225072
rect 280436 225020 280488 225072
rect 67364 224952 67416 225004
rect 204168 224952 204220 225004
rect 210516 224952 210568 225004
rect 210976 224952 211028 225004
rect 166356 224884 166408 224936
rect 166908 224884 166960 224936
rect 204352 224884 204404 224936
rect 50804 224204 50856 224256
rect 160744 224204 160796 224256
rect 191288 224204 191340 224256
rect 194600 224204 194652 224256
rect 206284 224204 206336 224256
rect 252560 224204 252612 224256
rect 253204 224204 253256 224256
rect 270592 224204 270644 224256
rect 165528 223524 165580 223576
rect 274916 223524 274968 223576
rect 56508 222844 56560 222896
rect 163688 222844 163740 222896
rect 164148 222844 164200 222896
rect 220084 222844 220136 222896
rect 252744 222844 252796 222896
rect 64604 222096 64656 222148
rect 153108 222096 153160 222148
rect 204168 222096 204220 222148
rect 265164 222096 265216 222148
rect 153108 221416 153160 221468
rect 187608 221416 187660 221468
rect 195980 221416 196032 221468
rect 252560 221416 252612 221468
rect 274824 221416 274876 221468
rect 102784 220736 102836 220788
rect 263692 220736 263744 220788
rect 53656 220056 53708 220108
rect 171876 220056 171928 220108
rect 222844 220056 222896 220108
rect 252652 220056 252704 220108
rect 256056 220056 256108 220108
rect 580356 220056 580408 220108
rect 160744 219376 160796 219428
rect 161388 219376 161440 219428
rect 278044 219376 278096 219428
rect 47584 218764 47636 218816
rect 106924 218764 106976 218816
rect 92572 218696 92624 218748
rect 153844 218696 153896 218748
rect 154028 218696 154080 218748
rect 256608 218696 256660 218748
rect 258540 218696 258592 218748
rect 71780 217948 71832 218000
rect 73068 217948 73120 218000
rect 167000 217948 167052 218000
rect 271880 217948 271932 218000
rect 172060 217880 172112 217932
rect 224224 217880 224276 217932
rect 106096 217268 106148 217320
rect 120172 217268 120224 217320
rect 239404 217268 239456 217320
rect 249156 217268 249208 217320
rect 171876 216656 171928 216708
rect 172060 216656 172112 216708
rect 98736 216588 98788 216640
rect 103612 216588 103664 216640
rect 264980 216588 265032 216640
rect 184296 216520 184348 216572
rect 247776 216520 247828 216572
rect 119344 215908 119396 215960
rect 159548 215908 159600 215960
rect 258724 215908 258776 215960
rect 273260 215908 273312 215960
rect 184296 215636 184348 215688
rect 184848 215636 184900 215688
rect 3976 214888 4028 214940
rect 7564 214888 7616 214940
rect 105636 214548 105688 214600
rect 244924 214548 244976 214600
rect 95240 213188 95292 213240
rect 117412 213188 117464 213240
rect 117412 212508 117464 212560
rect 258080 212508 258132 212560
rect 258632 212508 258684 212560
rect 50988 212440 51040 212492
rect 269396 212440 269448 212492
rect 149796 212372 149848 212424
rect 222384 212372 222436 212424
rect 222936 212372 222988 212424
rect 142988 210468 143040 210520
rect 236000 210468 236052 210520
rect 78588 210400 78640 210452
rect 106924 210400 106976 210452
rect 257344 210400 257396 210452
rect 173808 209720 173860 209772
rect 278964 209720 279016 209772
rect 97356 209108 97408 209160
rect 108120 209108 108172 209160
rect 57704 209040 57756 209092
rect 173808 209040 173860 209092
rect 107752 208360 107804 208412
rect 108120 208360 108172 208412
rect 263600 208360 263652 208412
rect 263968 208360 264020 208412
rect 86960 207680 87012 207732
rect 103612 207680 103664 207732
rect 104808 207680 104860 207732
rect 13820 207612 13872 207664
rect 189080 207612 189132 207664
rect 104808 207000 104860 207052
rect 269304 207000 269356 207052
rect 96620 206320 96672 206372
rect 109224 206320 109276 206372
rect 84108 206252 84160 206304
rect 113272 206252 113324 206304
rect 113916 206252 113968 206304
rect 227720 206252 227772 206304
rect 270684 206252 270736 206304
rect 109224 205708 109276 205760
rect 227720 205708 227772 205760
rect 113916 205640 113968 205692
rect 260932 205640 260984 205692
rect 77300 204892 77352 204944
rect 109132 204892 109184 204944
rect 255964 204892 256016 204944
rect 265072 204892 265124 204944
rect 159548 204212 159600 204264
rect 292672 204212 292724 204264
rect 203524 203532 203576 203584
rect 281816 203532 281868 203584
rect 98092 202784 98144 202836
rect 98828 202784 98880 202836
rect 3332 202172 3384 202224
rect 98092 202172 98144 202224
rect 175096 202172 175148 202224
rect 209136 202172 209188 202224
rect 38660 202104 38712 202156
rect 182824 202104 182876 202156
rect 192576 202104 192628 202156
rect 228364 202104 228416 202156
rect 54944 201424 54996 201476
rect 291292 201424 291344 201476
rect 243544 200744 243596 200796
rect 268384 200744 268436 200796
rect 249708 199384 249760 199436
rect 293960 199384 294012 199436
rect 129096 198636 129148 198688
rect 256700 198636 256752 198688
rect 195244 197956 195296 198008
rect 280344 197956 280396 198008
rect 23480 196596 23532 196648
rect 187056 196596 187108 196648
rect 200028 196596 200080 196648
rect 582472 196596 582524 196648
rect 244924 195916 244976 195968
rect 272524 195916 272576 195968
rect 90364 195236 90416 195288
rect 129096 195236 129148 195288
rect 137376 195236 137428 195288
rect 150440 195236 150492 195288
rect 164976 195236 165028 195288
rect 196624 195236 196676 195288
rect 272524 195236 272576 195288
rect 579988 195236 580040 195288
rect 162676 194488 162728 194540
rect 170404 194488 170456 194540
rect 131764 193876 131816 193928
rect 145564 193876 145616 193928
rect 61844 193808 61896 193860
rect 69020 193808 69072 193860
rect 123484 193808 123536 193860
rect 137468 193808 137520 193860
rect 138664 193808 138716 193860
rect 148508 193808 148560 193860
rect 170496 193808 170548 193860
rect 189724 193808 189776 193860
rect 49700 189728 49752 189780
rect 193312 189728 193364 189780
rect 213184 189728 213236 189780
rect 295432 189728 295484 189780
rect 3424 188980 3476 189032
rect 43444 188980 43496 189032
rect 232504 188300 232556 188352
rect 276296 188300 276348 188352
rect 48320 186940 48372 186992
rect 120816 186940 120868 186992
rect 195336 186940 195388 186992
rect 226340 186940 226392 186992
rect 133144 185648 133196 185700
rect 147128 185648 147180 185700
rect 45468 185580 45520 185632
rect 73436 185580 73488 185632
rect 118792 185580 118844 185632
rect 138756 185580 138808 185632
rect 145564 184968 145616 185020
rect 153936 184968 153988 185020
rect 195336 184152 195388 184204
rect 249064 184152 249116 184204
rect 122104 182860 122156 182912
rect 134708 182860 134760 182912
rect 89536 182792 89588 182844
rect 124312 182792 124364 182844
rect 69664 180820 69716 180872
rect 175924 180820 175976 180872
rect 214564 180140 214616 180192
rect 224960 180140 225012 180192
rect 91008 180072 91060 180124
rect 107660 180072 107712 180124
rect 122840 180072 122892 180124
rect 140136 180072 140188 180124
rect 207756 180072 207808 180124
rect 287244 180072 287296 180124
rect 191104 179732 191156 179784
rect 198924 179732 198976 179784
rect 1400 178644 1452 178696
rect 145656 178644 145708 178696
rect 198004 178644 198056 178696
rect 234620 178644 234672 178696
rect 241428 178644 241480 178696
rect 580172 178644 580224 178696
rect 240784 178032 240836 178084
rect 241428 178032 241480 178084
rect 85488 177284 85540 177336
rect 213184 177284 213236 177336
rect 228364 177284 228416 177336
rect 251824 177284 251876 177336
rect 84200 176672 84252 176724
rect 85488 176672 85540 176724
rect 93124 176672 93176 176724
rect 93676 176672 93728 176724
rect 220084 176672 220136 176724
rect 88984 175924 89036 175976
rect 121552 175924 121604 175976
rect 214012 175924 214064 175976
rect 214012 175244 214064 175296
rect 247684 175244 247736 175296
rect 255320 175244 255372 175296
rect 256608 175244 256660 175296
rect 583024 175244 583076 175296
rect 196072 175176 196124 175228
rect 196808 175176 196860 175228
rect 205732 174700 205784 174752
rect 206284 174700 206336 174752
rect 82084 174496 82136 174548
rect 82728 174496 82780 174548
rect 205732 174496 205784 174548
rect 88340 173884 88392 173936
rect 196808 173884 196860 173936
rect 137468 172592 137520 172644
rect 228364 172592 228416 172644
rect 205732 172524 205784 172576
rect 320180 172524 320232 172576
rect 85580 171844 85632 171896
rect 106280 171844 106332 171896
rect 91008 171776 91060 171828
rect 180156 171776 180208 171828
rect 221464 171776 221516 171828
rect 237380 171776 237432 171828
rect 256700 171776 256752 171828
rect 112444 171096 112496 171148
rect 230572 171096 230624 171148
rect 194876 170620 194928 170672
rect 195336 170620 195388 170672
rect 56324 170348 56376 170400
rect 194876 170348 194928 170400
rect 196716 170348 196768 170400
rect 205640 170348 205692 170400
rect 215392 170348 215444 170400
rect 259460 170348 259512 170400
rect 115296 169736 115348 169788
rect 204720 169736 204772 169788
rect 262680 168988 262732 169040
rect 276204 168988 276256 169040
rect 87696 168444 87748 168496
rect 200672 168444 200724 168496
rect 204260 168444 204312 168496
rect 204720 168444 204772 168496
rect 262312 168444 262364 168496
rect 262680 168444 262732 168496
rect 92664 168376 92716 168428
rect 222200 168376 222252 168428
rect 222844 168376 222896 168428
rect 76748 167628 76800 167680
rect 202880 167628 202932 167680
rect 203524 167628 203576 167680
rect 222292 167628 222344 167680
rect 238024 167628 238076 167680
rect 75920 167016 75972 167068
rect 76748 167016 76800 167068
rect 195980 167016 196032 167068
rect 196624 167016 196676 167068
rect 303620 167016 303672 167068
rect 169116 165656 169168 165708
rect 224224 165656 224276 165708
rect 82912 165588 82964 165640
rect 204996 165588 205048 165640
rect 199384 164840 199436 164892
rect 260840 164840 260892 164892
rect 65892 164296 65944 164348
rect 154028 164296 154080 164348
rect 82176 164228 82228 164280
rect 208400 164228 208452 164280
rect 224776 163480 224828 163532
rect 283104 163480 283156 163532
rect 60556 162936 60608 162988
rect 152648 162936 152700 162988
rect 2872 162868 2924 162920
rect 4804 162868 4856 162920
rect 92480 162868 92532 162920
rect 222292 162868 222344 162920
rect 133236 161984 133288 162036
rect 133696 161984 133748 162036
rect 133236 161508 133288 161560
rect 226524 161508 226576 161560
rect 87144 161440 87196 161492
rect 215392 161440 215444 161492
rect 231124 160760 231176 160812
rect 274732 160760 274784 160812
rect 97908 160692 97960 160744
rect 249800 160692 249852 160744
rect 97356 160148 97408 160200
rect 97908 160148 97960 160200
rect 91744 160080 91796 160132
rect 92296 160080 92348 160132
rect 218796 160080 218848 160132
rect 249616 159400 249668 159452
rect 202788 159332 202840 159384
rect 269212 159332 269264 159384
rect 278872 159332 278924 159384
rect 338764 159332 338816 159384
rect 198740 159196 198792 159248
rect 199384 159196 199436 159248
rect 72976 158788 73028 158840
rect 198740 158788 198792 158840
rect 91836 158720 91888 158772
rect 92388 158720 92440 158772
rect 221004 158720 221056 158772
rect 192484 158652 192536 158704
rect 249616 158652 249668 158704
rect 56416 157972 56468 158024
rect 74632 157972 74684 158024
rect 76564 157972 76616 158024
rect 107016 157972 107068 158024
rect 154028 157972 154080 158024
rect 187700 157972 187752 158024
rect 98000 157360 98052 157412
rect 98828 157360 98880 157412
rect 227720 157360 227772 157412
rect 187700 157292 187752 157344
rect 188896 157292 188948 157344
rect 214656 157292 214708 157344
rect 35808 156612 35860 156664
rect 67732 156612 67784 156664
rect 68928 156612 68980 156664
rect 68928 156000 68980 156052
rect 188436 156000 188488 156052
rect 210516 156000 210568 156052
rect 210976 156000 211028 156052
rect 229100 156000 229152 156052
rect 75184 155932 75236 155984
rect 201684 155932 201736 155984
rect 202788 155932 202840 155984
rect 218060 155932 218112 155984
rect 218888 155932 218940 155984
rect 246396 155932 246448 155984
rect 60464 155864 60516 155916
rect 60648 155864 60700 155916
rect 294696 155184 294748 155236
rect 583116 155184 583168 155236
rect 60464 154640 60516 154692
rect 154028 154640 154080 154692
rect 158720 154640 158772 154692
rect 160008 154640 160060 154692
rect 186964 154640 187016 154692
rect 187700 154640 187752 154692
rect 224960 154640 225012 154692
rect 88616 154572 88668 154624
rect 218704 154572 218756 154624
rect 93860 153892 93912 153944
rect 131120 153892 131172 153944
rect 223672 153892 223724 153944
rect 65984 153824 66036 153876
rect 158720 153824 158772 153876
rect 192484 153824 192536 153876
rect 218060 153824 218112 153876
rect 187516 153212 187568 153264
rect 191840 153212 191892 153264
rect 222384 152464 222436 152516
rect 222844 152464 222896 152516
rect 182916 151920 182968 151972
rect 222844 151920 222896 151972
rect 62028 151852 62080 151904
rect 131856 151852 131908 151904
rect 151268 151852 151320 151904
rect 208492 151852 208544 151904
rect 69756 151784 69808 151836
rect 160192 151784 160244 151836
rect 160744 151784 160796 151836
rect 220820 151784 220872 151836
rect 222108 151784 222160 151836
rect 302240 151784 302292 151836
rect 74816 151104 74868 151156
rect 177948 151104 178000 151156
rect 63408 151036 63460 151088
rect 167644 151036 167696 151088
rect 189632 151104 189684 151156
rect 201500 151104 201552 151156
rect 201592 151036 201644 151088
rect 207848 151036 207900 151088
rect 220820 151036 220872 151088
rect 204168 150424 204220 150476
rect 230664 150424 230716 150476
rect 148600 149744 148652 149796
rect 204168 149744 204220 149796
rect 206376 149744 206428 149796
rect 252468 149744 252520 149796
rect 86868 149676 86920 149728
rect 124864 149676 124916 149728
rect 216772 149676 216824 149728
rect 252468 149132 252520 149184
rect 256056 149132 256108 149184
rect 67548 149064 67600 149116
rect 111156 149064 111208 149116
rect 216864 149064 216916 149116
rect 217324 149064 217376 149116
rect 582748 149064 582800 149116
rect 193036 148996 193088 149048
rect 211068 148996 211120 149048
rect 218520 148996 218572 149048
rect 218704 148996 218756 149048
rect 267832 148996 267884 149048
rect 190368 148384 190420 148436
rect 193220 148384 193272 148436
rect 64696 148316 64748 148368
rect 192484 148316 192536 148368
rect 48228 147636 48280 147688
rect 104164 147636 104216 147688
rect 213000 147636 213052 147688
rect 233884 147636 233936 147688
rect 214012 147568 214064 147620
rect 216864 147568 216916 147620
rect 208400 146956 208452 147008
rect 209136 146956 209188 147008
rect 3148 146888 3200 146940
rect 95424 146888 95476 146940
rect 153936 146888 153988 146940
rect 154028 146888 154080 146940
rect 187700 146888 187752 146940
rect 252192 146888 252244 146940
rect 288716 146888 288768 146940
rect 327080 146888 327132 146940
rect 221464 146344 221516 146396
rect 256148 146344 256200 146396
rect 67272 146276 67324 146328
rect 97448 146276 97500 146328
rect 100024 146276 100076 146328
rect 100576 146276 100628 146328
rect 224960 146276 225012 146328
rect 4804 146208 4856 146260
rect 86868 146208 86920 146260
rect 87604 146208 87656 146260
rect 89628 146208 89680 146260
rect 95240 146208 95292 146260
rect 218796 146208 218848 146260
rect 221096 146208 221148 146260
rect 204904 145528 204956 145580
rect 234712 145528 234764 145580
rect 259368 145528 259420 145580
rect 277584 145528 277636 145580
rect 177856 144984 177908 145036
rect 209872 144984 209924 145036
rect 71780 144916 71832 144968
rect 72884 144916 72936 144968
rect 198372 144916 198424 144968
rect 228364 144916 228416 144968
rect 349804 144916 349856 144968
rect 85580 144712 85632 144764
rect 88984 144712 89036 144764
rect 90088 144712 90140 144764
rect 93124 144712 93176 144764
rect 186964 144372 187016 144424
rect 193588 144372 193640 144424
rect 175924 144236 175976 144288
rect 194140 144236 194192 144288
rect 102140 144168 102192 144220
rect 178776 144168 178828 144220
rect 224500 144168 224552 144220
rect 224868 144168 224920 144220
rect 238116 144168 238168 144220
rect 249064 144168 249116 144220
rect 262220 144168 262272 144220
rect 223672 144032 223724 144084
rect 224500 144032 224552 144084
rect 200120 143964 200172 144016
rect 200396 143964 200448 144016
rect 204260 143964 204312 144016
rect 204628 143964 204680 144016
rect 59268 143556 59320 143608
rect 167736 143556 167788 143608
rect 195428 143488 195480 143540
rect 197912 143488 197964 143540
rect 245016 143556 245068 143608
rect 219532 143488 219584 143540
rect 220176 143488 220228 143540
rect 259368 143488 259420 143540
rect 260104 143488 260156 143540
rect 60648 142808 60700 142860
rect 77944 142808 77996 142860
rect 120724 142808 120776 142860
rect 199016 142876 199068 142928
rect 218244 142876 218296 142928
rect 212908 142808 212960 142860
rect 259368 142808 259420 142860
rect 63132 142128 63184 142180
rect 88524 142128 88576 142180
rect 220084 142128 220136 142180
rect 225696 142128 225748 142180
rect 69848 142060 69900 142112
rect 76012 142060 76064 142112
rect 76012 141380 76064 141432
rect 159456 141380 159508 141432
rect 203156 141380 203208 141432
rect 69112 140836 69164 140888
rect 69848 140836 69900 140888
rect 205640 140836 205692 140888
rect 266360 140836 266412 140888
rect 267004 140836 267056 140888
rect 57796 140768 57848 140820
rect 91100 140768 91152 140820
rect 203432 140768 203484 140820
rect 289084 140768 289136 140820
rect 193036 140496 193088 140548
rect 194876 140496 194928 140548
rect 89076 140088 89128 140140
rect 120724 140088 120776 140140
rect 193404 140088 193456 140140
rect 210148 140564 210200 140616
rect 68652 140020 68704 140072
rect 80704 140020 80756 140072
rect 84476 140020 84528 140072
rect 118884 140020 118936 140072
rect 173256 140020 173308 140072
rect 184480 140020 184532 140072
rect 71320 139408 71372 139460
rect 73804 139408 73856 139460
rect 118884 139408 118936 139460
rect 205180 140428 205232 140480
rect 210056 140496 210108 140548
rect 212540 140428 212592 140480
rect 79416 139340 79468 139392
rect 215392 140428 215444 140480
rect 225144 140428 225196 140480
rect 287704 140020 287756 140072
rect 225144 139408 225196 139460
rect 249708 139408 249760 139460
rect 251180 139408 251232 139460
rect 226708 139204 226760 139256
rect 229192 139204 229244 139256
rect 66168 138660 66220 138712
rect 178684 138660 178736 138712
rect 236000 138660 236052 138712
rect 582656 138660 582708 138712
rect 93860 138048 93912 138100
rect 94320 138048 94372 138100
rect 65892 137980 65944 138032
rect 66168 137980 66220 138032
rect 2872 137912 2924 137964
rect 72976 137912 73028 137964
rect 73160 137912 73212 137964
rect 78496 137912 78548 137964
rect 79416 137912 79468 137964
rect 87052 137912 87104 137964
rect 193220 137912 193272 137964
rect 226708 137912 226760 137964
rect 234620 137912 234672 137964
rect 240876 137912 240928 137964
rect 58900 137232 58952 137284
rect 69204 137232 69256 137284
rect 91100 137232 91152 137284
rect 151360 137232 151412 137284
rect 247684 137232 247736 137284
rect 255320 137232 255372 137284
rect 256148 137232 256200 137284
rect 276020 137232 276072 137284
rect 91008 136824 91060 136876
rect 91836 136824 91888 136876
rect 79600 136620 79652 136672
rect 87052 136688 87104 136740
rect 81348 136620 81400 136672
rect 82176 136620 82228 136672
rect 85488 136620 85540 136672
rect 86224 136620 86276 136672
rect 91192 136552 91244 136604
rect 91744 136552 91796 136604
rect 170404 136552 170456 136604
rect 191564 136552 191616 136604
rect 159456 135940 159508 135992
rect 169024 135940 169076 135992
rect 160192 135872 160244 135924
rect 161388 135872 161440 135924
rect 175924 135872 175976 135924
rect 256056 135872 256108 135924
rect 298744 135872 298796 135924
rect 53104 135328 53156 135380
rect 91284 135328 91336 135380
rect 4804 135260 4856 135312
rect 91192 135260 91244 135312
rect 187700 135260 187752 135312
rect 191564 135260 191616 135312
rect 97908 135192 97960 135244
rect 137468 135192 137520 135244
rect 226708 135192 226760 135244
rect 231952 135192 232004 135244
rect 188436 134852 188488 134904
rect 191196 134852 191248 134904
rect 70308 134784 70360 134836
rect 75368 134784 75420 134836
rect 68560 134580 68612 134632
rect 69756 134580 69808 134632
rect 93768 134580 93820 134632
rect 189172 134512 189224 134564
rect 226616 134512 226668 134564
rect 309784 134512 309836 134564
rect 95148 133832 95200 133884
rect 177580 133832 177632 133884
rect 226616 133832 226668 133884
rect 237380 133832 237432 133884
rect 226708 133628 226760 133680
rect 231124 133628 231176 133680
rect 148508 133220 148560 133272
rect 187700 133220 187752 133272
rect 103704 133152 103756 133204
rect 148600 133152 148652 133204
rect 52184 132404 52236 132456
rect 66904 132404 66956 132456
rect 97908 132404 97960 132456
rect 142988 132404 143040 132456
rect 226708 132404 226760 132456
rect 249892 132404 249944 132456
rect 56324 132336 56376 132388
rect 66812 132336 66864 132388
rect 180156 131792 180208 131844
rect 190460 131792 190512 131844
rect 150440 131724 150492 131776
rect 182916 131724 182968 131776
rect 240784 131724 240836 131776
rect 335452 131724 335504 131776
rect 104900 131112 104952 131164
rect 111064 131112 111116 131164
rect 63132 131044 63184 131096
rect 66812 131044 66864 131096
rect 169208 131044 169260 131096
rect 189816 131044 189868 131096
rect 226708 131044 226760 131096
rect 230664 131044 230716 131096
rect 276112 131044 276164 131096
rect 226800 130976 226852 131028
rect 233240 130976 233292 131028
rect 267740 130976 267792 131028
rect 97540 130568 97592 130620
rect 102876 130568 102928 130620
rect 97724 130364 97776 130416
rect 181536 130364 181588 130416
rect 97908 129684 97960 129736
rect 106372 129684 106424 129736
rect 151360 129684 151412 129736
rect 191748 129684 191800 129736
rect 114560 129072 114612 129124
rect 148416 129072 148468 129124
rect 97448 129004 97500 129056
rect 160836 129004 160888 129056
rect 61752 128324 61804 128376
rect 66812 128324 66864 128376
rect 226432 128324 226484 128376
rect 299480 128324 299532 128376
rect 97632 128256 97684 128308
rect 140136 128256 140188 128308
rect 227904 127644 227956 127696
rect 267832 127644 267884 127696
rect 109132 127576 109184 127628
rect 133236 127576 133288 127628
rect 158076 127576 158128 127628
rect 183468 127576 183520 127628
rect 226708 127576 226760 127628
rect 340880 127576 340932 127628
rect 183468 126964 183520 127016
rect 191748 126964 191800 127016
rect 64512 126896 64564 126948
rect 66812 126896 66864 126948
rect 226708 126896 226760 126948
rect 249800 126896 249852 126948
rect 251088 126896 251140 126948
rect 97908 126828 97960 126880
rect 103704 126828 103756 126880
rect 97172 126216 97224 126268
rect 109132 126216 109184 126268
rect 179236 126216 179288 126268
rect 187516 126216 187568 126268
rect 191564 126216 191616 126268
rect 251088 126216 251140 126268
rect 351920 126216 351972 126268
rect 97908 125536 97960 125588
rect 155408 125536 155460 125588
rect 155868 125536 155920 125588
rect 156696 125536 156748 125588
rect 167736 125536 167788 125588
rect 190368 125536 190420 125588
rect 59268 124924 59320 124976
rect 66812 124924 66864 124976
rect 57796 124856 57848 124908
rect 66996 124856 67048 124908
rect 238116 124856 238168 124908
rect 305644 124856 305696 124908
rect 97816 124788 97868 124840
rect 100760 124788 100812 124840
rect 101588 124176 101640 124228
rect 155868 124176 155920 124228
rect 60464 124108 60516 124160
rect 66904 124108 66956 124160
rect 97908 124108 97960 124160
rect 150440 124108 150492 124160
rect 160744 124108 160796 124160
rect 180156 124108 180208 124160
rect 226708 124108 226760 124160
rect 230572 124108 230624 124160
rect 279424 124108 279476 124160
rect 582840 124108 582892 124160
rect 175924 124040 175976 124092
rect 191748 124040 191800 124092
rect 235264 123428 235316 123480
rect 243544 123428 243596 123480
rect 63316 122748 63368 122800
rect 66352 122748 66404 122800
rect 97908 122748 97960 122800
rect 153936 122748 153988 122800
rect 226524 122748 226576 122800
rect 240232 122748 240284 122800
rect 250536 122068 250588 122120
rect 285680 122068 285732 122120
rect 189080 121592 189132 121644
rect 191748 121592 191800 121644
rect 53748 121388 53800 121440
rect 66904 121388 66956 121440
rect 131856 121388 131908 121440
rect 188988 121388 189040 121440
rect 191012 121388 191064 121440
rect 226708 121388 226760 121440
rect 234712 121388 234764 121440
rect 61936 121320 61988 121372
rect 66812 121320 66864 121372
rect 97080 121320 97132 121372
rect 145656 121320 145708 121372
rect 159548 121320 159600 121372
rect 191196 121320 191248 121372
rect 240784 120776 240836 120828
rect 252560 120776 252612 120828
rect 232504 120708 232556 120760
rect 313280 120708 313332 120760
rect 96068 120300 96120 120352
rect 98828 120300 98880 120352
rect 64696 120028 64748 120080
rect 66812 120028 66864 120080
rect 97908 120028 97960 120080
rect 112444 120028 112496 120080
rect 184296 120028 184348 120080
rect 191748 120028 191800 120080
rect 59084 119960 59136 120012
rect 66904 119960 66956 120012
rect 104164 119348 104216 119400
rect 187700 119348 187752 119400
rect 284300 119348 284352 119400
rect 289820 119348 289872 119400
rect 52276 118600 52328 118652
rect 66628 118600 66680 118652
rect 97908 118600 97960 118652
rect 134708 118600 134760 118652
rect 186136 118600 186188 118652
rect 188988 118600 189040 118652
rect 167644 117920 167696 117972
rect 191748 117920 191800 117972
rect 226524 117376 226576 117428
rect 231124 117376 231176 117428
rect 99472 117308 99524 117360
rect 100668 117308 100720 117360
rect 160744 117308 160796 117360
rect 226616 117308 226668 117360
rect 244280 117308 244332 117360
rect 62028 117240 62080 117292
rect 66628 117240 66680 117292
rect 97356 117240 97408 117292
rect 178868 117240 178920 117292
rect 97908 117172 97960 117224
rect 177488 117172 177540 117224
rect 230388 116628 230440 116680
rect 262404 116628 262456 116680
rect 245016 116560 245068 116612
rect 285680 116560 285732 116612
rect 188436 116084 188488 116136
rect 191564 116084 191616 116136
rect 226708 115948 226760 116000
rect 229192 115948 229244 116000
rect 230388 115948 230440 116000
rect 50896 115880 50948 115932
rect 66812 115880 66864 115932
rect 97816 115880 97868 115932
rect 99472 115880 99524 115932
rect 226156 115880 226208 115932
rect 280160 115880 280212 115932
rect 186228 115608 186280 115660
rect 191748 115608 191800 115660
rect 63408 115540 63460 115592
rect 66904 115540 66956 115592
rect 97908 114520 97960 114572
rect 188344 114520 188396 114572
rect 60556 114452 60608 114504
rect 66812 114452 66864 114504
rect 187700 114452 187752 114504
rect 191748 114452 191800 114504
rect 226432 113840 226484 113892
rect 250536 113840 250588 113892
rect 7564 113772 7616 113824
rect 63408 113772 63460 113824
rect 66904 113772 66956 113824
rect 110512 113772 110564 113824
rect 134616 113772 134668 113824
rect 246396 113772 246448 113824
rect 270500 113772 270552 113824
rect 97540 113160 97592 113212
rect 169024 113160 169076 113212
rect 55128 113092 55180 113144
rect 66812 113092 66864 113144
rect 169668 112412 169720 112464
rect 191748 112412 191800 112464
rect 225696 112412 225748 112464
rect 252560 112412 252612 112464
rect 269120 112412 269172 112464
rect 96712 111868 96764 111920
rect 98644 111868 98696 111920
rect 102048 111868 102100 111920
rect 166264 111868 166316 111920
rect 169116 111868 169168 111920
rect 169668 111868 169720 111920
rect 97908 111800 97960 111852
rect 189724 111800 189776 111852
rect 226340 111800 226392 111852
rect 231952 111800 232004 111852
rect 295340 111800 295392 111852
rect 43996 111732 44048 111784
rect 66812 111732 66864 111784
rect 185584 111732 185636 111784
rect 191748 111732 191800 111784
rect 226708 111528 226760 111580
rect 230480 111528 230532 111580
rect 96804 111120 96856 111172
rect 100024 111120 100076 111172
rect 39948 111052 40000 111104
rect 59268 111052 59320 111104
rect 66904 111052 66956 111104
rect 100116 111052 100168 111104
rect 188436 111052 188488 111104
rect 226340 111052 226392 111104
rect 295340 111052 295392 111104
rect 324320 111052 324372 111104
rect 295432 110984 295484 111036
rect 2872 110780 2924 110832
rect 4804 110780 4856 110832
rect 190368 110440 190420 110492
rect 191840 110440 191892 110492
rect 295432 110440 295484 110492
rect 295984 110440 296036 110492
rect 97816 110372 97868 110424
rect 102048 110372 102100 110424
rect 111156 110372 111208 110424
rect 190644 110372 190696 110424
rect 231124 110372 231176 110424
rect 299664 110372 299716 110424
rect 307024 110372 307076 110424
rect 97908 110304 97960 110356
rect 173256 110304 173308 110356
rect 48228 109012 48280 109064
rect 53840 109012 53892 109064
rect 66904 109012 66956 109064
rect 54944 108944 54996 108996
rect 66812 108944 66864 108996
rect 165528 108944 165580 108996
rect 189080 108944 189132 108996
rect 187608 108876 187660 108928
rect 191748 108876 191800 108928
rect 226524 108876 226576 108928
rect 229100 108876 229152 108928
rect 98828 108332 98880 108384
rect 113272 108332 113324 108384
rect 97908 108264 97960 108316
rect 109040 108264 109092 108316
rect 109684 108264 109736 108316
rect 112444 108264 112496 108316
rect 165528 108264 165580 108316
rect 226984 108264 227036 108316
rect 263692 108264 263744 108316
rect 64604 107584 64656 107636
rect 66628 107584 66680 107636
rect 97908 107584 97960 107636
rect 177396 107584 177448 107636
rect 182824 107584 182876 107636
rect 190828 107584 190880 107636
rect 226708 107584 226760 107636
rect 285772 107584 285824 107636
rect 286232 107584 286284 107636
rect 286232 106904 286284 106956
rect 342904 106904 342956 106956
rect 97908 106496 97960 106548
rect 101680 106496 101732 106548
rect 7564 106292 7616 106344
rect 66812 106292 66864 106344
rect 160836 106224 160888 106276
rect 191196 106224 191248 106276
rect 46848 105544 46900 105596
rect 66168 105544 66220 105596
rect 66628 105544 66680 105596
rect 106188 105544 106240 105596
rect 120172 105544 120224 105596
rect 177396 105544 177448 105596
rect 178684 105544 178736 105596
rect 187608 105544 187660 105596
rect 191748 105544 191800 105596
rect 226340 105544 226392 105596
rect 240784 105544 240836 105596
rect 245016 105544 245068 105596
rect 273260 105544 273312 105596
rect 226708 105000 226760 105052
rect 230572 105000 230624 105052
rect 56508 104796 56560 104848
rect 66812 104796 66864 104848
rect 101312 104796 101364 104848
rect 101496 104796 101548 104848
rect 270408 104796 270460 104848
rect 274640 104796 274692 104848
rect 97908 104184 97960 104236
rect 106188 104184 106240 104236
rect 225696 104116 225748 104168
rect 255964 104116 256016 104168
rect 97908 103436 97960 103488
rect 101312 103436 101364 103488
rect 185584 103504 185636 103556
rect 226708 103504 226760 103556
rect 229100 103504 229152 103556
rect 270408 103504 270460 103556
rect 55036 103368 55088 103420
rect 66444 103368 66496 103420
rect 97908 103028 97960 103080
rect 99380 103028 99432 103080
rect 99380 102756 99432 102808
rect 182824 102756 182876 102808
rect 226708 102756 226760 102808
rect 230480 102756 230532 102808
rect 282920 102756 282972 102808
rect 321652 102756 321704 102808
rect 188528 102144 188580 102196
rect 191012 102144 191064 102196
rect 226708 102144 226760 102196
rect 237380 102144 237432 102196
rect 97908 102076 97960 102128
rect 129188 102076 129240 102128
rect 226340 102076 226392 102128
rect 266452 102076 266504 102128
rect 166908 101464 166960 101516
rect 180800 101464 180852 101516
rect 181904 101464 181956 101516
rect 55128 101396 55180 101448
rect 59176 101396 59228 101448
rect 66720 101396 66772 101448
rect 104164 101396 104216 101448
rect 117412 101396 117464 101448
rect 129188 101396 129240 101448
rect 153936 101396 153988 101448
rect 155868 101396 155920 101448
rect 186964 101396 187016 101448
rect 226708 101396 226760 101448
rect 277400 101396 277452 101448
rect 64696 100716 64748 100768
rect 66812 100716 66864 100768
rect 120724 100716 120776 100768
rect 163504 100716 163556 100768
rect 164148 100716 164200 100768
rect 181904 100716 181956 100768
rect 191748 100716 191800 100768
rect 97908 99968 97960 100020
rect 101404 99968 101456 100020
rect 185676 99968 185728 100020
rect 64788 99628 64840 99680
rect 66812 99628 66864 99680
rect 97540 99356 97592 99408
rect 129648 99356 129700 99408
rect 226340 99356 226392 99408
rect 327724 99356 327776 99408
rect 53656 99288 53708 99340
rect 66812 99288 66864 99340
rect 271880 99288 271932 99340
rect 580172 99288 580224 99340
rect 246488 98744 246540 98796
rect 269304 98744 269356 98796
rect 262864 98676 262916 98728
rect 271880 98676 271932 98728
rect 97540 98608 97592 98660
rect 107752 98608 107804 98660
rect 226616 98608 226668 98660
rect 237288 98608 237340 98660
rect 247684 98608 247736 98660
rect 184296 98064 184348 98116
rect 191748 98064 191800 98116
rect 97908 97996 97960 98048
rect 188804 97996 188856 98048
rect 180248 97928 180300 97980
rect 191656 97928 191708 97980
rect 101404 97248 101456 97300
rect 169116 97248 169168 97300
rect 227168 97248 227220 97300
rect 263600 97248 263652 97300
rect 96712 96976 96764 97028
rect 98736 96976 98788 97028
rect 3056 96636 3108 96688
rect 65524 96636 65576 96688
rect 99012 96636 99064 96688
rect 114652 96636 114704 96688
rect 115848 96636 115900 96688
rect 226708 96568 226760 96620
rect 264980 96568 265032 96620
rect 115848 95888 115900 95940
rect 191932 95888 191984 95940
rect 227996 95888 228048 95940
rect 244924 95888 244976 95940
rect 97908 95208 97960 95260
rect 177488 95208 177540 95260
rect 57704 95140 57756 95192
rect 66812 95140 66864 95192
rect 95976 94528 96028 94580
rect 110604 94528 110656 94580
rect 94872 94460 94924 94512
rect 124312 94460 124364 94512
rect 191840 94460 191892 94512
rect 158628 93848 158680 93900
rect 192024 93848 192076 93900
rect 57888 93780 57940 93832
rect 67180 93780 67232 93832
rect 67456 93780 67508 93832
rect 67732 93780 67784 93832
rect 97908 93780 97960 93832
rect 109224 93780 109276 93832
rect 224040 93372 224092 93424
rect 225144 93372 225196 93424
rect 222108 93304 222160 93356
rect 225696 93304 225748 93356
rect 247684 93100 247736 93152
rect 331220 93100 331272 93152
rect 88662 92692 88714 92744
rect 90134 92624 90186 92676
rect 91008 92624 91060 92676
rect 94872 92624 94924 92676
rect 93814 92556 93866 92608
rect 94504 92556 94556 92608
rect 95884 92556 95936 92608
rect 94688 92488 94740 92540
rect 104164 92488 104216 92540
rect 191932 92488 191984 92540
rect 207388 92488 207440 92540
rect 212908 92488 212960 92540
rect 242256 92488 242308 92540
rect 67364 92420 67416 92472
rect 184296 92420 184348 92472
rect 191840 92420 191892 92472
rect 217140 92420 217192 92472
rect 224868 92420 224920 92472
rect 227812 92420 227864 92472
rect 60648 92352 60700 92404
rect 79416 92352 79468 92404
rect 80612 92352 80664 92404
rect 99012 92352 99064 92404
rect 182088 92352 182140 92404
rect 202604 92352 202656 92404
rect 213276 92352 213328 92404
rect 226616 92352 226668 92404
rect 61844 90992 61896 91044
rect 70308 90992 70360 91044
rect 78956 90992 79008 91044
rect 111892 90992 111944 91044
rect 176568 90992 176620 91044
rect 195980 90992 196032 91044
rect 217140 90992 217192 91044
rect 246396 90992 246448 91044
rect 181996 90924 182048 90976
rect 194692 90924 194744 90976
rect 221372 90924 221424 90976
rect 225604 90924 225656 90976
rect 194692 90516 194744 90568
rect 195244 90516 195296 90568
rect 223764 90516 223816 90568
rect 224868 90516 224920 90568
rect 258724 90312 258776 90364
rect 291200 90312 291252 90364
rect 70308 89700 70360 89752
rect 73804 89700 73856 89752
rect 85212 89700 85264 89752
rect 93124 89700 93176 89752
rect 63408 89632 63460 89684
rect 100116 89632 100168 89684
rect 122196 89632 122248 89684
rect 217692 89632 217744 89684
rect 220636 89632 220688 89684
rect 245016 89632 245068 89684
rect 67272 89564 67324 89616
rect 94688 89564 94740 89616
rect 192024 89564 192076 89616
rect 199384 89564 199436 89616
rect 204444 89564 204496 89616
rect 205732 89564 205784 89616
rect 213368 88952 213420 89004
rect 235264 88952 235316 89004
rect 254584 88952 254636 89004
rect 583024 88952 583076 89004
rect 67456 88272 67508 88324
rect 100024 88272 100076 88324
rect 103520 88272 103572 88324
rect 214012 88272 214064 88324
rect 68928 88204 68980 88256
rect 80704 88204 80756 88256
rect 86132 88204 86184 88256
rect 111892 88204 111944 88256
rect 205548 88204 205600 88256
rect 207388 87592 207440 87644
rect 246304 87592 246356 87644
rect 89812 86912 89864 86964
rect 116676 86912 116728 86964
rect 218244 86912 218296 86964
rect 93308 86844 93360 86896
rect 124864 86844 124916 86896
rect 125508 86844 125560 86896
rect 205732 86844 205784 86896
rect 280252 86912 280304 86964
rect 580172 86912 580224 86964
rect 3516 85484 3568 85536
rect 53840 85484 53892 85536
rect 78404 85484 78456 85536
rect 106924 85484 106976 85536
rect 204996 85484 205048 85536
rect 214564 85484 214616 85536
rect 246488 85484 246540 85536
rect 198372 85416 198424 85468
rect 262864 85416 262916 85468
rect 88340 84124 88392 84176
rect 122196 84124 122248 84176
rect 169852 84124 169904 84176
rect 171048 84124 171100 84176
rect 193404 84124 193456 84176
rect 74540 84056 74592 84108
rect 101588 84056 101640 84108
rect 193404 83512 193456 83564
rect 226984 83512 227036 83564
rect 193036 83444 193088 83496
rect 259460 83444 259512 83496
rect 227076 82832 227128 82884
rect 241520 82832 241572 82884
rect 77300 82764 77352 82816
rect 108396 82764 108448 82816
rect 185584 82764 185636 82816
rect 229100 82764 229152 82816
rect 75920 82696 75972 82748
rect 94780 82696 94832 82748
rect 95148 82696 95200 82748
rect 186964 82696 187016 82748
rect 200120 82696 200172 82748
rect 201408 82696 201460 82748
rect 201408 82084 201460 82136
rect 214564 82084 214616 82136
rect 215392 81948 215444 82000
rect 216036 81948 216088 82000
rect 242164 82084 242216 82136
rect 85764 81336 85816 81388
rect 103612 81336 103664 81388
rect 109684 81336 109736 81388
rect 224960 81336 225012 81388
rect 69204 81268 69256 81320
rect 169852 81268 169904 81320
rect 201592 80656 201644 80708
rect 253204 80656 253256 80708
rect 201592 80044 201644 80096
rect 202144 80044 202196 80096
rect 54484 79976 54536 80028
rect 55128 79976 55180 80028
rect 188528 79976 188580 80028
rect 66076 79908 66128 79960
rect 112444 79908 112496 79960
rect 177488 79908 177540 79960
rect 227076 79908 227128 79960
rect 191564 79296 191616 79348
rect 280160 79296 280212 79348
rect 82820 78616 82872 78668
rect 178040 78616 178092 78668
rect 186964 78616 187016 78668
rect 190368 78616 190420 78668
rect 263600 78616 263652 78668
rect 264244 78616 264296 78668
rect 177396 78548 177448 78600
rect 230572 78548 230624 78600
rect 85580 77936 85632 77988
rect 105544 77936 105596 77988
rect 260104 77936 260156 77988
rect 295340 77936 295392 77988
rect 65524 77188 65576 77240
rect 102232 77188 102284 77240
rect 169024 77188 169076 77240
rect 229192 77188 229244 77240
rect 80704 76508 80756 76560
rect 100024 76508 100076 76560
rect 109040 76508 109092 76560
rect 135996 76508 136048 76560
rect 193128 76508 193180 76560
rect 338120 76508 338172 76560
rect 182824 75828 182876 75880
rect 230480 75828 230532 75880
rect 67640 75148 67692 75200
rect 171784 75148 171836 75200
rect 190184 75148 190236 75200
rect 248420 75148 248472 75200
rect 249064 75148 249116 75200
rect 85672 74468 85724 74520
rect 120080 74468 120132 74520
rect 213184 74468 213236 74520
rect 153936 74400 153988 74452
rect 237380 74400 237432 74452
rect 237380 73176 237432 73228
rect 238116 73176 238168 73228
rect 64788 73108 64840 73160
rect 190184 73108 190236 73160
rect 207020 73108 207072 73160
rect 258724 73176 258776 73228
rect 129648 73040 129700 73092
rect 227904 73040 227956 73092
rect 227904 71748 227956 71800
rect 228364 71748 228416 71800
rect 93124 71680 93176 71732
rect 106280 71680 106332 71732
rect 166264 71680 166316 71732
rect 231952 71680 232004 71732
rect 3516 71612 3568 71664
rect 95332 71612 95384 71664
rect 187608 71000 187660 71052
rect 288440 71000 288492 71052
rect 67548 70320 67600 70372
rect 180800 70320 180852 70372
rect 181444 70320 181496 70372
rect 160744 70252 160796 70304
rect 244280 70252 244332 70304
rect 244280 69844 244332 69896
rect 244924 69844 244976 69896
rect 222292 69028 222344 69080
rect 339500 69028 339552 69080
rect 124864 68960 124916 69012
rect 222200 68960 222252 69012
rect 222844 68960 222896 69012
rect 193312 68892 193364 68944
rect 193864 68892 193916 68944
rect 281540 68892 281592 68944
rect 88340 68280 88392 68332
rect 169760 68280 169812 68332
rect 97264 67532 97316 67584
rect 227720 67532 227772 67584
rect 65524 66852 65576 66904
rect 123484 66852 123536 66904
rect 190276 66852 190328 66904
rect 320272 66852 320324 66904
rect 71872 66172 71924 66224
rect 198004 66172 198056 66224
rect 200764 66172 200816 66224
rect 201408 66172 201460 66224
rect 250444 66172 250496 66224
rect 100024 66104 100076 66156
rect 207020 66104 207072 66156
rect 87052 64812 87104 64864
rect 215300 64812 215352 64864
rect 80060 64744 80112 64796
rect 205640 64744 205692 64796
rect 213184 64132 213236 64184
rect 333980 64132 334032 64184
rect 205640 63520 205692 63572
rect 206284 63520 206336 63572
rect 215300 63520 215352 63572
rect 215944 63520 215996 63572
rect 67732 63452 67784 63504
rect 193864 63452 193916 63504
rect 194784 62024 194836 62076
rect 287152 62024 287204 62076
rect 288348 62024 288400 62076
rect 86960 61956 87012 62008
rect 116032 61956 116084 62008
rect 216036 61956 216088 62008
rect 73804 61888 73856 61940
rect 194692 61888 194744 61940
rect 288348 61344 288400 61396
rect 345020 61344 345072 61396
rect 194692 60732 194744 60784
rect 195244 60732 195296 60784
rect 69112 60664 69164 60716
rect 194784 60664 194836 60716
rect 83464 60596 83516 60648
rect 107660 60596 107712 60648
rect 209780 60596 209832 60648
rect 211068 60596 211120 60648
rect 240876 60052 240928 60104
rect 278044 60052 278096 60104
rect 199384 59984 199436 60036
rect 244280 59984 244332 60036
rect 84844 59304 84896 59356
rect 211160 59304 211212 59356
rect 212448 59304 212500 59356
rect 70492 59236 70544 59288
rect 195980 59236 196032 59288
rect 196624 59236 196676 59288
rect 198740 58624 198792 58676
rect 240140 58624 240192 58676
rect 91008 57876 91060 57928
rect 219532 57876 219584 57928
rect 220084 57876 220136 57928
rect 212448 57808 212500 57860
rect 278688 57808 278740 57860
rect 278688 57196 278740 57248
rect 353300 57196 353352 57248
rect 74632 56516 74684 56568
rect 202144 56516 202196 56568
rect 211068 56516 211120 56568
rect 296720 56516 296772 56568
rect 298008 56516 298060 56568
rect 298008 55836 298060 55888
rect 322940 55836 322992 55888
rect 71780 54476 71832 54528
rect 151176 54476 151228 54528
rect 206284 54476 206336 54528
rect 232504 54476 232556 54528
rect 232596 54476 232648 54528
rect 324412 54476 324464 54528
rect 86960 53048 87012 53100
rect 153844 53048 153896 53100
rect 97264 51688 97316 51740
rect 131764 51688 131816 51740
rect 183468 51688 183520 51740
rect 281540 51688 281592 51740
rect 20 50328 72 50380
rect 97356 50328 97408 50380
rect 100760 50328 100812 50380
rect 146944 50328 146996 50380
rect 169576 50328 169628 50380
rect 335360 50328 335412 50380
rect 295984 49648 296036 49700
rect 296720 49648 296772 49700
rect 107660 49036 107712 49088
rect 126244 49036 126296 49088
rect 250536 49036 250588 49088
rect 260840 49036 260892 49088
rect 52460 48968 52512 49020
rect 133144 48968 133196 49020
rect 181444 48968 181496 49020
rect 251272 48968 251324 49020
rect 2872 47540 2924 47592
rect 147036 47540 147088 47592
rect 188436 46860 188488 46912
rect 580172 46860 580224 46912
rect 3516 46180 3568 46232
rect 54484 46180 54536 46232
rect 78680 46180 78732 46232
rect 142896 46180 142948 46232
rect 186136 43392 186188 43444
rect 249800 43392 249852 43444
rect 75920 42032 75972 42084
rect 137284 42032 137336 42084
rect 184756 42032 184808 42084
rect 298100 42032 298152 42084
rect 45560 40672 45612 40724
rect 156604 40672 156656 40724
rect 27712 39312 27764 39364
rect 159364 39312 159416 39364
rect 179236 39312 179288 39364
rect 309140 39312 309192 39364
rect 84200 37952 84252 38004
rect 122104 37952 122156 38004
rect 113180 37884 113232 37936
rect 160100 37884 160152 37936
rect 208400 37884 208452 37936
rect 278780 37884 278832 37936
rect 73160 36524 73212 36576
rect 155316 36524 155368 36576
rect 82820 35164 82872 35216
rect 145564 35164 145616 35216
rect 60740 33736 60792 33788
rect 174544 33736 174596 33788
rect 195244 33736 195296 33788
rect 311900 33736 311952 33788
rect 3516 33056 3568 33108
rect 53104 33056 53156 33108
rect 61752 32376 61804 32428
rect 125600 32376 125652 32428
rect 233884 32376 233936 32428
rect 316040 32376 316092 32428
rect 120080 29656 120132 29708
rect 157984 29656 158036 29708
rect 59360 29588 59412 29640
rect 130476 29588 130528 29640
rect 215944 29588 215996 29640
rect 266360 29588 266412 29640
rect 106280 28228 106332 28280
rect 162124 28228 162176 28280
rect 193864 28228 193916 28280
rect 291200 28228 291252 28280
rect 191656 26868 191708 26920
rect 322204 26868 322256 26920
rect 69112 25508 69164 25560
rect 152556 25508 152608 25560
rect 81440 24080 81492 24132
rect 164240 24080 164292 24132
rect 235264 24080 235316 24132
rect 287060 24080 287112 24132
rect 52552 22720 52604 22772
rect 161480 22720 161532 22772
rect 89720 21360 89772 21412
rect 148324 21360 148376 21412
rect 242164 21360 242216 21412
rect 284392 21360 284444 21412
rect 3424 20612 3476 20664
rect 90364 20612 90416 20664
rect 95240 19932 95292 19984
rect 151084 19932 151136 19984
rect 222844 19932 222896 19984
rect 302332 19932 302384 19984
rect 240784 18640 240836 18692
rect 276112 18640 276164 18692
rect 77300 18572 77352 18624
rect 155224 18572 155276 18624
rect 180156 18572 180208 18624
rect 242992 18572 243044 18624
rect 63500 17212 63552 17264
rect 177304 17212 177356 17264
rect 238024 17212 238076 17264
rect 269764 17212 269816 17264
rect 244924 15852 244976 15904
rect 256700 15852 256752 15904
rect 270408 15852 270460 15904
rect 330392 15852 330444 15904
rect 93124 14424 93176 14476
rect 137376 14424 137428 14476
rect 253204 14424 253256 14476
rect 321560 14424 321612 14476
rect 102232 13132 102284 13184
rect 159456 13132 159508 13184
rect 61568 13064 61620 13116
rect 140044 13064 140096 13116
rect 201408 13064 201460 13116
rect 340972 13064 341024 13116
rect 75184 11704 75236 11756
rect 135904 11704 135956 11756
rect 246396 11704 246448 11756
rect 291936 11704 291988 11756
rect 58440 10276 58492 10328
rect 138664 10276 138716 10328
rect 198004 10276 198056 10328
rect 342904 10276 342956 10328
rect 9956 8916 10008 8968
rect 184204 8916 184256 8968
rect 196624 8916 196676 8968
rect 258264 8916 258316 8968
rect 258724 8916 258776 8968
rect 274824 8916 274876 8968
rect 97448 7624 97500 7676
rect 141424 7624 141476 7676
rect 44272 7556 44324 7608
rect 97264 7556 97316 7608
rect 220084 7556 220136 7608
rect 346400 7556 346452 7608
rect 3424 6808 3476 6860
rect 7564 6808 7616 6860
rect 191748 6128 191800 6180
rect 293684 6128 293736 6180
rect 305644 5516 305696 5568
rect 309048 5516 309100 5568
rect 349804 5516 349856 5568
rect 350540 5516 350592 5568
rect 323584 4904 323636 4956
rect 326804 4904 326856 4956
rect 238116 4836 238168 4888
rect 239312 4836 239364 4888
rect 65524 4768 65576 4820
rect 149704 4768 149756 4820
rect 228364 4768 228416 4820
rect 278320 4768 278372 4820
rect 342996 4768 343048 4820
rect 346952 4768 347004 4820
rect 134524 4156 134576 4208
rect 136456 4156 136508 4208
rect 309784 4156 309836 4208
rect 315028 4156 315080 4208
rect 317328 4156 317380 4208
rect 321652 4156 321704 4208
rect 337476 4156 337528 4208
rect 340880 4156 340932 4208
rect 63224 4088 63276 4140
rect 65432 4088 65484 4140
rect 267004 4088 267056 4140
rect 267740 4088 267792 4140
rect 333888 4088 333940 4140
rect 335452 4088 335504 4140
rect 150624 3612 150676 3664
rect 152464 3612 152516 3664
rect 2780 3476 2832 3528
rect 4068 3476 4120 3528
rect 11060 3476 11112 3528
rect 12348 3476 12400 3528
rect 37188 3476 37240 3528
rect 47584 3476 47636 3528
rect 69020 3476 69072 3528
rect 70308 3476 70360 3528
rect 77392 3476 77444 3528
rect 79324 3476 79376 3528
rect 85580 3476 85632 3528
rect 86868 3476 86920 3528
rect 91560 3476 91612 3528
rect 98644 3476 98696 3528
rect 102140 3476 102192 3528
rect 103336 3476 103388 3528
rect 140044 3476 140096 3528
rect 148508 3544 148560 3596
rect 251180 3544 251232 3596
rect 252376 3544 252428 3596
rect 276020 3544 276072 3596
rect 277124 3544 277176 3596
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 232504 3476 232556 3528
rect 242900 3476 242952 3528
rect 287704 3476 287756 3528
rect 290188 3476 290240 3528
rect 291936 3476 291988 3528
rect 294880 3476 294932 3528
rect 299480 3476 299532 3528
rect 300768 3476 300820 3528
rect 309140 3476 309192 3528
rect 310244 3476 310296 3528
rect 319720 3476 319772 3528
rect 320180 3476 320232 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 20628 3408 20680 3460
rect 36544 3408 36596 3460
rect 51356 3408 51408 3460
rect 75184 3408 75236 3460
rect 80888 3408 80940 3460
rect 93124 3408 93176 3460
rect 99840 3408 99892 3460
rect 108304 3408 108356 3460
rect 104532 3340 104584 3392
rect 142804 3408 142856 3460
rect 214564 3408 214616 3460
rect 246396 3408 246448 3460
rect 298744 3408 298796 3460
rect 305552 3408 305604 3460
rect 322204 3408 322256 3460
rect 329196 3408 329248 3460
rect 334716 3408 334768 3460
rect 344560 3408 344612 3460
rect 278044 3340 278096 3392
rect 283104 3340 283156 3392
rect 346400 3340 346452 3392
rect 349252 3340 349304 3392
rect 260656 3272 260708 3324
rect 262312 3272 262364 3324
rect 327724 3272 327776 3324
rect 332692 3272 332744 3324
rect 338764 3272 338816 3324
rect 342168 3272 342220 3324
rect 348056 3272 348108 3324
rect 351920 3272 351972 3324
rect 581000 3272 581052 3324
rect 582564 3272 582616 3324
rect 269764 3068 269816 3120
rect 272432 3068 272484 3120
rect 299664 3068 299716 3120
rect 302240 3068 302292 3120
rect 246304 2932 246356 2984
rect 247592 2932 247644 2984
rect 289084 2932 289136 2984
rect 292580 2932 292632 2984
rect 307024 2932 307076 2984
rect 307944 2932 307996 2984
rect 351644 2864 351696 2916
rect 353300 2864 353352 2916
rect 7656 2048 7708 2100
rect 22744 2048 22796 2100
rect 93952 2048 94004 2100
rect 130384 2048 130436 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702506 8156 703520
rect 24320 702642 24348 703520
rect 24308 702636 24360 702642
rect 24308 702578 24360 702584
rect 8116 702500 8168 702506
rect 8116 702442 8168 702448
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 33784 683188 33836 683194
rect 33784 683130 33836 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 15844 670744 15896 670750
rect 15844 670686 15896 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3332 580984 3384 580990
rect 3332 580926 3384 580932
rect 3344 580009 3372 580926
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3436 576842 3464 632023
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 576836 3476 576842
rect 3424 576778 3476 576784
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553722 3464 553823
rect 3424 553716 3476 553722
rect 3424 553658 3476 553664
rect 7564 553716 7616 553722
rect 7564 553658 7616 553664
rect 7576 538218 7604 553658
rect 15856 541686 15884 670686
rect 33796 543726 33824 683130
rect 40052 588606 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 67640 702568 67692 702574
rect 67640 702510 67692 702516
rect 57244 618316 57296 618322
rect 57244 618258 57296 618264
rect 40040 588600 40092 588606
rect 40040 588542 40092 588548
rect 55128 582480 55180 582486
rect 55128 582422 55180 582428
rect 53748 579692 53800 579698
rect 53748 579634 53800 579640
rect 39304 565888 39356 565894
rect 39304 565830 39356 565836
rect 52368 565888 52420 565894
rect 52368 565830 52420 565836
rect 33784 543720 33836 543726
rect 33784 543662 33836 543668
rect 15844 541680 15896 541686
rect 15844 541622 15896 541628
rect 7564 538212 7616 538218
rect 7564 538154 7616 538160
rect 39316 536110 39344 565830
rect 50988 543788 51040 543794
rect 50988 543730 51040 543736
rect 39948 541680 40000 541686
rect 39948 541622 40000 541628
rect 39960 541006 39988 541622
rect 39948 541000 40000 541006
rect 39948 540942 40000 540948
rect 39304 536104 39356 536110
rect 39304 536046 39356 536052
rect 3424 528488 3476 528494
rect 3424 528430 3476 528436
rect 3436 527921 3464 528430
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3424 522300 3476 522306
rect 3424 522242 3476 522248
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 2780 514762 2832 514768
rect 3436 501809 3464 522242
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 475386 3372 475623
rect 3332 475380 3384 475386
rect 3332 475322 3384 475328
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 4816 439550 4844 514762
rect 35164 478168 35216 478174
rect 35164 478110 35216 478116
rect 35176 475386 35204 478110
rect 35164 475380 35216 475386
rect 35164 475322 35216 475328
rect 17224 462392 17276 462398
rect 17224 462334 17276 462340
rect 4804 439544 4856 439550
rect 4804 439486 4856 439492
rect 15844 436144 15896 436150
rect 15844 436086 15896 436092
rect 3424 434784 3476 434790
rect 3424 434726 3476 434732
rect 3436 423609 3464 434726
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 2778 410544 2834 410553
rect 2778 410479 2834 410488
rect 2792 410242 2820 410479
rect 2780 410236 2832 410242
rect 2780 410178 2832 410184
rect 4804 410236 4856 410242
rect 4804 410178 4856 410184
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 380905 3464 397423
rect 4816 391270 4844 410178
rect 4804 391264 4856 391270
rect 4804 391206 4856 391212
rect 3516 383716 3568 383722
rect 3516 383658 3568 383664
rect 3422 380896 3478 380905
rect 3422 380831 3478 380840
rect 3528 371385 3556 383658
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 15200 344344 15252 344350
rect 15200 344286 15252 344292
rect 11058 333296 11114 333305
rect 11058 333231 11114 333240
rect 8300 329112 8352 329118
rect 8300 329054 8352 329060
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 264926 3464 306167
rect 4080 305182 4108 319223
rect 5538 306504 5594 306513
rect 5538 306439 5594 306448
rect 4068 305176 4120 305182
rect 4068 305118 4120 305124
rect 4158 294536 4214 294545
rect 4158 294471 4214 294480
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3424 264920 3476 264926
rect 3424 264862 3476 264868
rect 4068 261520 4120 261526
rect 4068 261462 4120 261468
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3436 254153 3464 255206
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 241120 3476 241126
rect 3422 241088 3424 241097
rect 3476 241088 3478 241097
rect 3422 241023 3478 241032
rect 4080 219434 4108 261462
rect 3988 219406 4108 219434
rect 2778 215928 2834 215937
rect 2778 215863 2834 215872
rect 1400 178696 1452 178702
rect 1400 178638 1452 178644
rect 20 50380 72 50386
rect 20 50322 72 50328
rect 32 16574 60 50322
rect 1412 16574 1440 178638
rect 32 16546 152 16574
rect 1412 16546 1716 16574
rect 124 490 152 16546
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 16546
rect 2792 3534 2820 215863
rect 3988 214985 4016 219406
rect 3974 214976 4030 214985
rect 3974 214911 3976 214920
rect 4028 214911 4030 214920
rect 3976 214882 4028 214888
rect 3332 202224 3384 202230
rect 3332 202166 3384 202172
rect 3344 201929 3372 202166
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 2872 162920 2924 162926
rect 2870 162888 2872 162897
rect 2924 162888 2926 162897
rect 2870 162823 2926 162832
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 146946 3188 149767
rect 3148 146940 3200 146946
rect 3148 146882 3200 146888
rect 2872 137964 2924 137970
rect 2872 137906 2924 137912
rect 2884 136785 2912 137906
rect 2870 136776 2926 136785
rect 2870 136711 2926 136720
rect 3422 134872 3478 134881
rect 3422 134807 3478 134816
rect 2872 110832 2924 110838
rect 2872 110774 2924 110780
rect 2884 110673 2912 110774
rect 2870 110664 2926 110673
rect 2870 110599 2926 110608
rect 3054 97608 3110 97617
rect 3054 97543 3110 97552
rect 3068 96694 3096 97543
rect 3056 96688 3108 96694
rect 3056 96630 3108 96636
rect 3436 58585 3464 134807
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 3568 71632 3570 71641
rect 3514 71567 3570 71576
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 2872 47592 2924 47598
rect 2872 47534 2924 47540
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 47534
rect 3516 46232 3568 46238
rect 3516 46174 3568 46180
rect 3528 45529 3556 46174
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 294471
rect 4804 162920 4856 162926
rect 4804 162862 4856 162868
rect 4816 146266 4844 162862
rect 4804 146260 4856 146266
rect 4804 146202 4856 146208
rect 4804 135312 4856 135318
rect 4804 135254 4856 135260
rect 4816 110838 4844 135254
rect 4804 110832 4856 110838
rect 4804 110774 4856 110780
rect 5552 16574 5580 306439
rect 7564 305176 7616 305182
rect 7564 305118 7616 305124
rect 7576 279478 7604 305118
rect 7564 279472 7616 279478
rect 7564 279414 7616 279420
rect 7564 262268 7616 262274
rect 7564 262210 7616 262216
rect 7576 241126 7604 262210
rect 7564 241120 7616 241126
rect 7564 241062 7616 241068
rect 7564 214940 7616 214946
rect 7564 214882 7616 214888
rect 7576 113830 7604 214882
rect 7564 113824 7616 113830
rect 7564 113766 7616 113772
rect 7564 106344 7616 106350
rect 7564 106286 7616 106292
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 480 4108 3470
rect 5276 480 5304 16546
rect 6012 490 6040 16546
rect 7576 6866 7604 106286
rect 8312 16574 8340 329054
rect 8312 16546 8800 16574
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 6288 598 6500 626
rect 6288 490 6316 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 462 6316 490
rect 6472 480 6500 598
rect 7668 480 7696 2042
rect 8772 480 8800 16546
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 480 9996 8910
rect 11072 3534 11100 333231
rect 12438 300112 12494 300121
rect 12438 300047 12494 300056
rect 11150 298752 11206 298761
rect 11150 298687 11206 298696
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 298687
rect 12452 16574 12480 300047
rect 13820 207664 13872 207670
rect 13820 207606 13872 207612
rect 13832 16574 13860 207606
rect 15212 16574 15240 344286
rect 15856 319462 15884 436086
rect 17236 389230 17264 462334
rect 35176 391338 35204 475322
rect 39856 408468 39908 408474
rect 39856 408410 39908 408416
rect 36544 397520 36596 397526
rect 36544 397462 36596 397468
rect 35164 391332 35216 391338
rect 35164 391274 35216 391280
rect 17224 389224 17276 389230
rect 17224 389166 17276 389172
rect 36556 358766 36584 397462
rect 36544 358760 36596 358766
rect 36544 358702 36596 358708
rect 24858 347032 24914 347041
rect 24858 346967 24914 346976
rect 20718 338736 20774 338745
rect 20718 338671 20774 338680
rect 17958 335472 18014 335481
rect 17958 335407 18014 335416
rect 16578 331800 16634 331809
rect 16578 331735 16634 331744
rect 15844 319456 15896 319462
rect 15844 319398 15896 319404
rect 16592 16574 16620 331735
rect 17972 16574 18000 335407
rect 19338 155272 19394 155281
rect 19338 155207 19394 155216
rect 19352 16574 19380 155207
rect 20732 16574 20760 338671
rect 22742 334112 22798 334121
rect 22742 334047 22798 334056
rect 22098 324456 22154 324465
rect 22098 324391 22154 324400
rect 22112 16574 22140 324391
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 17972 16546 18276 16574
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12360 480 12388 3470
rect 13556 480 13584 16546
rect 14292 490 14320 16546
rect 14568 598 14780 626
rect 14568 490 14596 598
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 462 14596 490
rect 14752 480 14780 598
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 18248 480 18276 16546
rect 19444 480 19472 16546
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20640 480 20668 3402
rect 21836 480 21864 16546
rect 22572 490 22600 16546
rect 22756 2106 22784 334047
rect 22836 292596 22888 292602
rect 22836 292538 22888 292544
rect 22848 241466 22876 292538
rect 22836 241460 22888 241466
rect 22836 241402 22888 241408
rect 23480 196648 23532 196654
rect 23480 196590 23532 196596
rect 23492 16574 23520 196590
rect 24872 16574 24900 346967
rect 35164 345092 35216 345098
rect 35164 345034 35216 345040
rect 30378 330440 30434 330449
rect 30378 330375 30434 330384
rect 27618 327720 27674 327729
rect 27618 327655 27674 327664
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 22744 2100 22796 2106
rect 22744 2042 22796 2048
rect 22848 598 23060 626
rect 22848 490 22876 598
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 462 22876 490
rect 23032 480 23060 598
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 27632 6914 27660 327655
rect 28998 322144 29054 322153
rect 28998 322079 29054 322088
rect 27712 39364 27764 39370
rect 27712 39306 27764 39312
rect 27724 16574 27752 39306
rect 29012 16574 29040 322079
rect 30392 16574 30420 330375
rect 33140 326392 33192 326398
rect 33140 326334 33192 326340
rect 32404 316736 32456 316742
rect 32404 316678 32456 316684
rect 32416 264926 32444 316678
rect 32404 264920 32456 264926
rect 32404 264862 32456 264868
rect 32416 253230 32444 264862
rect 32404 253224 32456 253230
rect 32404 253166 32456 253172
rect 31758 233880 31814 233889
rect 31758 233815 31814 233824
rect 31772 16574 31800 233815
rect 33152 16574 33180 326334
rect 34520 301504 34572 301510
rect 34520 301446 34572 301452
rect 34532 16574 34560 301446
rect 35176 288386 35204 345034
rect 37278 318880 37334 318889
rect 37278 318815 37334 318824
rect 36542 296032 36598 296041
rect 36542 295967 36598 295976
rect 35164 288380 35216 288386
rect 35164 288322 35216 288328
rect 35808 279472 35860 279478
rect 35808 279414 35860 279420
rect 35820 156670 35848 279414
rect 35808 156664 35860 156670
rect 35808 156606 35860 156612
rect 35898 30968 35954 30977
rect 35898 30903 35954 30912
rect 35912 16574 35940 30903
rect 27724 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 34532 16546 34836 16574
rect 35912 16546 36032 16574
rect 27632 6886 27752 6914
rect 26514 6216 26570 6225
rect 26514 6151 26570 6160
rect 26528 480 26556 6151
rect 27724 480 27752 6886
rect 28460 490 28488 16546
rect 28736 598 28948 626
rect 28736 490 28764 598
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28460 462 28764 490
rect 28920 480 28948 598
rect 30116 480 30144 16546
rect 30852 490 30880 16546
rect 31128 598 31340 626
rect 31128 490 31156 598
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 462 31156 490
rect 31312 480 31340 598
rect 31956 490 31984 16546
rect 32232 598 32444 626
rect 32232 490 32260 598
rect 31270 -960 31382 480
rect 31956 462 32260 490
rect 32416 480 32444 598
rect 33612 480 33640 16546
rect 34808 480 34836 16546
rect 36004 480 36032 16546
rect 36556 3466 36584 295967
rect 37292 16574 37320 318815
rect 37924 284368 37976 284374
rect 37924 284310 37976 284316
rect 37936 267714 37964 284310
rect 37924 267708 37976 267714
rect 37924 267650 37976 267656
rect 39868 255921 39896 408410
rect 39960 386306 39988 540942
rect 43444 538348 43496 538354
rect 43444 538290 43496 538296
rect 43456 478174 43484 538290
rect 48228 532024 48280 532030
rect 48228 531966 48280 531972
rect 43444 478168 43496 478174
rect 43444 478110 43496 478116
rect 48240 455530 48268 531966
rect 51000 511970 51028 543730
rect 50988 511964 51040 511970
rect 50988 511906 51040 511912
rect 48228 455524 48280 455530
rect 48228 455466 48280 455472
rect 40684 448588 40736 448594
rect 40684 448530 40736 448536
rect 40696 389298 40724 448530
rect 41328 425740 41380 425746
rect 41328 425682 41380 425688
rect 40684 389292 40736 389298
rect 40684 389234 40736 389240
rect 39948 386300 40000 386306
rect 39948 386242 40000 386248
rect 40038 323640 40094 323649
rect 40038 323575 40094 323584
rect 39946 260128 40002 260137
rect 39946 260063 40002 260072
rect 39854 255912 39910 255921
rect 39854 255847 39910 255856
rect 38660 202156 38712 202162
rect 38660 202098 38712 202104
rect 38672 16574 38700 202098
rect 39960 111110 39988 260063
rect 39948 111104 40000 111110
rect 39948 111046 40000 111052
rect 40052 16574 40080 323575
rect 41340 269822 41368 425682
rect 48136 420980 48188 420986
rect 48136 420922 48188 420928
rect 44088 410576 44140 410582
rect 44088 410518 44140 410524
rect 41420 336864 41472 336870
rect 41420 336806 41472 336812
rect 41328 269816 41380 269822
rect 41328 269758 41380 269764
rect 41432 16574 41460 336806
rect 43444 280220 43496 280226
rect 43444 280162 43496 280168
rect 43456 255270 43484 280162
rect 43996 260160 44048 260166
rect 43996 260102 44048 260108
rect 43444 255264 43496 255270
rect 43444 255206 43496 255212
rect 43444 234660 43496 234666
rect 43444 234602 43496 234608
rect 43456 189038 43484 234602
rect 43444 189032 43496 189038
rect 43444 188974 43496 188980
rect 42798 188320 42854 188329
rect 42798 188255 42854 188264
rect 42812 16574 42840 188255
rect 44008 111790 44036 260102
rect 44100 257378 44128 410518
rect 48148 387025 48176 420922
rect 48240 408474 48268 455466
rect 51000 440881 51028 511906
rect 52380 460934 52408 565830
rect 53656 536104 53708 536110
rect 53656 536046 53708 536052
rect 52196 460906 52408 460934
rect 52196 458318 52224 460906
rect 52184 458312 52236 458318
rect 52184 458254 52236 458260
rect 50986 440872 51042 440881
rect 50986 440807 51042 440816
rect 50988 422340 51040 422346
rect 50988 422282 51040 422288
rect 50896 416084 50948 416090
rect 50896 416026 50948 416032
rect 49608 408536 49660 408542
rect 49608 408478 49660 408484
rect 48228 408468 48280 408474
rect 48228 408410 48280 408416
rect 48134 387016 48190 387025
rect 48134 386951 48190 386960
rect 46756 376032 46808 376038
rect 46756 375974 46808 375980
rect 44180 342916 44232 342922
rect 44180 342858 44232 342864
rect 44088 257372 44140 257378
rect 44088 257314 44140 257320
rect 43996 111784 44048 111790
rect 43996 111726 44048 111732
rect 44192 16574 44220 342858
rect 45468 288448 45520 288454
rect 45468 288390 45520 288396
rect 45480 185638 45508 288390
rect 46768 238746 46796 375974
rect 48148 265033 48176 386951
rect 48228 371884 48280 371890
rect 48228 371826 48280 371832
rect 48134 265024 48190 265033
rect 48134 264959 48190 264968
rect 46846 255912 46902 255921
rect 46846 255847 46902 255856
rect 46860 254590 46888 255847
rect 46848 254584 46900 254590
rect 46848 254526 46900 254532
rect 46756 238740 46808 238746
rect 46756 238682 46808 238688
rect 45468 185632 45520 185638
rect 45468 185574 45520 185580
rect 46860 105602 46888 254526
rect 48136 250504 48188 250510
rect 48136 250446 48188 250452
rect 47584 218816 47636 218822
rect 47584 218758 47636 218764
rect 46848 105596 46900 105602
rect 46848 105538 46900 105544
rect 46938 43480 46994 43489
rect 46938 43415 46994 43424
rect 45560 40724 45612 40730
rect 45560 40666 45612 40672
rect 45572 16574 45600 40666
rect 46952 16574 46980 43415
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 42812 16546 43116 16574
rect 44192 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 36544 3460 36596 3466
rect 36544 3402 36596 3408
rect 37200 480 37228 3470
rect 38396 480 38424 16546
rect 39132 490 39160 16546
rect 39408 598 39620 626
rect 39408 490 39436 598
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 462 39436 490
rect 39592 480 39620 598
rect 40236 490 40264 16546
rect 40512 598 40724 626
rect 40512 490 40540 598
rect 39550 -960 39662 480
rect 40236 462 40540 490
rect 40696 480 40724 598
rect 41892 480 41920 16546
rect 43088 480 43116 16546
rect 44272 7608 44324 7614
rect 44272 7550 44324 7556
rect 44284 480 44312 7550
rect 45020 490 45048 16546
rect 45296 598 45508 626
rect 45296 490 45324 598
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 462 45324 490
rect 45480 480 45508 598
rect 46676 480 46704 16546
rect 47412 490 47440 16546
rect 47596 3534 47624 218758
rect 48148 151814 48176 250446
rect 48240 240106 48268 371826
rect 49516 262268 49568 262274
rect 49516 262210 49568 262216
rect 48228 240100 48280 240106
rect 48228 240042 48280 240048
rect 49528 227798 49556 262210
rect 49620 256018 49648 408478
rect 50908 289105 50936 416026
rect 50894 289096 50950 289105
rect 50894 289031 50950 289040
rect 50804 269816 50856 269822
rect 50804 269758 50856 269764
rect 50816 268025 50844 269758
rect 50802 268016 50858 268025
rect 50802 267951 50858 267960
rect 50710 265024 50766 265033
rect 50710 264959 50766 264968
rect 49608 256012 49660 256018
rect 49608 255954 49660 255960
rect 49516 227792 49568 227798
rect 49516 227734 49568 227740
rect 49700 189780 49752 189786
rect 49700 189722 49752 189728
rect 48320 186992 48372 186998
rect 48320 186934 48372 186940
rect 48148 151786 48268 151814
rect 48240 147694 48268 151786
rect 48228 147688 48280 147694
rect 48228 147630 48280 147636
rect 48240 109070 48268 147630
rect 48228 109064 48280 109070
rect 48228 109006 48280 109012
rect 48332 16574 48360 186934
rect 49712 16574 49740 189722
rect 50724 171134 50752 264959
rect 50816 224262 50844 267951
rect 50908 261594 50936 289031
rect 51000 267714 51028 422282
rect 52196 411262 52224 458254
rect 52274 434752 52330 434761
rect 52274 434687 52330 434696
rect 52184 411256 52236 411262
rect 52184 411198 52236 411204
rect 52196 410582 52224 411198
rect 52184 410576 52236 410582
rect 52184 410518 52236 410524
rect 52288 308417 52316 434687
rect 52368 432676 52420 432682
rect 52368 432618 52420 432624
rect 52274 308408 52330 308417
rect 52274 308343 52330 308352
rect 52184 285796 52236 285802
rect 52184 285738 52236 285744
rect 50988 267708 51040 267714
rect 50988 267650 51040 267656
rect 50896 261588 50948 261594
rect 50896 261530 50948 261536
rect 50988 236700 51040 236706
rect 50988 236642 51040 236648
rect 50804 224256 50856 224262
rect 50804 224198 50856 224204
rect 51000 212498 51028 236642
rect 50988 212492 51040 212498
rect 50988 212434 51040 212440
rect 50724 171106 50936 171134
rect 50908 150521 50936 171106
rect 50894 150512 50950 150521
rect 50894 150447 50950 150456
rect 50908 115938 50936 150447
rect 50896 115932 50948 115938
rect 50896 115874 50948 115880
rect 51000 88233 51028 212434
rect 52196 132462 52224 285738
rect 52288 277370 52316 308343
rect 52380 283626 52408 432618
rect 53668 432614 53696 536046
rect 53760 434042 53788 579634
rect 53748 434036 53800 434042
rect 53748 433978 53800 433984
rect 53656 432608 53708 432614
rect 53656 432550 53708 432556
rect 53668 403646 53696 432550
rect 53748 423700 53800 423706
rect 53748 423642 53800 423648
rect 53656 403640 53708 403646
rect 53656 403582 53708 403588
rect 53656 398880 53708 398886
rect 53656 398822 53708 398828
rect 53564 285728 53616 285734
rect 53564 285670 53616 285676
rect 52368 283620 52420 283626
rect 52368 283562 52420 283568
rect 52276 277364 52328 277370
rect 52276 277306 52328 277312
rect 53470 270736 53526 270745
rect 53470 270671 53526 270680
rect 52276 269068 52328 269074
rect 52276 269010 52328 269016
rect 52288 149705 52316 269010
rect 52274 149696 52330 149705
rect 52274 149631 52330 149640
rect 52184 132456 52236 132462
rect 52184 132398 52236 132404
rect 52288 118658 52316 149631
rect 53484 139505 53512 270671
rect 53576 141409 53604 285670
rect 53668 249082 53696 398822
rect 53760 269074 53788 423642
rect 55036 414044 55088 414050
rect 55036 413986 55088 413992
rect 54300 284980 54352 284986
rect 54300 284922 54352 284928
rect 54312 284374 54340 284922
rect 54300 284368 54352 284374
rect 54300 284310 54352 284316
rect 54852 284368 54904 284374
rect 54852 284310 54904 284316
rect 53748 269068 53800 269074
rect 53748 269010 53800 269016
rect 53840 257372 53892 257378
rect 53840 257314 53892 257320
rect 53852 256766 53880 257314
rect 53840 256760 53892 256766
rect 53840 256702 53892 256708
rect 53656 249076 53708 249082
rect 53656 249018 53708 249024
rect 53656 247104 53708 247110
rect 53656 247046 53708 247052
rect 53668 220114 53696 247046
rect 54864 233170 54892 284310
rect 55048 262857 55076 413986
rect 55140 413302 55168 582422
rect 56416 553444 56468 553450
rect 56416 553386 56468 553392
rect 56428 416090 56456 553386
rect 57256 536790 57284 618258
rect 66168 611380 66220 611386
rect 66168 611322 66220 611328
rect 65984 585200 66036 585206
rect 65984 585142 66036 585148
rect 61936 579760 61988 579766
rect 61936 579702 61988 579708
rect 59268 567248 59320 567254
rect 59268 567190 59320 567196
rect 57796 539640 57848 539646
rect 57796 539582 57848 539588
rect 57244 536784 57296 536790
rect 57244 536726 57296 536732
rect 57702 533352 57758 533361
rect 57702 533287 57758 533296
rect 56506 425096 56562 425105
rect 56506 425031 56562 425040
rect 56416 416084 56468 416090
rect 56416 416026 56468 416032
rect 55128 413296 55180 413302
rect 55128 413238 55180 413244
rect 55034 262848 55090 262857
rect 55034 262783 55090 262792
rect 55140 258738 55168 413238
rect 56416 283620 56468 283626
rect 56416 283562 56468 283568
rect 55128 258732 55180 258738
rect 55128 258674 55180 258680
rect 54944 256760 54996 256766
rect 54944 256702 54996 256708
rect 54852 233164 54904 233170
rect 54852 233106 54904 233112
rect 53656 220108 53708 220114
rect 53656 220050 53708 220056
rect 53562 141400 53618 141409
rect 53562 141335 53618 141344
rect 53470 139496 53526 139505
rect 53470 139431 53526 139440
rect 53104 135380 53156 135386
rect 53104 135322 53156 135328
rect 52276 118652 52328 118658
rect 52276 118594 52328 118600
rect 50986 88224 51042 88233
rect 50986 88159 51042 88168
rect 52460 49020 52512 49026
rect 52460 48962 52512 48968
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 47688 598 47900 626
rect 47688 490 47716 598
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 462 47716 490
rect 47872 480 47900 598
rect 48516 490 48544 16546
rect 48792 598 49004 626
rect 48792 490 48820 598
rect 47830 -960 47942 480
rect 48516 462 48820 490
rect 48976 480 49004 598
rect 50172 480 50200 16546
rect 52472 6914 52500 48962
rect 53116 33114 53144 135322
rect 53668 99346 53696 220050
rect 54956 201482 54984 256702
rect 55036 251864 55088 251870
rect 55036 251806 55088 251812
rect 54944 201476 54996 201482
rect 54944 201418 54996 201424
rect 54956 143585 54984 201418
rect 54942 143576 54998 143585
rect 54942 143511 54998 143520
rect 53746 139496 53802 139505
rect 53746 139431 53802 139440
rect 53760 121446 53788 139431
rect 53748 121440 53800 121446
rect 53748 121382 53800 121388
rect 53840 109064 53892 109070
rect 53840 109006 53892 109012
rect 53656 99340 53708 99346
rect 53656 99282 53708 99288
rect 53852 85542 53880 109006
rect 54956 109002 54984 143511
rect 55048 138145 55076 251806
rect 55128 227792 55180 227798
rect 55128 227734 55180 227740
rect 55034 138136 55090 138145
rect 55034 138071 55090 138080
rect 54944 108996 54996 109002
rect 54944 108938 54996 108944
rect 55048 103426 55076 138071
rect 55140 113150 55168 227734
rect 56428 171134 56456 283562
rect 56520 270502 56548 425031
rect 57716 395350 57744 533287
rect 57704 395344 57756 395350
rect 57704 395286 57756 395292
rect 57704 392012 57756 392018
rect 57704 391954 57756 391960
rect 57716 365634 57744 391954
rect 57808 389201 57836 539582
rect 59176 533384 59228 533390
rect 59176 533326 59228 533332
rect 57888 406428 57940 406434
rect 57888 406370 57940 406376
rect 57794 389192 57850 389201
rect 57794 389127 57850 389136
rect 57704 365628 57756 365634
rect 57704 365570 57756 365576
rect 56508 270496 56560 270502
rect 56508 270438 56560 270444
rect 56600 253972 56652 253978
rect 56600 253914 56652 253920
rect 56612 252498 56640 253914
rect 56520 252470 56640 252498
rect 56520 222902 56548 252470
rect 57716 244254 57744 365570
rect 57794 275224 57850 275233
rect 57794 275159 57850 275168
rect 57704 244248 57756 244254
rect 57704 244190 57756 244196
rect 57704 242956 57756 242962
rect 57704 242898 57756 242904
rect 56508 222896 56560 222902
rect 56508 222838 56560 222844
rect 56336 171106 56456 171134
rect 56336 170406 56364 171106
rect 56324 170400 56376 170406
rect 56324 170342 56376 170348
rect 56336 132394 56364 170342
rect 56416 158024 56468 158030
rect 56416 157966 56468 157972
rect 56324 132388 56376 132394
rect 56324 132330 56376 132336
rect 55128 113144 55180 113150
rect 55128 113086 55180 113092
rect 55036 103420 55088 103426
rect 55036 103362 55088 103368
rect 55128 101448 55180 101454
rect 55128 101390 55180 101396
rect 53840 85536 53892 85542
rect 53840 85478 53892 85484
rect 55140 80034 55168 101390
rect 56428 90953 56456 157966
rect 56520 104854 56548 222838
rect 57716 209098 57744 242898
rect 57704 209092 57756 209098
rect 57704 209034 57756 209040
rect 56508 104848 56560 104854
rect 56508 104790 56560 104796
rect 57716 95198 57744 209034
rect 57808 140826 57836 275159
rect 57900 254726 57928 406370
rect 59084 400240 59136 400246
rect 59084 400182 59136 400188
rect 59096 287054 59124 400182
rect 59188 388482 59216 533326
rect 59280 528562 59308 567190
rect 60648 558952 60700 558958
rect 60648 558894 60700 558900
rect 59268 528556 59320 528562
rect 59268 528498 59320 528504
rect 59268 436212 59320 436218
rect 59268 436154 59320 436160
rect 59176 388476 59228 388482
rect 59176 388418 59228 388424
rect 59096 287026 59216 287054
rect 59188 284617 59216 287026
rect 59174 284608 59230 284617
rect 59174 284543 59230 284552
rect 58900 284368 58952 284374
rect 58900 284310 58952 284316
rect 57888 254720 57940 254726
rect 57888 254662 57940 254668
rect 57900 253978 57928 254662
rect 57888 253972 57940 253978
rect 57888 253914 57940 253920
rect 57888 241528 57940 241534
rect 57888 241470 57940 241476
rect 57796 140820 57848 140826
rect 57796 140762 57848 140768
rect 57808 124914 57836 140762
rect 57796 124908 57848 124914
rect 57796 124850 57848 124856
rect 57704 95192 57756 95198
rect 57704 95134 57756 95140
rect 57900 93838 57928 241470
rect 58912 137290 58940 284310
rect 59084 270496 59136 270502
rect 59084 270438 59136 270444
rect 59096 269822 59124 270438
rect 59084 269816 59136 269822
rect 59084 269758 59136 269764
rect 58992 258732 59044 258738
rect 58992 258674 59044 258680
rect 59004 230489 59032 258674
rect 58990 230480 59046 230489
rect 58990 230415 59046 230424
rect 59096 153241 59124 269758
rect 59188 250073 59216 284543
rect 59280 283257 59308 436154
rect 60556 429276 60608 429282
rect 60556 429218 60608 429224
rect 60464 291848 60516 291854
rect 60464 291790 60516 291796
rect 59266 283248 59322 283257
rect 59266 283183 59322 283192
rect 59174 250064 59230 250073
rect 59174 249999 59230 250008
rect 59176 247036 59228 247042
rect 59176 246978 59228 246984
rect 59082 153232 59138 153241
rect 59082 153167 59138 153176
rect 58900 137284 58952 137290
rect 58900 137226 58952 137232
rect 59096 120018 59124 153167
rect 59084 120012 59136 120018
rect 59084 119954 59136 119960
rect 59188 101454 59216 246978
rect 60476 241369 60504 291790
rect 60568 271998 60596 429218
rect 60660 398818 60688 558894
rect 61842 519480 61898 519489
rect 61842 519415 61898 519424
rect 61752 434036 61804 434042
rect 61752 433978 61804 433984
rect 61660 418260 61712 418266
rect 61660 418202 61712 418208
rect 60648 398812 60700 398818
rect 60648 398754 60700 398760
rect 60648 314696 60700 314702
rect 60648 314638 60700 314644
rect 60660 279478 60688 314638
rect 60648 279472 60700 279478
rect 60648 279414 60700 279420
rect 60648 273284 60700 273290
rect 60648 273226 60700 273232
rect 60556 271992 60608 271998
rect 60556 271934 60608 271940
rect 60556 263900 60608 263906
rect 60556 263842 60608 263848
rect 60462 241360 60518 241369
rect 60462 241295 60518 241304
rect 60568 162994 60596 263842
rect 60556 162988 60608 162994
rect 60556 162930 60608 162936
rect 60464 155916 60516 155922
rect 60464 155858 60516 155864
rect 60476 154698 60504 155858
rect 60464 154692 60516 154698
rect 60464 154634 60516 154640
rect 59268 143608 59320 143614
rect 59268 143550 59320 143556
rect 59280 124982 59308 143550
rect 59268 124976 59320 124982
rect 59268 124918 59320 124924
rect 60476 124166 60504 154634
rect 60464 124160 60516 124166
rect 60464 124102 60516 124108
rect 60568 114510 60596 162930
rect 60660 155922 60688 273226
rect 60740 267708 60792 267714
rect 60740 267650 60792 267656
rect 60752 266529 60780 267650
rect 60738 266520 60794 266529
rect 60738 266455 60794 266464
rect 61672 263906 61700 418202
rect 61764 309806 61792 433978
rect 61856 393446 61884 519415
rect 61948 515438 61976 579702
rect 64788 572756 64840 572762
rect 64788 572698 64840 572704
rect 63408 564460 63460 564466
rect 63408 564402 63460 564408
rect 62028 557592 62080 557598
rect 62028 557534 62080 557540
rect 61936 515432 61988 515438
rect 61936 515374 61988 515380
rect 61936 460964 61988 460970
rect 61936 460906 61988 460912
rect 61948 418130 61976 460906
rect 62040 460222 62068 557534
rect 63316 554804 63368 554810
rect 63316 554746 63368 554752
rect 63328 522986 63356 554746
rect 63316 522980 63368 522986
rect 63316 522922 63368 522928
rect 62028 460216 62080 460222
rect 62028 460158 62080 460164
rect 63224 448588 63276 448594
rect 63224 448530 63276 448536
rect 63130 439512 63186 439521
rect 63130 439447 63186 439456
rect 63144 425105 63172 439447
rect 63130 425096 63186 425105
rect 63130 425031 63186 425040
rect 63236 418266 63264 448530
rect 63316 430636 63368 430642
rect 63316 430578 63368 430584
rect 63224 418260 63276 418266
rect 63224 418202 63276 418208
rect 61936 418124 61988 418130
rect 61936 418066 61988 418072
rect 61936 411324 61988 411330
rect 61936 411266 61988 411272
rect 61844 393440 61896 393446
rect 61844 393382 61896 393388
rect 61752 309800 61804 309806
rect 61752 309742 61804 309748
rect 61764 306374 61792 309742
rect 61764 306346 61884 306374
rect 61856 276010 61884 306346
rect 61948 282169 61976 411266
rect 63224 404388 63276 404394
rect 63224 404330 63276 404336
rect 61934 282160 61990 282169
rect 61934 282095 61990 282104
rect 61844 276004 61896 276010
rect 61844 275946 61896 275952
rect 61752 271992 61804 271998
rect 61752 271934 61804 271940
rect 61660 263900 61712 263906
rect 61660 263842 61712 263848
rect 61764 159361 61792 271934
rect 61948 259418 61976 282095
rect 62028 266416 62080 266422
rect 62028 266358 62080 266364
rect 61936 259412 61988 259418
rect 61936 259354 61988 259360
rect 61844 193860 61896 193866
rect 61844 193802 61896 193808
rect 61750 159352 61806 159361
rect 61750 159287 61806 159296
rect 61764 158817 61792 159287
rect 61750 158808 61806 158817
rect 61750 158743 61806 158752
rect 60648 155916 60700 155922
rect 60648 155858 60700 155864
rect 60648 142860 60700 142866
rect 60648 142802 60700 142808
rect 60556 114504 60608 114510
rect 60556 114446 60608 114452
rect 59268 111104 59320 111110
rect 59268 111046 59320 111052
rect 59176 101448 59228 101454
rect 59176 101390 59228 101396
rect 57888 93832 57940 93838
rect 57888 93774 57940 93780
rect 56414 90944 56470 90953
rect 56414 90879 56470 90888
rect 56598 80744 56654 80753
rect 56598 80679 56654 80688
rect 54484 80028 54536 80034
rect 54484 79970 54536 79976
rect 55128 80028 55180 80034
rect 55128 79970 55180 79976
rect 54496 46238 54524 79970
rect 54484 46232 54536 46238
rect 54484 46174 54536 46180
rect 53838 44840 53894 44849
rect 53838 44775 53894 44784
rect 53104 33108 53156 33114
rect 53104 33050 53156 33056
rect 52552 22772 52604 22778
rect 52552 22714 52604 22720
rect 52564 16574 52592 22714
rect 53852 16574 53880 44775
rect 55218 28248 55274 28257
rect 55218 28183 55274 28192
rect 55232 16574 55260 28183
rect 56612 16574 56640 80679
rect 59280 70281 59308 111046
rect 60660 92410 60688 142802
rect 61752 128376 61804 128382
rect 61752 128318 61804 128324
rect 60648 92404 60700 92410
rect 60648 92346 60700 92352
rect 59266 70272 59322 70281
rect 59266 70207 59322 70216
rect 60740 33788 60792 33794
rect 60740 33730 60792 33736
rect 59360 29640 59412 29646
rect 59360 29582 59412 29588
rect 59372 16574 59400 29582
rect 60752 16574 60780 33730
rect 61764 32434 61792 128318
rect 61856 91050 61884 193802
rect 61934 158808 61990 158817
rect 61934 158743 61990 158752
rect 61948 121378 61976 158743
rect 62040 151910 62068 266358
rect 63236 253910 63264 404330
rect 63328 273290 63356 430578
rect 63420 391513 63448 564402
rect 64696 560380 64748 560386
rect 64696 560322 64748 560328
rect 64708 529145 64736 560322
rect 64694 529136 64750 529145
rect 64694 529071 64750 529080
rect 64696 440904 64748 440910
rect 64696 440846 64748 440852
rect 64708 426494 64736 440846
rect 64696 426488 64748 426494
rect 64696 426430 64748 426436
rect 64604 421116 64656 421122
rect 64604 421058 64656 421064
rect 63406 391504 63462 391513
rect 63406 391439 63462 391448
rect 63316 273284 63368 273290
rect 63316 273226 63368 273232
rect 63314 272096 63370 272105
rect 63314 272031 63370 272040
rect 63224 253904 63276 253910
rect 63224 253846 63276 253852
rect 63222 179480 63278 179489
rect 63222 179415 63278 179424
rect 62028 151904 62080 151910
rect 62028 151846 62080 151852
rect 61936 121372 61988 121378
rect 61936 121314 61988 121320
rect 62040 117298 62068 151846
rect 63132 142180 63184 142186
rect 63132 142122 63184 142128
rect 63144 131102 63172 142122
rect 63132 131096 63184 131102
rect 63132 131038 63184 131044
rect 63236 124409 63264 179415
rect 63328 160721 63356 272031
rect 64616 266422 64644 421058
rect 64708 270638 64736 426430
rect 64800 406434 64828 572698
rect 65996 569945 66024 585142
rect 66180 576842 66208 611322
rect 67364 582412 67416 582418
rect 67364 582354 67416 582360
rect 66902 580000 66958 580009
rect 66902 579935 66958 579944
rect 66916 579766 66944 579935
rect 66904 579760 66956 579766
rect 66904 579702 66956 579708
rect 66168 576836 66220 576842
rect 66168 576778 66220 576784
rect 66180 575929 66208 576778
rect 66166 575920 66222 575929
rect 66166 575855 66222 575864
rect 67376 575113 67404 582354
rect 67454 581088 67510 581097
rect 67454 581023 67510 581032
rect 67362 575104 67418 575113
rect 67362 575039 67418 575048
rect 67376 574122 67404 575039
rect 66076 574116 66128 574122
rect 66076 574058 66128 574064
rect 67364 574116 67416 574122
rect 67364 574058 67416 574064
rect 65982 569936 66038 569945
rect 65982 569871 66038 569880
rect 65890 563408 65946 563417
rect 65890 563343 65946 563352
rect 65904 535401 65932 563343
rect 65982 548312 66038 548321
rect 65982 548247 66038 548256
rect 65890 535392 65946 535401
rect 65890 535327 65946 535336
rect 65996 517274 66024 548247
rect 66088 537538 66116 574058
rect 66810 573200 66866 573209
rect 66810 573135 66866 573144
rect 66824 572762 66852 573135
rect 66812 572756 66864 572762
rect 66812 572698 66864 572704
rect 67468 572665 67496 581023
rect 67546 577280 67602 577289
rect 67546 577215 67602 577224
rect 67454 572656 67510 572665
rect 67454 572591 67510 572600
rect 67454 570208 67510 570217
rect 67454 570143 67510 570152
rect 66902 567488 66958 567497
rect 66902 567423 66958 567432
rect 66916 567254 66944 567423
rect 66904 567248 66956 567254
rect 66904 567190 66956 567196
rect 66442 564904 66498 564913
rect 66442 564839 66498 564848
rect 66456 564466 66484 564839
rect 66444 564460 66496 564466
rect 66444 564402 66496 564408
rect 66810 560688 66866 560697
rect 66810 560623 66866 560632
rect 66824 560386 66852 560623
rect 66812 560380 66864 560386
rect 66812 560322 66864 560328
rect 66810 559328 66866 559337
rect 66810 559263 66866 559272
rect 66824 558958 66852 559263
rect 66812 558952 66864 558958
rect 66812 558894 66864 558900
rect 66810 557968 66866 557977
rect 66810 557903 66866 557912
rect 66824 557598 66852 557903
rect 66812 557592 66864 557598
rect 66812 557534 66864 557540
rect 66534 555248 66590 555257
rect 66534 555183 66590 555192
rect 66548 554810 66576 555183
rect 66536 554804 66588 554810
rect 66536 554746 66588 554752
rect 66902 553616 66958 553625
rect 66902 553551 66958 553560
rect 66916 553450 66944 553551
rect 66904 553444 66956 553450
rect 66904 553386 66956 553392
rect 66166 546816 66222 546825
rect 66166 546751 66222 546760
rect 66076 537532 66128 537538
rect 66076 537474 66128 537480
rect 65984 517268 66036 517274
rect 65984 517210 66036 517216
rect 66180 462913 66208 546751
rect 67362 545456 67418 545465
rect 67362 545391 67418 545400
rect 66810 544096 66866 544105
rect 66810 544031 66866 544040
rect 66824 543794 66852 544031
rect 66812 543788 66864 543794
rect 66812 543730 66864 543736
rect 66260 543720 66312 543726
rect 66260 543662 66312 543668
rect 66272 543425 66300 543662
rect 66258 543416 66314 543425
rect 66258 543351 66314 543360
rect 66258 541376 66314 541385
rect 66258 541311 66314 541320
rect 66272 541006 66300 541311
rect 66260 541000 66312 541006
rect 66260 540942 66312 540948
rect 66258 540016 66314 540025
rect 66258 539951 66314 539960
rect 66272 539646 66300 539951
rect 66260 539640 66312 539646
rect 66260 539582 66312 539588
rect 67376 538801 67404 545391
rect 67362 538792 67418 538801
rect 67362 538727 67418 538736
rect 66166 462904 66222 462913
rect 66166 462839 66222 462848
rect 66076 453076 66128 453082
rect 66076 453018 66128 453024
rect 66088 435305 66116 453018
rect 67468 451897 67496 570143
rect 67454 451888 67510 451897
rect 67454 451823 67510 451832
rect 66168 443012 66220 443018
rect 66168 442954 66220 442960
rect 66074 435296 66130 435305
rect 66074 435231 66130 435240
rect 65892 434852 65944 434858
rect 65892 434794 65944 434800
rect 65800 430704 65852 430710
rect 65800 430646 65852 430652
rect 65812 425746 65840 430646
rect 65800 425740 65852 425746
rect 65800 425682 65852 425688
rect 65904 414089 65932 434794
rect 65982 432576 66038 432585
rect 65982 432511 66038 432520
rect 65890 414080 65946 414089
rect 65890 414015 65946 414024
rect 64788 406428 64840 406434
rect 64788 406370 64840 406376
rect 65892 398812 65944 398818
rect 65892 398754 65944 398760
rect 65904 375358 65932 398754
rect 65996 397361 66024 432511
rect 66088 430710 66116 435231
rect 66076 430704 66128 430710
rect 66076 430646 66128 430652
rect 66180 430522 66208 442954
rect 67364 438932 67416 438938
rect 67364 438874 67416 438880
rect 67272 437504 67324 437510
rect 67272 437446 67324 437452
rect 66812 434036 66864 434042
rect 66812 433978 66864 433984
rect 66824 433401 66852 433978
rect 66810 433392 66866 433401
rect 66810 433327 66866 433336
rect 66088 430494 66208 430522
rect 66088 429282 66116 430494
rect 66166 430400 66222 430409
rect 66166 430335 66222 430344
rect 66076 429276 66128 429282
rect 66076 429218 66128 429224
rect 66074 403744 66130 403753
rect 66074 403679 66130 403688
rect 65982 397352 66038 397361
rect 65982 397287 66038 397296
rect 65996 393446 66024 393477
rect 65984 393440 66036 393446
rect 65982 393408 65984 393417
rect 66036 393408 66038 393417
rect 65982 393343 66038 393352
rect 65996 382974 66024 393343
rect 65984 382968 66036 382974
rect 65984 382910 66036 382916
rect 65982 376000 66038 376009
rect 65982 375935 66038 375944
rect 65892 375352 65944 375358
rect 65892 375294 65944 375300
rect 64788 289128 64840 289134
rect 64788 289070 64840 289076
rect 64696 270632 64748 270638
rect 64696 270574 64748 270580
rect 64604 266416 64656 266422
rect 64604 266358 64656 266364
rect 63408 264988 63460 264994
rect 63408 264930 63460 264936
rect 63314 160712 63370 160721
rect 63314 160647 63370 160656
rect 63222 124400 63278 124409
rect 63222 124335 63278 124344
rect 63328 122806 63356 160647
rect 63420 151094 63448 264930
rect 64604 256012 64656 256018
rect 64604 255954 64656 255960
rect 64616 222154 64644 255954
rect 64604 222148 64656 222154
rect 64604 222090 64656 222096
rect 63408 151088 63460 151094
rect 63408 151030 63460 151036
rect 63316 122800 63368 122806
rect 63316 122742 63368 122748
rect 62028 117292 62080 117298
rect 62028 117234 62080 117240
rect 63420 115598 63448 151030
rect 64510 138272 64566 138281
rect 64510 138207 64566 138216
rect 64524 126954 64552 138207
rect 64512 126948 64564 126954
rect 64512 126890 64564 126896
rect 63408 115592 63460 115598
rect 63408 115534 63460 115540
rect 63408 113824 63460 113830
rect 63408 113766 63460 113772
rect 61844 91044 61896 91050
rect 61844 90986 61896 90992
rect 63420 89690 63448 113766
rect 64616 107642 64644 222090
rect 64708 148374 64736 270574
rect 64800 251174 64828 289070
rect 65890 283248 65946 283257
rect 65890 283183 65946 283192
rect 65904 278322 65932 283183
rect 65892 278316 65944 278322
rect 65892 278258 65944 278264
rect 65890 276040 65946 276049
rect 65890 275975 65946 275984
rect 64880 251184 64932 251190
rect 64800 251146 64880 251174
rect 64880 251126 64932 251132
rect 64788 249076 64840 249082
rect 64788 249018 64840 249024
rect 64696 148368 64748 148374
rect 64696 148310 64748 148316
rect 64708 120086 64736 148310
rect 64696 120080 64748 120086
rect 64696 120022 64748 120028
rect 64604 107636 64656 107642
rect 64604 107578 64656 107584
rect 64696 100768 64748 100774
rect 64696 100710 64748 100716
rect 63408 89684 63460 89690
rect 63408 89626 63460 89632
rect 64708 85513 64736 100710
rect 64800 99686 64828 249018
rect 64892 247042 64920 251126
rect 64880 247036 64932 247042
rect 64880 246978 64932 246984
rect 65904 164354 65932 275975
rect 65996 238649 66024 375935
rect 66088 251870 66116 403679
rect 66180 272649 66208 430335
rect 66626 429312 66682 429321
rect 66626 429247 66628 429256
rect 66680 429247 66682 429256
rect 66628 429218 66680 429224
rect 66810 427408 66866 427417
rect 66810 427343 66866 427352
rect 66824 426494 66852 427343
rect 66812 426488 66864 426494
rect 66812 426430 66864 426436
rect 66628 425740 66680 425746
rect 66628 425682 66680 425688
rect 66640 425241 66668 425682
rect 66626 425232 66682 425241
rect 66626 425167 66682 425176
rect 66810 424144 66866 424153
rect 66810 424079 66866 424088
rect 66824 423706 66852 424079
rect 66812 423700 66864 423706
rect 66812 423642 66864 423648
rect 66258 423328 66314 423337
rect 66258 423263 66314 423272
rect 66272 422346 66300 423263
rect 66260 422340 66312 422346
rect 66260 422282 66312 422288
rect 67178 422240 67234 422249
rect 67178 422175 67234 422184
rect 66902 421152 66958 421161
rect 67192 421122 67220 422175
rect 66902 421087 66958 421096
rect 67180 421116 67232 421122
rect 66916 420986 66944 421087
rect 67180 421058 67232 421064
rect 66904 420980 66956 420986
rect 66904 420922 66956 420928
rect 66626 418976 66682 418985
rect 66626 418911 66682 418920
rect 66640 418266 66668 418911
rect 66628 418260 66680 418266
rect 66628 418202 66680 418208
rect 66994 418160 67050 418169
rect 66994 418095 66996 418104
rect 67048 418095 67050 418104
rect 66996 418066 67048 418072
rect 66812 416084 66864 416090
rect 66812 416026 66864 416032
rect 66824 415993 66852 416026
rect 66810 415984 66866 415993
rect 66810 415919 66866 415928
rect 66810 414896 66866 414905
rect 66810 414831 66866 414840
rect 66824 414050 66852 414831
rect 66812 414044 66864 414050
rect 66812 413986 66864 413992
rect 66628 413296 66680 413302
rect 66628 413238 66680 413244
rect 66640 413001 66668 413238
rect 66626 412992 66682 413001
rect 66626 412927 66682 412936
rect 67008 412634 67036 418066
rect 67008 412606 67220 412634
rect 66902 411904 66958 411913
rect 66902 411839 66958 411848
rect 66916 411330 66944 411839
rect 66904 411324 66956 411330
rect 66904 411266 66956 411272
rect 66812 411256 66864 411262
rect 66812 411198 66864 411204
rect 66824 410825 66852 411198
rect 66810 410816 66866 410825
rect 66810 410751 66866 410760
rect 66810 408912 66866 408921
rect 66810 408847 66866 408856
rect 66824 408542 66852 408847
rect 66812 408536 66864 408542
rect 66812 408478 66864 408484
rect 66904 408468 66956 408474
rect 66904 408410 66956 408416
rect 66916 407833 66944 408410
rect 66902 407824 66958 407833
rect 66902 407759 66958 407768
rect 66810 406736 66866 406745
rect 66810 406671 66866 406680
rect 66824 406434 66852 406671
rect 66812 406428 66864 406434
rect 66812 406370 66864 406376
rect 66810 404560 66866 404569
rect 66810 404495 66866 404504
rect 66824 404394 66852 404495
rect 66812 404388 66864 404394
rect 66812 404330 66864 404336
rect 66810 401568 66866 401577
rect 66810 401503 66866 401512
rect 66824 400246 66852 401503
rect 66812 400240 66864 400246
rect 66812 400182 66864 400188
rect 66810 399664 66866 399673
rect 66810 399599 66866 399608
rect 66824 398886 66852 399599
rect 66812 398880 66864 398886
rect 66812 398822 66864 398828
rect 66536 398812 66588 398818
rect 66536 398754 66588 398760
rect 66548 398585 66576 398754
rect 66534 398576 66590 398585
rect 66534 398511 66590 398520
rect 67088 397520 67140 397526
rect 67086 397488 67088 397497
rect 67140 397488 67142 397497
rect 67086 397423 67142 397432
rect 66810 392320 66866 392329
rect 66810 392255 66866 392264
rect 66824 392018 66852 392255
rect 66812 392012 66864 392018
rect 66812 391954 66864 391960
rect 67192 345014 67220 412606
rect 67284 405657 67312 437446
rect 67376 420073 67404 438874
rect 67362 420064 67418 420073
rect 67362 419999 67418 420008
rect 67468 417081 67496 451823
rect 67560 437510 67588 577215
rect 67652 566681 67680 702510
rect 71044 700324 71096 700330
rect 71044 700266 71096 700272
rect 69848 593428 69900 593434
rect 69848 593370 69900 593376
rect 69860 581074 69888 593370
rect 71056 582418 71084 700266
rect 72988 699825 73016 703520
rect 85580 702636 85632 702642
rect 85580 702578 85632 702584
rect 72974 699816 73030 699825
rect 72974 699751 73030 699760
rect 74540 656940 74592 656946
rect 74540 656882 74592 656888
rect 74552 596174 74580 656882
rect 81440 621036 81492 621042
rect 81440 620978 81492 620984
rect 75918 599312 75974 599321
rect 75918 599247 75974 599256
rect 75932 596174 75960 599247
rect 74552 596146 74672 596174
rect 75932 596146 76512 596174
rect 71780 591320 71832 591326
rect 71780 591262 71832 591268
rect 71044 582412 71096 582418
rect 71044 582354 71096 582360
rect 71792 581074 71820 591262
rect 74264 583772 74316 583778
rect 74264 583714 74316 583720
rect 73526 582584 73582 582593
rect 73526 582519 73582 582528
rect 73540 581074 73568 582519
rect 74276 581074 74304 583714
rect 69860 581046 70288 581074
rect 71792 581046 72128 581074
rect 73232 581046 73568 581074
rect 74152 581046 74304 581074
rect 74644 581074 74672 596146
rect 76288 581120 76340 581126
rect 74644 581046 75408 581074
rect 75992 581068 76288 581074
rect 75992 581062 76340 581068
rect 76484 581074 76512 596146
rect 78128 588668 78180 588674
rect 78128 588610 78180 588616
rect 78140 581074 78168 588610
rect 79968 583840 80020 583846
rect 79968 583782 80020 583788
rect 79980 581074 80008 583782
rect 80704 582412 80756 582418
rect 80704 582354 80756 582360
rect 75992 581046 76328 581062
rect 76484 581046 76912 581074
rect 77832 581046 78168 581074
rect 79672 581046 80008 581074
rect 75380 580961 75408 581046
rect 75366 580952 75422 580961
rect 75366 580887 75422 580896
rect 79980 580825 80008 581046
rect 80244 581052 80296 581058
rect 80244 580994 80296 581000
rect 80256 580938 80284 580994
rect 80716 580938 80744 582354
rect 81452 581346 81480 620978
rect 84108 597576 84160 597582
rect 84108 597518 84160 597524
rect 82726 582720 82782 582729
rect 84120 582690 84148 597518
rect 85592 596174 85620 702578
rect 89180 702434 89208 703520
rect 96620 702500 96672 702506
rect 96620 702442 96672 702448
rect 88352 702406 89208 702434
rect 86960 599616 87012 599622
rect 86960 599558 87012 599564
rect 85592 596146 85896 596174
rect 82726 582655 82782 582664
rect 84108 582684 84160 582690
rect 81452 581318 81526 581346
rect 81498 581060 81526 581318
rect 82740 581074 82768 582655
rect 84108 582626 84160 582632
rect 85028 582684 85080 582690
rect 85028 582626 85080 582632
rect 83004 582480 83056 582486
rect 83004 582422 83056 582428
rect 82432 581046 82768 581074
rect 83016 581074 83044 582422
rect 85040 581074 85068 582626
rect 85868 581074 85896 596146
rect 86972 581074 87000 599558
rect 88352 592090 88380 702406
rect 94688 605872 94740 605878
rect 94688 605814 94740 605820
rect 88982 603256 89038 603265
rect 88982 603191 89038 603200
rect 88260 592062 88380 592090
rect 88260 588674 88288 592062
rect 88248 588668 88300 588674
rect 88248 588610 88300 588616
rect 88996 583234 89024 603191
rect 94700 596174 94728 605814
rect 94700 596146 95004 596174
rect 92480 594856 92532 594862
rect 92480 594798 92532 594804
rect 89720 592680 89772 592686
rect 89720 592622 89772 592628
rect 88248 583228 88300 583234
rect 88248 583170 88300 583176
rect 88984 583228 89036 583234
rect 88984 583170 89036 583176
rect 88260 581074 88288 583170
rect 83016 581046 83352 581074
rect 85040 581046 85376 581074
rect 85868 581058 86632 581074
rect 85868 581052 86644 581058
rect 85868 581046 86592 581052
rect 86972 581046 87216 581074
rect 88136 581046 88288 581074
rect 89732 581074 89760 592622
rect 91376 589348 91428 589354
rect 91376 589290 91428 589296
rect 91008 582480 91060 582486
rect 91008 582422 91060 582428
rect 91020 581074 91048 582422
rect 89732 581046 89976 581074
rect 90896 581046 91048 581074
rect 91388 581074 91416 589290
rect 92492 581074 92520 594798
rect 94870 583400 94926 583409
rect 94870 583335 94926 583344
rect 93766 581224 93822 581233
rect 93766 581159 93822 581168
rect 93780 581074 93808 581159
rect 94884 581074 94912 583335
rect 91388 581046 91816 581074
rect 92492 581046 92736 581074
rect 93656 581046 93808 581074
rect 94576 581046 94912 581074
rect 86592 580994 86644 581000
rect 80256 580910 80744 580938
rect 70950 580816 71006 580825
rect 69032 580774 69368 580802
rect 69032 580718 69060 580774
rect 79966 580816 80022 580825
rect 71006 580774 71208 580802
rect 78752 580774 79088 580802
rect 70950 580751 71006 580760
rect 79060 580718 79088 580774
rect 84658 580816 84714 580825
rect 84456 580774 84658 580802
rect 79966 580751 80022 580760
rect 89258 580816 89314 580825
rect 89056 580774 89258 580802
rect 84658 580751 84714 580760
rect 89258 580751 89314 580760
rect 69020 580712 69072 580718
rect 69020 580654 69072 580660
rect 79048 580712 79100 580718
rect 79048 580654 79100 580660
rect 94976 579630 95004 596146
rect 95332 588600 95384 588606
rect 95332 588542 95384 588548
rect 94964 579624 95016 579630
rect 94964 579566 95016 579572
rect 67730 575920 67786 575929
rect 67730 575855 67786 575864
rect 67638 566672 67694 566681
rect 67638 566607 67694 566616
rect 67652 565894 67680 566607
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67638 556608 67694 556617
rect 67638 556543 67694 556552
rect 67652 538898 67680 556543
rect 67640 538892 67692 538898
rect 67640 538834 67692 538840
rect 67744 529281 67772 575855
rect 95238 563680 95294 563689
rect 95238 563615 95294 563624
rect 95148 558884 95200 558890
rect 95146 558852 95148 558861
rect 95200 558852 95202 558861
rect 95146 558787 95202 558796
rect 94686 558648 94742 558657
rect 94686 558583 94742 558592
rect 67822 552256 67878 552265
rect 67822 552191 67878 552200
rect 67836 539850 67864 552191
rect 67824 539844 67876 539850
rect 67824 539786 67876 539792
rect 71780 539844 71832 539850
rect 71780 539786 71832 539792
rect 68816 539158 68968 539186
rect 68940 535537 68968 539158
rect 69400 539158 69736 539186
rect 70656 539158 70716 539186
rect 69400 536110 69428 539158
rect 69662 539064 69718 539073
rect 69662 538999 69718 539008
rect 69676 536217 69704 538999
rect 70688 538218 70716 539158
rect 70964 539158 71576 539186
rect 70676 538212 70728 538218
rect 70676 538154 70728 538160
rect 70688 536858 70716 538154
rect 70676 536852 70728 536858
rect 70676 536794 70728 536800
rect 69662 536208 69718 536217
rect 69662 536143 69718 536152
rect 69388 536104 69440 536110
rect 69388 536046 69440 536052
rect 68926 535528 68982 535537
rect 68926 535463 68982 535472
rect 67730 529272 67786 529281
rect 67730 529207 67786 529216
rect 70964 528554 70992 539158
rect 71044 536852 71096 536858
rect 71044 536794 71096 536800
rect 70504 528526 70992 528554
rect 69664 517268 69716 517274
rect 69664 517210 69716 517216
rect 68926 467936 68982 467945
rect 68926 467871 68982 467880
rect 68284 458856 68336 458862
rect 68284 458798 68336 458804
rect 67640 445732 67692 445738
rect 67640 445674 67692 445680
rect 67548 437504 67600 437510
rect 67548 437446 67600 437452
rect 67548 434716 67600 434722
rect 67548 434658 67600 434664
rect 67560 431497 67588 434658
rect 67546 431488 67602 431497
rect 67546 431423 67602 431432
rect 67560 430642 67588 431423
rect 67548 430636 67600 430642
rect 67548 430578 67600 430584
rect 67454 417072 67510 417081
rect 67454 417007 67510 417016
rect 67652 409737 67680 445674
rect 67732 441652 67784 441658
rect 67732 441594 67784 441600
rect 68296 441614 68324 458798
rect 68940 450634 68968 467871
rect 68928 450628 68980 450634
rect 68928 450570 68980 450576
rect 67744 428233 67772 441594
rect 68296 441586 68416 441614
rect 68388 434761 68416 441586
rect 69676 438841 69704 517210
rect 70308 456816 70360 456822
rect 70308 456758 70360 456764
rect 70320 441614 70348 456758
rect 70504 453082 70532 528526
rect 71056 523734 71084 536794
rect 71044 523728 71096 523734
rect 71044 523670 71096 523676
rect 70492 453076 70544 453082
rect 70492 453018 70544 453024
rect 70872 448662 70900 448693
rect 70860 448656 70912 448662
rect 70858 448624 70860 448633
rect 70912 448624 70914 448633
rect 70858 448559 70914 448568
rect 70872 445738 70900 448559
rect 71136 446412 71188 446418
rect 71136 446354 71188 446360
rect 70860 445732 70912 445738
rect 70860 445674 70912 445680
rect 70400 444440 70452 444446
rect 70400 444382 70452 444388
rect 69952 441586 70348 441614
rect 70412 441614 70440 444382
rect 71148 441614 71176 446354
rect 70412 441586 71084 441614
rect 71148 441586 71360 441614
rect 69662 438832 69718 438841
rect 69662 438767 69718 438776
rect 69676 436218 69704 438767
rect 69664 436212 69716 436218
rect 69664 436154 69716 436160
rect 68374 434752 68430 434761
rect 68374 434687 68430 434696
rect 68388 434330 68416 434687
rect 69294 434344 69350 434353
rect 68388 434302 68816 434330
rect 69952 434330 69980 441586
rect 71056 437474 71084 441586
rect 71056 437446 71176 437474
rect 70032 436212 70084 436218
rect 70032 436154 70084 436160
rect 69350 434302 69980 434330
rect 70044 434330 70072 436154
rect 70860 436144 70912 436150
rect 70860 436086 70912 436092
rect 70044 434302 70288 434330
rect 69294 434279 69350 434288
rect 68652 434104 68704 434110
rect 68652 434046 68704 434052
rect 70872 434058 70900 436086
rect 71148 434330 71176 437446
rect 71332 434722 71360 441586
rect 71320 434716 71372 434722
rect 71320 434658 71372 434664
rect 71148 434302 71576 434330
rect 71792 434110 71820 539786
rect 94136 539708 94188 539714
rect 94136 539650 94188 539656
rect 88156 539640 88208 539646
rect 73066 539608 73122 539617
rect 76746 539608 76802 539617
rect 73122 539566 73200 539594
rect 73066 539543 73122 539552
rect 71884 539158 72496 539186
rect 71884 525094 71912 539158
rect 72422 535528 72478 535537
rect 72422 535463 72478 535472
rect 71872 525088 71924 525094
rect 71872 525030 71924 525036
rect 72436 518226 72464 535463
rect 73172 533390 73200 539566
rect 76802 539566 77096 539594
rect 88156 539582 88208 539588
rect 76746 539543 76802 539552
rect 73416 539158 73476 539186
rect 73448 538214 73476 539158
rect 73264 538186 73476 538214
rect 73632 539158 74336 539186
rect 74552 539158 75256 539186
rect 76024 539158 76176 539186
rect 77312 539158 78016 539186
rect 78936 539158 79272 539186
rect 80040 539158 80100 539186
rect 73264 536790 73292 538186
rect 73252 536784 73304 536790
rect 73252 536726 73304 536732
rect 73264 536110 73292 536726
rect 73252 536104 73304 536110
rect 73252 536046 73304 536052
rect 73160 533384 73212 533390
rect 73160 533326 73212 533332
rect 73632 528554 73660 539158
rect 73172 528526 73660 528554
rect 72424 518220 72476 518226
rect 72424 518162 72476 518168
rect 73172 454753 73200 528526
rect 74552 460970 74580 539158
rect 75828 533384 75880 533390
rect 75828 533326 75880 533332
rect 75734 461000 75790 461009
rect 74540 460964 74592 460970
rect 75734 460935 75790 460944
rect 74540 460906 74592 460912
rect 74552 460193 74580 460906
rect 74538 460184 74594 460193
rect 74538 460119 74594 460128
rect 75184 455388 75236 455394
rect 75184 455330 75236 455336
rect 73158 454744 73214 454753
rect 73158 454679 73214 454688
rect 74446 452976 74502 452985
rect 74446 452911 74502 452920
rect 73160 447840 73212 447846
rect 73160 447782 73212 447788
rect 73172 441614 73200 447782
rect 73172 441586 73384 441614
rect 73356 434330 73384 441586
rect 73356 434302 73784 434330
rect 71780 434104 71832 434110
rect 67730 428224 67786 428233
rect 67730 428159 67786 428168
rect 67638 409728 67694 409737
rect 67638 409663 67694 409672
rect 67270 405648 67326 405657
rect 67270 405583 67326 405592
rect 67640 403640 67692 403646
rect 67640 403582 67692 403588
rect 67362 400480 67418 400489
rect 67362 400415 67418 400424
rect 67284 395350 67312 395381
rect 67272 395344 67324 395350
rect 67270 395312 67272 395321
rect 67324 395312 67326 395321
rect 67270 395247 67326 395256
rect 67284 386345 67312 395247
rect 67376 388482 67404 400415
rect 67652 398834 67680 403582
rect 67822 402656 67878 402665
rect 67822 402591 67878 402600
rect 67560 398806 67680 398834
rect 67454 397488 67510 397497
rect 67454 397423 67510 397432
rect 67364 388476 67416 388482
rect 67364 388418 67416 388424
rect 67270 386336 67326 386345
rect 67270 386271 67326 386280
rect 67468 383625 67496 397423
rect 67560 396409 67588 398806
rect 67546 396400 67602 396409
rect 67546 396335 67602 396344
rect 67730 394496 67786 394505
rect 67730 394431 67786 394440
rect 67640 390176 67692 390182
rect 67640 390118 67692 390124
rect 67454 383616 67510 383625
rect 67454 383551 67510 383560
rect 67652 357377 67680 390118
rect 67744 367062 67772 394431
rect 67836 378049 67864 402591
rect 68560 391332 68612 391338
rect 68560 391274 68612 391280
rect 68572 391134 68600 391274
rect 68560 391128 68612 391134
rect 68560 391070 68612 391076
rect 67822 378040 67878 378049
rect 67822 377975 67878 377984
rect 67732 367056 67784 367062
rect 67732 366998 67784 367004
rect 67638 357368 67694 357377
rect 67638 357303 67694 357312
rect 67192 344986 67496 345014
rect 67468 340950 67496 344986
rect 67456 340944 67508 340950
rect 67456 340886 67508 340892
rect 67364 305652 67416 305658
rect 67364 305594 67416 305600
rect 66260 283620 66312 283626
rect 66260 283562 66312 283568
rect 66272 282985 66300 283562
rect 66258 282976 66314 282985
rect 66258 282911 66314 282920
rect 66720 280220 66772 280226
rect 66720 280162 66772 280168
rect 66732 277394 66760 280162
rect 66812 279472 66864 279478
rect 66812 279414 66864 279420
rect 66824 278905 66852 279414
rect 66810 278896 66866 278905
rect 66810 278831 66866 278840
rect 66732 277366 66852 277394
rect 66166 272640 66222 272649
rect 66166 272575 66222 272584
rect 66720 269068 66772 269074
rect 66720 269010 66772 269016
rect 66732 268297 66760 269010
rect 66718 268288 66774 268297
rect 66718 268223 66774 268232
rect 66258 265024 66314 265033
rect 66258 264959 66260 264968
rect 66312 264959 66314 264968
rect 66260 264930 66312 264936
rect 66258 264208 66314 264217
rect 66258 264143 66314 264152
rect 66272 263906 66300 264143
rect 66260 263900 66312 263906
rect 66260 263842 66312 263848
rect 66258 263392 66314 263401
rect 66180 263350 66258 263378
rect 66180 261526 66208 263350
rect 66258 263327 66314 263336
rect 66350 262848 66406 262857
rect 66350 262783 66406 262792
rect 66258 262576 66314 262585
rect 66258 262511 66314 262520
rect 66272 262274 66300 262511
rect 66260 262268 66312 262274
rect 66260 262210 66312 262216
rect 66258 261760 66314 261769
rect 66258 261695 66314 261704
rect 66272 261594 66300 261695
rect 66260 261588 66312 261594
rect 66260 261530 66312 261536
rect 66168 261520 66220 261526
rect 66168 261462 66220 261468
rect 66272 260166 66300 261530
rect 66364 260953 66392 262783
rect 66350 260944 66406 260953
rect 66350 260879 66406 260888
rect 66260 260160 66312 260166
rect 66260 260102 66312 260108
rect 66628 259412 66680 259418
rect 66628 259354 66680 259360
rect 66352 258732 66404 258738
rect 66352 258674 66404 258680
rect 66364 258058 66392 258674
rect 66640 258505 66668 259354
rect 66626 258496 66682 258505
rect 66626 258431 66682 258440
rect 66352 258052 66404 258058
rect 66352 257994 66404 258000
rect 66258 257680 66314 257689
rect 66258 257615 66314 257624
rect 66272 256766 66300 257615
rect 66260 256760 66312 256766
rect 66260 256702 66312 256708
rect 66718 255232 66774 255241
rect 66718 255167 66774 255176
rect 66732 254590 66760 255167
rect 66720 254584 66772 254590
rect 66720 254526 66772 254532
rect 66628 253904 66680 253910
rect 66628 253846 66680 253852
rect 66640 252793 66668 253846
rect 66166 252784 66222 252793
rect 66166 252719 66222 252728
rect 66626 252784 66682 252793
rect 66626 252719 66682 252728
rect 66076 251864 66128 251870
rect 66076 251806 66128 251812
rect 65982 238640 66038 238649
rect 65982 238575 66038 238584
rect 65892 164348 65944 164354
rect 65892 164290 65944 164296
rect 65904 161474 65932 164290
rect 65904 161446 66116 161474
rect 65984 153876 66036 153882
rect 65984 153818 66036 153824
rect 65892 138032 65944 138038
rect 65892 137974 65944 137980
rect 65904 103193 65932 137974
rect 65996 133657 66024 153818
rect 65982 133648 66038 133657
rect 65982 133583 66038 133592
rect 66088 126041 66116 161446
rect 66180 138718 66208 252719
rect 66626 251968 66682 251977
rect 66626 251903 66682 251912
rect 66640 251870 66668 251903
rect 66628 251864 66680 251870
rect 66628 251806 66680 251812
rect 66260 251184 66312 251190
rect 66258 251152 66260 251161
rect 66312 251152 66314 251161
rect 66258 251087 66314 251096
rect 66626 247888 66682 247897
rect 66626 247823 66682 247832
rect 66640 247110 66668 247823
rect 66628 247104 66680 247110
rect 66628 247046 66680 247052
rect 66534 243808 66590 243817
rect 66534 243743 66590 243752
rect 66548 242962 66576 243743
rect 66536 242956 66588 242962
rect 66536 242898 66588 242904
rect 66168 138712 66220 138718
rect 66168 138654 66220 138660
rect 66180 138038 66208 138654
rect 66168 138032 66220 138038
rect 66168 137974 66220 137980
rect 66824 132494 66852 277366
rect 66904 277364 66956 277370
rect 66904 277306 66956 277312
rect 66916 276457 66944 277306
rect 66902 276448 66958 276457
rect 66902 276383 66958 276392
rect 66904 276004 66956 276010
rect 66904 275946 66956 275952
rect 66916 275641 66944 275946
rect 66902 275632 66958 275641
rect 66902 275567 66958 275576
rect 66902 274000 66958 274009
rect 66902 273935 66958 273944
rect 66916 273290 66944 273935
rect 66904 273284 66956 273290
rect 66904 273226 66956 273232
rect 67272 273284 67324 273290
rect 67272 273226 67324 273232
rect 66902 272368 66958 272377
rect 66902 272303 66958 272312
rect 66916 271998 66944 272303
rect 66904 271992 66956 271998
rect 66904 271934 66956 271940
rect 66902 270736 66958 270745
rect 66902 270671 66958 270680
rect 66916 270638 66944 270671
rect 66904 270632 66956 270638
rect 66904 270574 66956 270580
rect 66902 269920 66958 269929
rect 66902 269855 66958 269864
rect 66916 269822 66944 269855
rect 66904 269816 66956 269822
rect 66904 269758 66956 269764
rect 66902 266656 66958 266665
rect 66902 266591 66958 266600
rect 66916 266422 66944 266591
rect 66904 266416 66956 266422
rect 66904 266358 66956 266364
rect 67284 260137 67312 273226
rect 66994 260128 67050 260137
rect 66994 260063 67050 260072
rect 67270 260128 67326 260137
rect 67270 260063 67326 260072
rect 66902 256048 66958 256057
rect 66902 255983 66904 255992
rect 66956 255983 66958 255992
rect 66904 255954 66956 255960
rect 66904 254720 66956 254726
rect 66904 254662 66956 254668
rect 66916 254425 66944 254662
rect 66902 254416 66958 254425
rect 66902 254351 66958 254360
rect 66902 253600 66958 253609
rect 66902 253535 66958 253544
rect 66916 253230 66944 253535
rect 66904 253224 66956 253230
rect 66904 253166 66956 253172
rect 67008 250510 67036 260063
rect 67376 256873 67404 305594
rect 67468 263401 67496 340886
rect 68664 306374 68692 434046
rect 70872 434030 71024 434058
rect 72700 434104 72752 434110
rect 71780 434046 71832 434052
rect 72312 434042 72648 434058
rect 72752 434052 73048 434058
rect 72700 434046 73048 434052
rect 72312 434036 72660 434042
rect 72312 434030 72608 434036
rect 72712 434030 73048 434046
rect 72608 433978 72660 433984
rect 73988 433696 74040 433702
rect 74460 433650 74488 452911
rect 75196 436150 75224 455330
rect 75748 441614 75776 460935
rect 75840 455394 75868 533326
rect 76024 502314 76052 539158
rect 76012 502308 76064 502314
rect 76012 502250 76064 502256
rect 77208 502308 77260 502314
rect 77208 502250 77260 502256
rect 77220 501634 77248 502250
rect 77208 501628 77260 501634
rect 77208 501570 77260 501576
rect 75828 455388 75880 455394
rect 75828 455330 75880 455336
rect 77116 445052 77168 445058
rect 77116 444994 77168 445000
rect 77128 441614 77156 444994
rect 77220 442950 77248 501570
rect 77312 450566 77340 539158
rect 79244 537742 79272 539158
rect 80072 538393 80100 539158
rect 80164 539158 80960 539186
rect 81880 539158 82216 539186
rect 82800 539158 83136 539186
rect 83720 539158 84056 539186
rect 80058 538384 80114 538393
rect 80058 538319 80114 538328
rect 79968 538212 80020 538218
rect 79968 538154 80020 538160
rect 79980 537742 80008 538154
rect 79232 537736 79284 537742
rect 79232 537678 79284 537684
rect 79968 537736 80020 537742
rect 79968 537678 80020 537684
rect 79980 472666 80008 537678
rect 80164 528554 80192 539158
rect 81990 538792 82046 538801
rect 81990 538727 82046 538736
rect 81440 536104 81492 536110
rect 81440 536046 81492 536052
rect 81452 533458 81480 536046
rect 81440 533452 81492 533458
rect 81440 533394 81492 533400
rect 82004 530602 82032 538727
rect 82188 536722 82216 539158
rect 82176 536716 82228 536722
rect 82176 536658 82228 536664
rect 82728 534744 82780 534750
rect 82728 534686 82780 534692
rect 81992 530596 82044 530602
rect 81992 530538 82044 530544
rect 80072 528526 80192 528554
rect 79968 472660 80020 472666
rect 79968 472602 80020 472608
rect 79324 471300 79376 471306
rect 79324 471242 79376 471248
rect 77668 452668 77720 452674
rect 77668 452610 77720 452616
rect 77300 450560 77352 450566
rect 77300 450502 77352 450508
rect 77680 447846 77708 452610
rect 77668 447840 77720 447846
rect 77668 447782 77720 447788
rect 78680 443080 78732 443086
rect 78680 443022 78732 443028
rect 77208 442944 77260 442950
rect 77208 442886 77260 442892
rect 75380 441586 75776 441614
rect 76944 441586 77156 441614
rect 78692 441614 78720 443022
rect 78692 441586 78904 441614
rect 75184 436144 75236 436150
rect 75184 436086 75236 436092
rect 74040 433644 74488 433650
rect 73988 433638 74488 433644
rect 74000 433622 74488 433638
rect 74814 433664 74870 433673
rect 75380 433650 75408 441586
rect 75458 436112 75514 436121
rect 75458 436047 75514 436056
rect 75472 434330 75500 436047
rect 75472 434302 75808 434330
rect 74870 433622 75408 433650
rect 76194 433664 76250 433673
rect 74814 433599 74870 433608
rect 76944 433650 76972 441586
rect 78588 440292 78640 440298
rect 78588 440234 78640 440240
rect 78220 436416 78272 436422
rect 78220 436358 78272 436364
rect 78232 433809 78260 436358
rect 78600 434602 78628 440234
rect 78554 434574 78628 434602
rect 78554 434316 78582 434574
rect 78876 434330 78904 441586
rect 79336 436422 79364 471242
rect 80072 457473 80100 528526
rect 80058 457464 80114 457473
rect 80058 457399 80114 457408
rect 82740 455462 82768 534686
rect 83108 532098 83136 539158
rect 83464 538892 83516 538898
rect 83464 538834 83516 538840
rect 83096 532092 83148 532098
rect 83096 532034 83148 532040
rect 82728 455456 82780 455462
rect 82728 455398 82780 455404
rect 82740 451274 82768 455398
rect 82648 451246 82768 451274
rect 80060 450628 80112 450634
rect 80060 450570 80112 450576
rect 79324 436416 79376 436422
rect 79324 436358 79376 436364
rect 80072 436257 80100 450570
rect 82648 441614 82676 451246
rect 83476 444514 83504 538834
rect 84028 538121 84056 539158
rect 84304 539158 84640 539186
rect 85560 539158 85620 539186
rect 84014 538112 84070 538121
rect 84014 538047 84070 538056
rect 84304 533361 84332 539158
rect 85592 538286 85620 539158
rect 85684 539158 86480 539186
rect 87400 539158 87736 539186
rect 85580 538280 85632 538286
rect 85580 538222 85632 538228
rect 84290 533352 84346 533361
rect 84290 533287 84346 533296
rect 85684 528554 85712 539158
rect 85764 538280 85816 538286
rect 85764 538222 85816 538228
rect 85776 530641 85804 538222
rect 87708 536790 87736 539158
rect 87696 536784 87748 536790
rect 87696 536726 87748 536732
rect 88168 536722 88196 539582
rect 88320 539158 88380 539186
rect 88156 536716 88208 536722
rect 88156 536658 88208 536664
rect 88352 535537 88380 539158
rect 88536 539158 89240 539186
rect 89824 539158 90160 539186
rect 91204 539158 91264 539186
rect 91848 539158 92184 539186
rect 93104 539158 93440 539186
rect 94024 539158 94084 539186
rect 88338 535528 88394 535537
rect 86224 535492 86276 535498
rect 88338 535463 88394 535472
rect 86224 535434 86276 535440
rect 85762 530632 85818 530641
rect 85762 530567 85818 530576
rect 85592 528526 85712 528554
rect 85488 476808 85540 476814
rect 85488 476750 85540 476756
rect 83464 444508 83516 444514
rect 83464 444450 83516 444456
rect 83188 442944 83240 442950
rect 83188 442886 83240 442892
rect 82464 441586 82676 441614
rect 80334 436520 80390 436529
rect 80334 436455 80390 436464
rect 80058 436248 80114 436257
rect 80058 436183 80114 436192
rect 80072 434602 80100 436183
rect 80026 434574 80100 434602
rect 78876 434302 79304 434330
rect 80026 434316 80054 434574
rect 80348 434330 80376 436455
rect 81164 436212 81216 436218
rect 81164 436154 81216 436160
rect 80348 434302 80592 434330
rect 80978 434072 81034 434081
rect 81176 434058 81204 436154
rect 81034 434030 81328 434058
rect 80978 434007 81034 434016
rect 77482 433800 77538 433809
rect 77280 433758 77482 433786
rect 77482 433735 77538 433744
rect 78218 433800 78274 433809
rect 78218 433735 78274 433744
rect 78126 433664 78182 433673
rect 76250 433622 76972 433650
rect 77832 433622 78126 433650
rect 76194 433599 76250 433608
rect 78126 433599 78182 433608
rect 81898 433664 81954 433673
rect 82464 433650 82492 441586
rect 82910 433664 82966 433673
rect 81954 433622 82492 433650
rect 82800 433622 82910 433650
rect 81898 433599 81954 433608
rect 83200 433650 83228 442886
rect 83476 434602 83504 444450
rect 85500 441614 85528 476750
rect 85592 460902 85620 528526
rect 85580 460896 85632 460902
rect 85580 460838 85632 460844
rect 85672 460216 85724 460222
rect 85672 460158 85724 460164
rect 85224 441586 85528 441614
rect 85684 441614 85712 460158
rect 86236 445058 86264 535434
rect 88248 535424 88300 535430
rect 88248 535366 88300 535372
rect 86224 445052 86276 445058
rect 86224 444994 86276 445000
rect 86868 445052 86920 445058
rect 86868 444994 86920 445000
rect 86880 444514 86908 444994
rect 86868 444508 86920 444514
rect 86868 444450 86920 444456
rect 88260 441726 88288 535366
rect 88536 528554 88564 539158
rect 89824 535498 89852 539158
rect 89812 535492 89864 535498
rect 89812 535434 89864 535440
rect 91008 535492 91060 535498
rect 91008 535434 91060 535440
rect 88352 528526 88564 528554
rect 88352 527134 88380 528526
rect 88340 527128 88392 527134
rect 88340 527070 88392 527076
rect 88982 482896 89038 482905
rect 88982 482831 89038 482840
rect 88996 481681 89024 482831
rect 88982 481672 89038 481681
rect 88982 481607 89038 481616
rect 88248 441720 88300 441726
rect 88248 441662 88300 441668
rect 85684 441586 85896 441614
rect 83738 440872 83794 440881
rect 83738 440807 83794 440816
rect 83476 434574 83550 434602
rect 83522 434316 83550 434574
rect 82966 433622 83228 433650
rect 83752 433650 83780 440807
rect 83830 433664 83886 433673
rect 83752 433622 83830 433650
rect 82910 433599 82966 433608
rect 84566 433664 84622 433673
rect 83886 433622 84088 433650
rect 83830 433599 83886 433608
rect 85224 433650 85252 441586
rect 85868 437474 85896 441586
rect 85868 437446 85988 437474
rect 85854 433800 85910 433809
rect 85560 433758 85854 433786
rect 85854 433735 85910 433744
rect 85960 433673 85988 437446
rect 88260 436150 88288 441662
rect 88430 436384 88486 436393
rect 88430 436319 88486 436328
rect 87328 436144 87380 436150
rect 87328 436086 87380 436092
rect 88248 436144 88300 436150
rect 88248 436086 88300 436092
rect 87340 434330 87368 436086
rect 87032 434302 87368 434330
rect 88444 434194 88472 436319
rect 88996 436218 89024 481607
rect 91020 469266 91048 535434
rect 91204 471306 91232 539158
rect 91848 535498 91876 539158
rect 93412 536761 93440 539158
rect 93398 536752 93454 536761
rect 93398 536687 93454 536696
rect 91836 535492 91888 535498
rect 91836 535434 91888 535440
rect 94056 531350 94084 539158
rect 93124 531344 93176 531350
rect 93124 531286 93176 531292
rect 94044 531344 94096 531350
rect 94044 531286 94096 531292
rect 93136 522306 93164 531286
rect 93124 522300 93176 522306
rect 93124 522242 93176 522248
rect 92572 515432 92624 515438
rect 92572 515374 92624 515380
rect 91192 471300 91244 471306
rect 91192 471242 91244 471248
rect 90364 469260 90416 469266
rect 90364 469202 90416 469208
rect 91008 469260 91060 469266
rect 91008 469202 91060 469208
rect 90376 458862 90404 469202
rect 90364 458856 90416 458862
rect 90364 458798 90416 458804
rect 89350 436792 89406 436801
rect 89350 436727 89406 436736
rect 88984 436212 89036 436218
rect 88984 436154 89036 436160
rect 89364 434330 89392 436727
rect 89902 436248 89958 436257
rect 89902 436183 89958 436192
rect 89056 434302 89392 434330
rect 88320 434166 88472 434194
rect 89916 434058 89944 436183
rect 92584 434602 92612 515374
rect 93952 483676 94004 483682
rect 93952 483618 94004 483624
rect 93964 441614 93992 483618
rect 94148 476814 94176 539650
rect 94594 538928 94650 538937
rect 94594 538863 94650 538872
rect 94608 538354 94636 538863
rect 94596 538348 94648 538354
rect 94596 538290 94648 538296
rect 94700 534750 94728 558583
rect 94778 540288 94834 540297
rect 94778 540223 94834 540232
rect 94792 539714 94820 540223
rect 94780 539708 94832 539714
rect 94780 539650 94832 539656
rect 94688 534744 94740 534750
rect 94688 534686 94740 534692
rect 94504 522300 94556 522306
rect 94504 522242 94556 522248
rect 94136 476808 94188 476814
rect 94136 476750 94188 476756
rect 94516 465594 94544 522242
rect 95252 512689 95280 563615
rect 95344 558890 95372 588542
rect 95882 582584 95938 582593
rect 95882 582519 95938 582528
rect 95896 576162 95924 582519
rect 95884 576156 95936 576162
rect 95884 576098 95936 576104
rect 95422 565856 95478 565865
rect 95422 565791 95478 565800
rect 95332 558884 95384 558890
rect 95332 558826 95384 558832
rect 95330 555520 95386 555529
rect 95330 555455 95386 555464
rect 95344 520985 95372 555455
rect 95436 535430 95464 565791
rect 96632 552129 96660 702442
rect 105464 700330 105492 703520
rect 137848 702642 137876 703520
rect 154132 702846 154160 703520
rect 154120 702840 154172 702846
rect 154120 702782 154172 702788
rect 137836 702636 137888 702642
rect 137836 702578 137888 702584
rect 170324 702574 170352 703520
rect 202800 703050 202828 703520
rect 218992 703050 219020 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 218980 703044 219032 703050
rect 218980 702986 219032 702992
rect 179328 702976 179380 702982
rect 179328 702918 179380 702924
rect 170312 702568 170364 702574
rect 170312 702510 170364 702516
rect 166356 702500 166408 702506
rect 166356 702442 166408 702448
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 164148 618316 164200 618322
rect 164148 618258 164200 618264
rect 161388 616888 161440 616894
rect 161388 616830 161440 616836
rect 155592 615528 155644 615534
rect 155592 615470 155644 615476
rect 147588 614236 147640 614242
rect 147588 614178 147640 614184
rect 137928 610088 137980 610094
rect 137928 610030 137980 610036
rect 98644 605872 98696 605878
rect 98644 605814 98696 605820
rect 97264 596216 97316 596222
rect 97264 596158 97316 596164
rect 96712 579624 96764 579630
rect 96712 579566 96764 579572
rect 96724 569129 96752 579566
rect 96894 578912 96950 578921
rect 96894 578847 96950 578856
rect 96908 578270 96936 578847
rect 96896 578264 96948 578270
rect 96896 578206 96948 578212
rect 97276 572665 97304 596158
rect 98552 583840 98604 583846
rect 98552 583782 98604 583788
rect 98564 578202 98592 583782
rect 98656 583409 98684 605814
rect 115204 604512 115256 604518
rect 115204 604454 115256 604460
rect 104164 601724 104216 601730
rect 104164 601666 104216 601672
rect 98642 583400 98698 583409
rect 98642 583335 98698 583344
rect 98552 578196 98604 578202
rect 98552 578138 98604 578144
rect 97906 577552 97962 577561
rect 97962 577510 98040 577538
rect 97906 577487 97962 577496
rect 97908 576836 97960 576842
rect 97908 576778 97960 576784
rect 97920 576745 97948 576778
rect 97906 576736 97962 576745
rect 97906 576671 97962 576680
rect 97906 575104 97962 575113
rect 97906 575039 97962 575048
rect 97920 574802 97948 575039
rect 97908 574796 97960 574802
rect 97908 574738 97960 574744
rect 97538 573472 97594 573481
rect 97538 573407 97594 573416
rect 97552 573034 97580 573407
rect 98012 573374 98040 577510
rect 98000 573368 98052 573374
rect 98000 573310 98052 573316
rect 97540 573028 97592 573034
rect 97540 572970 97592 572976
rect 97262 572656 97318 572665
rect 97262 572591 97318 572600
rect 97722 571432 97778 571441
rect 97722 571367 97724 571376
rect 97776 571367 97778 571376
rect 97724 571338 97776 571344
rect 97906 570072 97962 570081
rect 97906 570007 97962 570016
rect 97920 569974 97948 570007
rect 97908 569968 97960 569974
rect 97908 569910 97960 569916
rect 97908 569220 97960 569226
rect 97908 569162 97960 569168
rect 97920 569129 97948 569162
rect 96710 569120 96766 569129
rect 96710 569055 96766 569064
rect 97906 569120 97962 569129
rect 97906 569055 97962 569064
rect 97908 567248 97960 567254
rect 97906 567216 97908 567225
rect 97960 567216 97962 567225
rect 97906 567151 97962 567160
rect 97906 562592 97962 562601
rect 97906 562527 97962 562536
rect 97920 562358 97948 562527
rect 97908 562352 97960 562358
rect 97908 562294 97960 562300
rect 96802 561096 96858 561105
rect 96802 561031 96858 561040
rect 97906 561096 97962 561105
rect 97906 561031 97962 561040
rect 96710 556880 96766 556889
rect 96710 556815 96766 556824
rect 96618 552120 96674 552129
rect 96618 552055 96674 552064
rect 95424 535424 95476 535430
rect 95424 535366 95476 535372
rect 96724 526425 96752 556815
rect 96816 533390 96844 561031
rect 97920 560998 97948 561031
rect 97908 560992 97960 560998
rect 97908 560934 97960 560940
rect 96894 559600 96950 559609
rect 96894 559535 96950 559544
rect 96908 558958 96936 559535
rect 96896 558952 96948 558958
rect 96896 558894 96948 558900
rect 97906 556880 97962 556889
rect 97906 556815 97908 556824
rect 97960 556815 97962 556824
rect 97908 556786 97960 556792
rect 96986 554160 97042 554169
rect 96986 554095 97042 554104
rect 96894 541784 96950 541793
rect 96894 541719 96950 541728
rect 96804 533384 96856 533390
rect 96804 533326 96856 533332
rect 96908 532030 96936 541719
rect 96896 532024 96948 532030
rect 96896 531966 96948 531972
rect 96710 526416 96766 526425
rect 96710 526351 96766 526360
rect 95330 520976 95386 520985
rect 95330 520911 95386 520920
rect 95238 512680 95294 512689
rect 95238 512615 95294 512624
rect 94594 500168 94650 500177
rect 94594 500103 94650 500112
rect 94608 483682 94636 500103
rect 94596 483676 94648 483682
rect 94596 483618 94648 483624
rect 94504 465588 94556 465594
rect 94504 465530 94556 465536
rect 95148 465588 95200 465594
rect 95148 465530 95200 465536
rect 95160 465118 95188 465530
rect 95148 465112 95200 465118
rect 95148 465054 95200 465060
rect 95160 450634 95188 465054
rect 96528 458856 96580 458862
rect 96528 458798 96580 458804
rect 95148 450628 95200 450634
rect 95148 450570 95200 450576
rect 95240 446480 95292 446486
rect 95240 446422 95292 446428
rect 93964 441586 94176 441614
rect 94044 436688 94096 436694
rect 94044 436630 94096 436636
rect 92538 434574 92612 434602
rect 92538 434194 92566 434574
rect 94056 434330 94084 436630
rect 93840 434302 94084 434330
rect 94148 434330 94176 441586
rect 95252 434602 95280 446422
rect 96540 441614 96568 458798
rect 96712 450628 96764 450634
rect 96712 450570 96764 450576
rect 96448 441586 96568 441614
rect 96724 441614 96752 450570
rect 96724 441586 96936 441614
rect 95252 434574 95326 434602
rect 94148 434302 94576 434330
rect 95298 434316 95326 434574
rect 95698 434344 95754 434353
rect 96448 434330 96476 441586
rect 96710 436112 96766 436121
rect 96710 436047 96766 436056
rect 95754 434302 96476 434330
rect 95698 434279 95754 434288
rect 92754 434208 92810 434217
rect 92538 434180 92754 434194
rect 92552 434166 92754 434180
rect 96724 434194 96752 436047
rect 96908 434330 96936 441586
rect 97000 436121 97028 554095
rect 97906 552800 97962 552809
rect 97906 552735 97962 552744
rect 97814 552120 97870 552129
rect 97920 552090 97948 552735
rect 97814 552055 97870 552064
rect 97908 552084 97960 552090
rect 97828 549914 97856 552055
rect 97908 552026 97960 552032
rect 97816 549908 97868 549914
rect 97816 549850 97868 549856
rect 97078 545728 97134 545737
rect 97078 545663 97134 545672
rect 97092 545290 97120 545663
rect 97080 545284 97132 545290
rect 97080 545226 97132 545232
rect 97538 544368 97594 544377
rect 97538 544303 97594 544312
rect 97552 543794 97580 544303
rect 97540 543788 97592 543794
rect 97540 543730 97592 543736
rect 97538 543008 97594 543017
rect 97538 542943 97594 542952
rect 97552 542434 97580 542943
rect 97540 542428 97592 542434
rect 97540 542370 97592 542376
rect 97906 541784 97962 541793
rect 97906 541719 97962 541728
rect 97920 541686 97948 541719
rect 97908 541680 97960 541686
rect 97908 541622 97960 541628
rect 98012 528494 98040 573310
rect 100760 573028 100812 573034
rect 100760 572970 100812 572976
rect 100772 572014 100800 572970
rect 100760 572008 100812 572014
rect 100760 571950 100812 571956
rect 101404 571396 101456 571402
rect 101404 571338 101456 571344
rect 101416 551993 101444 571338
rect 102048 552084 102100 552090
rect 102048 552026 102100 552032
rect 101402 551984 101458 551993
rect 101402 551919 101458 551928
rect 102060 548554 102088 552026
rect 102048 548548 102100 548554
rect 102048 548490 102100 548496
rect 99380 546508 99432 546514
rect 99380 546450 99432 546456
rect 99392 538286 99420 546450
rect 100024 545284 100076 545290
rect 100024 545226 100076 545232
rect 99380 538280 99432 538286
rect 99380 538222 99432 538228
rect 100036 532030 100064 545226
rect 104176 538354 104204 601666
rect 106922 581224 106978 581233
rect 106922 581159 106978 581168
rect 105544 581052 105596 581058
rect 105544 580994 105596 581000
rect 105556 570654 105584 580994
rect 105544 570648 105596 570654
rect 105544 570590 105596 570596
rect 106188 562352 106240 562358
rect 106188 562294 106240 562300
rect 106200 551342 106228 562294
rect 106188 551336 106240 551342
rect 106188 551278 106240 551284
rect 106936 545766 106964 581159
rect 108304 581120 108356 581126
rect 108304 581062 108356 581068
rect 106924 545760 106976 545766
rect 106924 545702 106976 545708
rect 104256 543788 104308 543794
rect 104256 543730 104308 543736
rect 104164 538348 104216 538354
rect 104164 538290 104216 538296
rect 102784 533452 102836 533458
rect 102784 533394 102836 533400
rect 100024 532024 100076 532030
rect 100024 531966 100076 531972
rect 98000 528488 98052 528494
rect 98000 528430 98052 528436
rect 99380 518220 99432 518226
rect 99380 518162 99432 518168
rect 98644 464364 98696 464370
rect 98644 464306 98696 464312
rect 98366 438152 98422 438161
rect 98366 438087 98422 438096
rect 96986 436112 97042 436121
rect 96986 436047 97042 436056
rect 98380 434330 98408 438087
rect 98656 436694 98684 464306
rect 99392 441614 99420 518162
rect 102796 476814 102824 533394
rect 104268 488510 104296 543730
rect 104256 488504 104308 488510
rect 104256 488446 104308 488452
rect 104268 487218 104296 488446
rect 104256 487212 104308 487218
rect 104256 487154 104308 487160
rect 104808 487212 104860 487218
rect 104808 487154 104860 487160
rect 102140 476808 102192 476814
rect 102140 476750 102192 476756
rect 102784 476808 102836 476814
rect 102784 476750 102836 476756
rect 101404 472660 101456 472666
rect 101404 472602 101456 472608
rect 101416 451314 101444 472602
rect 101404 451308 101456 451314
rect 101404 451250 101456 451256
rect 101416 444514 101444 451250
rect 101404 444508 101456 444514
rect 101404 444450 101456 444456
rect 102152 441614 102180 476750
rect 104164 444508 104216 444514
rect 104164 444450 104216 444456
rect 104176 441614 104204 444450
rect 99392 441586 99696 441614
rect 102152 441586 102640 441614
rect 98644 436688 98696 436694
rect 98644 436630 98696 436636
rect 96908 434302 97336 434330
rect 98072 434302 98408 434330
rect 99668 434330 99696 441586
rect 102508 436824 102560 436830
rect 102508 436766 102560 436772
rect 100206 434344 100262 434353
rect 99668 434302 100206 434330
rect 102520 434330 102548 436766
rect 102304 434302 102548 434330
rect 102612 434330 102640 441586
rect 103992 441586 104204 441614
rect 103796 439544 103848 439550
rect 103796 439486 103848 439492
rect 103808 438870 103836 439486
rect 103796 438864 103848 438870
rect 103796 438806 103848 438812
rect 103992 434330 104020 441586
rect 104820 439006 104848 487154
rect 106924 474836 106976 474842
rect 106924 474778 106976 474784
rect 105544 472048 105596 472054
rect 105544 471990 105596 471996
rect 105556 460902 105584 471990
rect 105544 460896 105596 460902
rect 105544 460838 105596 460844
rect 105556 459950 105584 460838
rect 104900 459944 104952 459950
rect 104900 459886 104952 459892
rect 105544 459944 105596 459950
rect 105544 459886 105596 459892
rect 104912 441614 104940 459886
rect 106278 450528 106334 450537
rect 106278 450463 106334 450472
rect 104912 441586 105400 441614
rect 104808 439000 104860 439006
rect 104808 438942 104860 438948
rect 104440 438864 104492 438870
rect 104440 438806 104492 438812
rect 102612 434302 103040 434330
rect 103592 434302 104020 434330
rect 100206 434279 100262 434288
rect 96600 434166 96752 434194
rect 92754 434143 92810 434152
rect 104452 434058 104480 438806
rect 104898 434616 104954 434625
rect 104898 434551 104954 434560
rect 104912 434330 104940 434551
rect 105372 434330 105400 441586
rect 106292 434602 106320 450463
rect 106936 438870 106964 474778
rect 108316 451274 108344 581062
rect 111064 576156 111116 576162
rect 111064 576098 111116 576104
rect 109684 532092 109736 532098
rect 109684 532034 109736 532040
rect 109696 474065 109724 532034
rect 111076 479534 111104 576098
rect 112536 569968 112588 569974
rect 112536 569910 112588 569916
rect 112548 548554 112576 569910
rect 113824 558952 113876 558958
rect 113824 558894 113876 558900
rect 112444 548548 112496 548554
rect 112444 548490 112496 548496
rect 112536 548548 112588 548554
rect 112536 548490 112588 548496
rect 111064 479528 111116 479534
rect 111064 479470 111116 479476
rect 111076 478922 111104 479470
rect 110420 478916 110472 478922
rect 110420 478858 110472 478864
rect 111064 478916 111116 478922
rect 111064 478858 111116 478864
rect 109038 474056 109094 474065
rect 109038 473991 109094 474000
rect 109682 474056 109738 474065
rect 109682 473991 109738 474000
rect 107948 451246 108344 451274
rect 107948 450634 107976 451246
rect 107936 450628 107988 450634
rect 107936 450570 107988 450576
rect 107948 441614 107976 450570
rect 109052 441614 109080 473991
rect 110432 441614 110460 478858
rect 111064 471300 111116 471306
rect 111064 471242 111116 471248
rect 107948 441586 108160 441614
rect 109052 441586 109448 441614
rect 110432 441586 110920 441614
rect 107660 439000 107712 439006
rect 107660 438942 107712 438948
rect 106924 438864 106976 438870
rect 106924 438806 106976 438812
rect 107672 436121 107700 438942
rect 107658 436112 107714 436121
rect 107658 436047 107714 436056
rect 106292 434574 106366 434602
rect 104912 434302 105064 434330
rect 105372 434302 105800 434330
rect 106338 434316 106366 434574
rect 107672 434330 107700 436047
rect 108132 434330 108160 441586
rect 109420 434330 109448 441586
rect 110788 436756 110840 436762
rect 110788 436698 110840 436704
rect 110800 434330 110828 436698
rect 107672 434302 107824 434330
rect 108132 434302 108560 434330
rect 109420 434302 109848 434330
rect 110584 434302 110828 434330
rect 110892 434330 110920 441586
rect 111076 436830 111104 471242
rect 112456 462398 112484 548490
rect 113836 467906 113864 558894
rect 115216 556850 115244 604454
rect 133694 598224 133750 598233
rect 133694 598159 133750 598168
rect 133708 597582 133736 598159
rect 133696 597576 133748 597582
rect 133696 597518 133748 597524
rect 125508 589960 125560 589966
rect 125508 589902 125560 589908
rect 125520 589354 125548 589902
rect 124220 589348 124272 589354
rect 124220 589290 124272 589296
rect 125508 589348 125560 589354
rect 125508 589290 125560 589296
rect 122196 585200 122248 585206
rect 122196 585142 122248 585148
rect 122104 583772 122156 583778
rect 122104 583714 122156 583720
rect 119342 582720 119398 582729
rect 119342 582655 119398 582664
rect 116584 575544 116636 575550
rect 116584 575486 116636 575492
rect 115204 556844 115256 556850
rect 115204 556786 115256 556792
rect 116122 554024 116178 554033
rect 116122 553959 116178 553968
rect 114744 551336 114796 551342
rect 114744 551278 114796 551284
rect 114468 468512 114520 468518
rect 114468 468454 114520 468460
rect 114480 467906 114508 468454
rect 113824 467900 113876 467906
rect 113824 467842 113876 467848
rect 114468 467900 114520 467906
rect 114468 467842 114520 467848
rect 112444 462392 112496 462398
rect 112444 462334 112496 462340
rect 111064 436824 111116 436830
rect 111064 436766 111116 436772
rect 112456 434790 112484 462334
rect 113824 450560 113876 450566
rect 113824 450502 113876 450508
rect 113836 449857 113864 450502
rect 113822 449848 113878 449857
rect 113822 449783 113878 449792
rect 112444 434784 112496 434790
rect 112444 434726 112496 434732
rect 112456 434330 112484 434726
rect 110892 434302 111320 434330
rect 112456 434302 112944 434330
rect 89792 434030 89944 434058
rect 104328 434030 104480 434058
rect 101218 433800 101274 433809
rect 101274 433758 101568 433786
rect 101218 433735 101274 433744
rect 84622 433622 85252 433650
rect 85946 433664 86002 433673
rect 84566 433599 84622 433608
rect 87234 433664 87290 433673
rect 86002 433622 86296 433650
rect 85946 433599 86002 433608
rect 89994 433664 90050 433673
rect 87290 433622 87584 433650
rect 87234 433599 87290 433608
rect 90730 433664 90786 433673
rect 90050 433622 90344 433650
rect 89994 433599 90050 433608
rect 91558 433664 91614 433673
rect 90786 433622 91080 433650
rect 90730 433599 90786 433608
rect 93030 433664 93086 433673
rect 91614 433622 91816 433650
rect 91558 433599 91614 433608
rect 98458 433664 98514 433673
rect 93086 433622 93288 433650
rect 93030 433599 93086 433608
rect 99838 433664 99894 433673
rect 98514 433622 98808 433650
rect 99544 433622 99838 433650
rect 98458 433599 98514 433608
rect 99838 433599 99894 433608
rect 100666 433664 100722 433673
rect 106738 433664 106794 433673
rect 100722 433622 100832 433650
rect 100666 433599 100722 433608
rect 109498 433664 109554 433673
rect 106794 433622 107088 433650
rect 109296 433622 109498 433650
rect 106738 433599 106794 433608
rect 109498 433599 109554 433608
rect 111706 433664 111762 433673
rect 111762 433622 112056 433650
rect 111706 433599 111762 433608
rect 112916 431254 112944 434302
rect 112904 431248 112956 431254
rect 112904 431190 112956 431196
rect 113270 426048 113326 426057
rect 113270 425983 113326 425992
rect 113178 420880 113234 420889
rect 113178 420815 113234 420824
rect 113086 407144 113142 407153
rect 113086 407079 113088 407088
rect 113140 407079 113142 407088
rect 113088 407050 113140 407056
rect 112720 391332 112772 391338
rect 112720 391274 112772 391280
rect 93952 390992 94004 390998
rect 72422 390960 72478 390969
rect 72128 390918 72422 390946
rect 72422 390895 72478 390904
rect 84382 390960 84438 390969
rect 87142 390960 87198 390969
rect 84382 390895 84438 390904
rect 86972 390918 87142 390946
rect 80150 390824 80206 390833
rect 80150 390759 80206 390768
rect 80978 390824 81034 390833
rect 83186 390824 83242 390833
rect 81034 390782 81328 390810
rect 80978 390759 81034 390768
rect 83186 390759 83242 390768
rect 77206 390416 77262 390425
rect 68802 390182 68830 390388
rect 69124 390374 69368 390402
rect 69768 390374 70104 390402
rect 68790 390176 68842 390182
rect 68790 390118 68842 390124
rect 69020 387048 69072 387054
rect 69020 386990 69072 386996
rect 69032 360194 69060 386990
rect 69124 364342 69152 390374
rect 69768 387054 69796 390374
rect 70826 390130 70854 390388
rect 70964 390374 71576 390402
rect 72528 390374 72864 390402
rect 73172 390374 73600 390402
rect 73724 390374 74336 390402
rect 74552 390374 75072 390402
rect 75196 390374 75624 390402
rect 75932 390374 76360 390402
rect 77096 390374 77206 390402
rect 70826 390102 70900 390130
rect 70872 387870 70900 390102
rect 70860 387864 70912 387870
rect 70860 387806 70912 387812
rect 69756 387048 69808 387054
rect 69756 386990 69808 386996
rect 70964 373994 70992 390374
rect 71044 388476 71096 388482
rect 71044 388418 71096 388424
rect 70412 373966 70992 373994
rect 70412 369073 70440 373966
rect 70398 369064 70454 369073
rect 70398 368999 70454 369008
rect 71056 368422 71084 388418
rect 71688 388408 71740 388414
rect 71688 388350 71740 388356
rect 71700 388006 71728 388350
rect 72528 388006 72556 390374
rect 71688 388000 71740 388006
rect 71688 387942 71740 387948
rect 72516 388000 72568 388006
rect 72516 387942 72568 387948
rect 71700 384985 71728 387942
rect 72516 387864 72568 387870
rect 72516 387806 72568 387812
rect 72422 385112 72478 385121
rect 72422 385047 72478 385056
rect 71686 384976 71742 384985
rect 71686 384911 71742 384920
rect 71688 369164 71740 369170
rect 71688 369106 71740 369112
rect 71700 369073 71728 369106
rect 71686 369064 71742 369073
rect 71686 368999 71742 369008
rect 71044 368416 71096 368422
rect 71044 368358 71096 368364
rect 69112 364336 69164 364342
rect 69112 364278 69164 364284
rect 69020 360188 69072 360194
rect 69020 360130 69072 360136
rect 69664 360188 69716 360194
rect 69664 360130 69716 360136
rect 68664 306346 68876 306374
rect 68284 287768 68336 287774
rect 68284 287710 68336 287716
rect 67548 283076 67600 283082
rect 67548 283018 67600 283024
rect 67560 279721 67588 283018
rect 67914 280528 67970 280537
rect 67914 280463 67970 280472
rect 67546 279712 67602 279721
rect 67546 279647 67602 279656
rect 67548 278316 67600 278322
rect 67548 278258 67600 278264
rect 67560 278089 67588 278258
rect 67546 278080 67602 278089
rect 67546 278015 67602 278024
rect 67454 263392 67510 263401
rect 67454 263327 67510 263336
rect 67362 256864 67418 256873
rect 67362 256799 67418 256808
rect 67272 253224 67324 253230
rect 67272 253166 67324 253172
rect 66996 250504 67048 250510
rect 66996 250446 67048 250452
rect 66904 249076 66956 249082
rect 66904 249018 66956 249024
rect 66916 248713 66944 249018
rect 66902 248704 66958 248713
rect 66902 248639 66958 248648
rect 66904 244248 66956 244254
rect 66904 244190 66956 244196
rect 66916 243001 66944 244190
rect 66902 242992 66958 243001
rect 66902 242927 66958 242936
rect 66902 242176 66958 242185
rect 66902 242111 66958 242120
rect 66916 241534 66944 242111
rect 66904 241528 66956 241534
rect 66904 241470 66956 241476
rect 67284 146334 67312 253166
rect 67822 249520 67878 249529
rect 67822 249455 67878 249464
rect 67362 247072 67418 247081
rect 67362 247007 67418 247016
rect 67376 225010 67404 247007
rect 67454 246256 67510 246265
rect 67454 246191 67510 246200
rect 67468 234569 67496 246191
rect 67638 240136 67694 240145
rect 67638 240071 67694 240080
rect 67454 234560 67510 234569
rect 67454 234495 67510 234504
rect 67364 225004 67416 225010
rect 67364 224946 67416 224952
rect 67272 146328 67324 146334
rect 67272 146270 67324 146276
rect 66732 132466 66852 132494
rect 66732 129849 66760 132466
rect 66904 132456 66956 132462
rect 66904 132398 66956 132404
rect 66812 132388 66864 132394
rect 66812 132330 66864 132336
rect 66824 131209 66852 132330
rect 66916 132025 66944 132398
rect 66902 132016 66958 132025
rect 66902 131951 66958 131960
rect 66810 131200 66866 131209
rect 66810 131135 66866 131144
rect 66812 131096 66864 131102
rect 66812 131038 66864 131044
rect 66824 130665 66852 131038
rect 66810 130656 66866 130665
rect 66810 130591 66866 130600
rect 66718 129840 66774 129849
rect 66718 129775 66774 129784
rect 66810 129024 66866 129033
rect 66810 128959 66866 128968
rect 66824 128382 66852 128959
rect 66812 128376 66864 128382
rect 66812 128318 66864 128324
rect 66812 126948 66864 126954
rect 66812 126890 66864 126896
rect 66824 126857 66852 126890
rect 66810 126848 66866 126857
rect 66810 126783 66866 126792
rect 66074 126032 66130 126041
rect 66074 125967 66130 125976
rect 66812 124976 66864 124982
rect 66812 124918 66864 124924
rect 66824 124409 66852 124918
rect 66996 124908 67048 124914
rect 66996 124850 67048 124856
rect 66810 124400 66866 124409
rect 66810 124335 66866 124344
rect 66904 124160 66956 124166
rect 66904 124102 66956 124108
rect 66916 123049 66944 124102
rect 67008 123865 67036 124850
rect 66994 123856 67050 123865
rect 66994 123791 67050 123800
rect 66902 123040 66958 123049
rect 66902 122975 66958 122984
rect 66352 122800 66404 122806
rect 66352 122742 66404 122748
rect 66364 122233 66392 122742
rect 66350 122224 66406 122233
rect 66350 122159 66406 122168
rect 66904 121440 66956 121446
rect 66810 121408 66866 121417
rect 66904 121382 66956 121388
rect 66810 121343 66812 121352
rect 66864 121343 66866 121352
rect 66812 121314 66864 121320
rect 66916 120601 66944 121382
rect 66902 120592 66958 120601
rect 66902 120527 66958 120536
rect 66812 120080 66864 120086
rect 66810 120048 66812 120057
rect 66864 120048 66866 120057
rect 66810 119983 66866 119992
rect 66904 120012 66956 120018
rect 66904 119954 66956 119960
rect 66916 119241 66944 119954
rect 66902 119232 66958 119241
rect 66902 119167 66958 119176
rect 66628 118652 66680 118658
rect 66628 118594 66680 118600
rect 66640 117609 66668 118594
rect 66626 117600 66682 117609
rect 66626 117535 66682 117544
rect 66628 117292 66680 117298
rect 66628 117234 66680 117240
rect 66640 116249 66668 117234
rect 66626 116240 66682 116249
rect 66626 116175 66682 116184
rect 66812 115932 66864 115938
rect 66812 115874 66864 115880
rect 66824 115433 66852 115874
rect 66904 115592 66956 115598
rect 66904 115534 66956 115540
rect 66810 115424 66866 115433
rect 66810 115359 66866 115368
rect 66916 114617 66944 115534
rect 66902 114608 66958 114617
rect 66902 114543 66958 114552
rect 66812 114504 66864 114510
rect 66812 114446 66864 114452
rect 66824 113801 66852 114446
rect 66904 113824 66956 113830
rect 66810 113792 66866 113801
rect 66904 113766 66956 113772
rect 66810 113727 66866 113736
rect 66916 113257 66944 113766
rect 66902 113248 66958 113257
rect 66902 113183 66958 113192
rect 66812 113144 66864 113150
rect 66812 113086 66864 113092
rect 66824 112441 66852 113086
rect 66810 112432 66866 112441
rect 66810 112367 66866 112376
rect 66812 111784 66864 111790
rect 66812 111726 66864 111732
rect 66824 111625 66852 111726
rect 66810 111616 66866 111625
rect 66810 111551 66866 111560
rect 66904 111104 66956 111110
rect 66904 111046 66956 111052
rect 66916 110809 66944 111046
rect 66902 110800 66958 110809
rect 66902 110735 66958 110744
rect 66902 110256 66958 110265
rect 66902 110191 66958 110200
rect 66916 109070 66944 110191
rect 66904 109064 66956 109070
rect 66904 109006 66956 109012
rect 66812 108996 66864 109002
rect 66812 108938 66864 108944
rect 66074 108624 66130 108633
rect 66074 108559 66130 108568
rect 65890 103184 65946 103193
rect 65890 103119 65946 103128
rect 64788 99680 64840 99686
rect 64788 99622 64840 99628
rect 64694 85504 64750 85513
rect 64694 85439 64750 85448
rect 64800 73166 64828 99622
rect 65524 96688 65576 96694
rect 65524 96630 65576 96636
rect 65536 77246 65564 96630
rect 66088 79966 66116 108559
rect 66824 107817 66852 108938
rect 66810 107808 66866 107817
rect 66810 107743 66866 107752
rect 66628 107636 66680 107642
rect 66628 107578 66680 107584
rect 66640 106457 66668 107578
rect 66810 106992 66866 107001
rect 66810 106927 66866 106936
rect 66626 106448 66682 106457
rect 66626 106383 66682 106392
rect 66824 106350 66852 106927
rect 66812 106344 66864 106350
rect 66812 106286 66864 106292
rect 66626 105632 66682 105641
rect 66168 105596 66220 105602
rect 66626 105567 66628 105576
rect 66168 105538 66220 105544
rect 66680 105567 66682 105576
rect 66628 105538 66680 105544
rect 66076 79960 66128 79966
rect 66076 79902 66128 79908
rect 66180 78577 66208 105538
rect 66812 104848 66864 104854
rect 66810 104816 66812 104825
rect 66864 104816 66866 104825
rect 66810 104751 66866 104760
rect 67284 104009 67312 146270
rect 67270 104000 67326 104009
rect 67270 103935 67326 103944
rect 66444 103420 66496 103426
rect 66444 103362 66496 103368
rect 66456 102649 66484 103362
rect 66442 102640 66498 102649
rect 66442 102575 66498 102584
rect 66718 101824 66774 101833
rect 66718 101759 66774 101768
rect 66732 101454 66760 101759
rect 66720 101448 66772 101454
rect 66720 101390 66772 101396
rect 66810 101008 66866 101017
rect 66810 100943 66866 100952
rect 66824 100774 66852 100943
rect 66812 100768 66864 100774
rect 66812 100710 66864 100716
rect 66812 99680 66864 99686
rect 66810 99648 66812 99657
rect 66864 99648 66866 99657
rect 66810 99583 66866 99592
rect 66812 99340 66864 99346
rect 66812 99282 66864 99288
rect 66824 98841 66852 99282
rect 66810 98832 66866 98841
rect 66810 98767 66866 98776
rect 67376 98025 67404 224946
rect 67468 113174 67496 234495
rect 67546 149152 67602 149161
rect 67546 149087 67548 149096
rect 67600 149087 67602 149096
rect 67548 149058 67600 149064
rect 67652 113174 67680 240071
rect 67836 237386 67864 249455
rect 67824 237380 67876 237386
rect 67824 237322 67876 237328
rect 67928 236609 67956 280463
rect 68296 273290 68324 287710
rect 68466 285968 68522 285977
rect 68466 285903 68522 285912
rect 68480 277394 68508 285903
rect 68652 283280 68704 283286
rect 68652 283222 68704 283228
rect 68560 282192 68612 282198
rect 68558 282160 68560 282169
rect 68612 282160 68614 282169
rect 68558 282095 68614 282104
rect 68480 277366 68600 277394
rect 68284 273284 68336 273290
rect 68284 273226 68336 273232
rect 68190 258768 68246 258777
rect 68190 258703 68246 258712
rect 68204 258058 68232 258703
rect 68192 258052 68244 258058
rect 68192 257994 68244 258000
rect 68572 237998 68600 277366
rect 68664 240650 68692 283222
rect 68848 282690 68876 306346
rect 69202 304192 69258 304201
rect 69202 304127 69258 304136
rect 69020 285864 69072 285870
rect 69020 285806 69072 285812
rect 69032 285734 69060 285806
rect 69020 285728 69072 285734
rect 69020 285670 69072 285676
rect 69032 283778 69060 285670
rect 69216 283801 69244 304127
rect 69676 303657 69704 360130
rect 71964 345636 72016 345642
rect 71964 345578 72016 345584
rect 71042 313984 71098 313993
rect 71042 313919 71098 313928
rect 70306 307728 70362 307737
rect 70306 307663 70362 307672
rect 69662 303648 69718 303657
rect 69662 303583 69718 303592
rect 69664 294024 69716 294030
rect 69664 293966 69716 293972
rect 68986 283750 69060 283778
rect 69202 283792 69258 283801
rect 68986 283492 69014 283750
rect 69202 283727 69258 283736
rect 69388 283280 69440 283286
rect 69440 283228 69552 283234
rect 69388 283222 69552 283228
rect 69400 283206 69552 283222
rect 69676 283014 69704 293966
rect 70076 283792 70132 283801
rect 70076 283727 70132 283736
rect 70090 283506 70118 283727
rect 70214 283520 70270 283529
rect 70090 283492 70214 283506
rect 70104 283478 70214 283492
rect 70214 283455 70270 283464
rect 70320 283286 70348 307663
rect 71056 288386 71084 313919
rect 71136 307148 71188 307154
rect 71136 307090 71188 307096
rect 70584 288380 70636 288386
rect 70584 288322 70636 288328
rect 71044 288380 71096 288386
rect 71044 288322 71096 288328
rect 70596 283778 70624 288322
rect 71148 283778 71176 307090
rect 71872 290488 71924 290494
rect 71872 290430 71924 290436
rect 71884 284374 71912 290430
rect 71872 284368 71924 284374
rect 71872 284310 71924 284316
rect 70596 283750 70670 283778
rect 71148 283750 71222 283778
rect 70642 283492 70670 283750
rect 71194 283370 71222 283750
rect 71884 283506 71912 284310
rect 71976 283801 72004 345578
rect 72436 285734 72464 385047
rect 72528 378146 72556 387806
rect 73066 387696 73122 387705
rect 73066 387631 73122 387640
rect 72516 378140 72568 378146
rect 72516 378082 72568 378088
rect 73080 345642 73108 387631
rect 73172 361554 73200 390374
rect 73724 373994 73752 390374
rect 73264 373966 73752 373994
rect 73264 365702 73292 373966
rect 74552 373318 74580 390374
rect 75196 383654 75224 390374
rect 75932 386356 75960 390374
rect 77206 390351 77262 390360
rect 77496 390374 77832 390402
rect 78048 390374 78384 390402
rect 78784 390374 79120 390402
rect 79520 390374 79856 390402
rect 77220 388793 77248 390351
rect 77206 388784 77262 388793
rect 77206 388719 77262 388728
rect 77390 388512 77446 388521
rect 77390 388447 77446 388456
rect 77208 387864 77260 387870
rect 77208 387806 77260 387812
rect 75840 386328 75960 386356
rect 75196 383626 75316 383654
rect 75184 382968 75236 382974
rect 75184 382910 75236 382916
rect 74540 373312 74592 373318
rect 74540 373254 74592 373260
rect 75196 366994 75224 382910
rect 75288 380866 75316 383626
rect 75276 380860 75328 380866
rect 75276 380802 75328 380808
rect 75184 366988 75236 366994
rect 75184 366930 75236 366936
rect 73252 365696 73304 365702
rect 73252 365638 73304 365644
rect 73160 361548 73212 361554
rect 73160 361490 73212 361496
rect 75840 356046 75868 386328
rect 77220 376650 77248 387806
rect 77208 376644 77260 376650
rect 77208 376586 77260 376592
rect 77220 376106 77248 376586
rect 75920 376100 75972 376106
rect 75920 376042 75972 376048
rect 77208 376100 77260 376106
rect 77208 376042 77260 376048
rect 75932 371890 75960 376042
rect 77208 373380 77260 373386
rect 77208 373322 77260 373328
rect 75920 371884 75972 371890
rect 75920 371826 75972 371832
rect 75184 356040 75236 356046
rect 75184 355982 75236 355988
rect 75828 356040 75880 356046
rect 75828 355982 75880 355988
rect 73068 345636 73120 345642
rect 73068 345578 73120 345584
rect 73080 345098 73108 345578
rect 73068 345092 73120 345098
rect 73068 345034 73120 345040
rect 73804 312588 73856 312594
rect 73804 312530 73856 312536
rect 73068 302252 73120 302258
rect 73068 302194 73120 302200
rect 73080 292574 73108 302194
rect 72712 292546 73108 292574
rect 72424 285728 72476 285734
rect 72424 285670 72476 285676
rect 71962 283792 72018 283801
rect 71962 283727 72018 283736
rect 72712 283506 72740 292546
rect 73816 285870 73844 312530
rect 74632 307080 74684 307086
rect 74632 307022 74684 307028
rect 74644 287842 74672 307022
rect 75196 291854 75224 355982
rect 77220 321473 77248 373322
rect 77206 321464 77262 321473
rect 77206 321399 77262 321408
rect 77220 321065 77248 321399
rect 75918 321056 75974 321065
rect 75918 320991 75974 321000
rect 77206 321056 77262 321065
rect 77206 320991 77262 321000
rect 75276 317416 75328 317422
rect 75276 317358 75328 317364
rect 75184 291848 75236 291854
rect 75184 291790 75236 291796
rect 74632 287836 74684 287842
rect 74632 287778 74684 287784
rect 73804 285864 73856 285870
rect 73804 285806 73856 285812
rect 72836 283792 72892 283801
rect 72836 283727 72892 283736
rect 71760 283478 71912 283506
rect 71976 283478 72740 283506
rect 72850 283492 72878 283727
rect 73816 283506 73844 285806
rect 74630 285560 74686 285569
rect 74630 285495 74686 285504
rect 74644 284345 74672 285495
rect 75288 284481 75316 317358
rect 75932 306374 75960 320991
rect 77404 307154 77432 388447
rect 77496 381546 77524 390374
rect 78048 387870 78076 390374
rect 78036 387864 78088 387870
rect 78036 387806 78088 387812
rect 78680 387048 78732 387054
rect 78680 386990 78732 386996
rect 77484 381540 77536 381546
rect 77484 381482 77536 381488
rect 78692 376038 78720 386990
rect 78784 382974 78812 390374
rect 79520 387054 79548 390374
rect 79508 387048 79560 387054
rect 79508 386990 79560 386996
rect 78772 382968 78824 382974
rect 78772 382910 78824 382916
rect 78680 376032 78732 376038
rect 80164 376009 80192 390759
rect 83200 390674 83228 390759
rect 83200 390646 83352 390674
rect 82174 390552 82230 390561
rect 81728 390510 82174 390538
rect 80592 390374 80928 390402
rect 80242 388512 80298 388521
rect 80242 388447 80298 388456
rect 78680 375974 78732 375980
rect 80150 376000 80206 376009
rect 80150 375935 80206 375944
rect 78586 313984 78642 313993
rect 78586 313919 78642 313928
rect 77392 307148 77444 307154
rect 77392 307090 77444 307096
rect 77298 306640 77354 306649
rect 77298 306575 77354 306584
rect 75932 306346 76328 306374
rect 75458 292632 75514 292641
rect 75458 292567 75514 292576
rect 75368 287836 75420 287842
rect 75368 287778 75420 287784
rect 75274 284472 75330 284481
rect 75274 284407 75330 284416
rect 74630 284336 74686 284345
rect 74630 284271 74686 284280
rect 73816 283478 73968 283506
rect 70964 283356 71222 283370
rect 70964 283342 71208 283356
rect 70308 283280 70360 283286
rect 70964 283257 70992 283342
rect 71976 283257 72004 283478
rect 74644 283370 74672 284271
rect 75288 283370 75316 284407
rect 75380 283506 75408 287778
rect 75472 285569 75500 292567
rect 76196 289468 76248 289474
rect 76196 289410 76248 289416
rect 76208 288454 76236 289410
rect 76196 288448 76248 288454
rect 76196 288390 76248 288396
rect 75458 285560 75514 285569
rect 75458 285495 75514 285504
rect 76208 283778 76236 288390
rect 76162 283750 76236 283778
rect 75380 283478 75624 283506
rect 76162 283492 76190 283750
rect 76300 283506 76328 306346
rect 76562 303648 76618 303657
rect 76562 303583 76618 303592
rect 76576 289474 76604 303583
rect 76564 289468 76616 289474
rect 76564 289410 76616 289416
rect 77312 283778 77340 306575
rect 78600 296714 78628 313919
rect 80256 312594 80284 388447
rect 80900 385665 80928 390374
rect 81728 389230 81756 390510
rect 82174 390487 82230 390496
rect 82616 390374 82768 390402
rect 81716 389224 81768 389230
rect 81716 389166 81768 389172
rect 81438 388512 81494 388521
rect 82740 388482 82768 390374
rect 81438 388447 81494 388456
rect 82728 388476 82780 388482
rect 80886 385656 80942 385665
rect 80886 385591 80942 385600
rect 81452 317422 81480 388447
rect 82728 388418 82780 388424
rect 83200 387938 83228 390646
rect 83476 390374 84088 390402
rect 83188 387932 83240 387938
rect 83188 387874 83240 387880
rect 83476 387002 83504 390374
rect 84396 389174 84424 390895
rect 84824 390374 84976 390402
rect 84304 389146 84424 389174
rect 84108 387932 84160 387938
rect 84108 387874 84160 387880
rect 83554 387288 83610 387297
rect 83554 387223 83610 387232
rect 82832 386974 83504 387002
rect 82832 379506 82860 386974
rect 82820 379500 82872 379506
rect 82820 379442 82872 379448
rect 83568 373994 83596 387223
rect 83476 373966 83596 373994
rect 82726 339552 82782 339561
rect 82726 339487 82728 339496
rect 82780 339487 82782 339496
rect 82728 339458 82780 339464
rect 81440 317416 81492 317422
rect 81440 317358 81492 317364
rect 82726 316704 82782 316713
rect 82726 316639 82782 316648
rect 80244 312588 80296 312594
rect 80244 312530 80296 312536
rect 79966 311128 80022 311137
rect 79966 311063 80022 311072
rect 78508 296686 78628 296714
rect 78508 292574 78536 296686
rect 78232 292546 78536 292574
rect 78232 284481 78260 292546
rect 79980 288454 80008 311063
rect 80060 305040 80112 305046
rect 80060 304982 80112 304988
rect 79232 288448 79284 288454
rect 79232 288390 79284 288396
rect 79968 288448 80020 288454
rect 79968 288390 80020 288396
rect 78588 287700 78640 287706
rect 78588 287642 78640 287648
rect 78218 284472 78274 284481
rect 78218 284407 78274 284416
rect 77266 283750 77340 283778
rect 76300 283478 76728 283506
rect 77266 283492 77294 283750
rect 78232 283506 78260 284407
rect 78600 283506 78628 287642
rect 79244 283506 79272 288390
rect 79322 287056 79378 287065
rect 79322 286991 79378 287000
rect 79336 285977 79364 286991
rect 79322 285968 79378 285977
rect 79322 285903 79378 285912
rect 77832 283478 78260 283506
rect 78384 283478 78628 283506
rect 78936 283478 79272 283506
rect 79336 283506 79364 285903
rect 80072 283778 80100 304982
rect 82634 300248 82690 300257
rect 82634 300183 82690 300192
rect 80886 289912 80942 289921
rect 80886 289847 80942 289856
rect 80428 286476 80480 286482
rect 80428 286418 80480 286424
rect 80440 285841 80468 286418
rect 80426 285832 80482 285841
rect 80426 285767 80482 285776
rect 80026 283750 80100 283778
rect 79336 283478 79488 283506
rect 80026 283492 80054 283750
rect 80900 283506 80928 289847
rect 81256 286476 81308 286482
rect 81256 286418 81308 286424
rect 80592 283478 80928 283506
rect 81268 283370 81296 286418
rect 81992 286136 82044 286142
rect 81992 286078 82044 286084
rect 82004 283506 82032 286078
rect 82648 285841 82676 300183
rect 82740 286142 82768 316639
rect 82912 311160 82964 311166
rect 82912 311102 82964 311108
rect 82924 306374 82952 311102
rect 82924 306346 83412 306374
rect 82728 286136 82780 286142
rect 82728 286078 82780 286084
rect 83094 285968 83150 285977
rect 83094 285903 83150 285912
rect 82634 285832 82690 285841
rect 82634 285767 82690 285776
rect 82648 283506 82676 285767
rect 83108 283506 83136 285903
rect 83384 285818 83412 306346
rect 83476 286482 83504 373966
rect 84120 372502 84148 387874
rect 84304 373386 84332 389146
rect 84948 386374 84976 390374
rect 85040 390374 85376 390402
rect 85592 390374 86112 390402
rect 85040 388385 85068 390374
rect 85026 388376 85082 388385
rect 85026 388311 85082 388320
rect 84936 386368 84988 386374
rect 84936 386310 84988 386316
rect 84292 373380 84344 373386
rect 84292 373322 84344 373328
rect 84108 372496 84160 372502
rect 84108 372438 84160 372444
rect 85592 371142 85620 390374
rect 86834 390130 86862 390388
rect 86834 390102 86908 390130
rect 86880 387161 86908 390102
rect 86866 387152 86922 387161
rect 86866 387087 86922 387096
rect 86972 376553 87000 390918
rect 87142 390895 87198 390904
rect 87878 390960 87934 390969
rect 87934 390918 88136 390946
rect 93952 390934 94004 390940
rect 94964 390992 95016 390998
rect 107292 390992 107344 390998
rect 99654 390960 99710 390969
rect 95016 390940 95128 390946
rect 94964 390934 95128 390940
rect 87878 390895 87934 390904
rect 92018 390416 92074 390425
rect 87064 390374 87584 390402
rect 88352 390374 88872 390402
rect 89272 390374 89608 390402
rect 89732 390374 90344 390402
rect 91080 390374 91324 390402
rect 87064 383382 87092 390374
rect 88248 387796 88300 387802
rect 88248 387738 88300 387744
rect 87052 383376 87104 383382
rect 87052 383318 87104 383324
rect 86958 376544 87014 376553
rect 86958 376479 87014 376488
rect 85580 371136 85632 371142
rect 85580 371078 85632 371084
rect 84106 370560 84162 370569
rect 84106 370495 84162 370504
rect 84014 304192 84070 304201
rect 84014 304127 84070 304136
rect 83464 286476 83516 286482
rect 83464 286418 83516 286424
rect 83384 285790 83504 285818
rect 81696 283478 82032 283506
rect 82248 283478 82676 283506
rect 82800 283478 83136 283506
rect 83476 283506 83504 285790
rect 83476 283478 83904 283506
rect 74520 283342 74672 283370
rect 75072 283342 75316 283370
rect 81144 283342 81296 283370
rect 84028 283286 84056 304127
rect 84120 285977 84148 370495
rect 84200 350600 84252 350606
rect 84200 350542 84252 350548
rect 84106 285968 84162 285977
rect 84106 285903 84162 285912
rect 84212 283506 84240 350542
rect 88260 350538 88288 387738
rect 88352 374678 88380 390374
rect 89272 386306 89300 390374
rect 88432 386300 88484 386306
rect 88432 386242 88484 386248
rect 89260 386300 89312 386306
rect 89260 386242 89312 386248
rect 88444 379409 88472 386242
rect 89626 385792 89682 385801
rect 89626 385727 89682 385736
rect 88430 379400 88486 379409
rect 88430 379335 88486 379344
rect 88340 374672 88392 374678
rect 88340 374614 88392 374620
rect 88248 350532 88300 350538
rect 88248 350474 88300 350480
rect 88260 317393 88288 350474
rect 88984 324964 89036 324970
rect 88984 324906 89036 324912
rect 87602 317384 87658 317393
rect 87602 317319 87658 317328
rect 88246 317384 88302 317393
rect 88246 317319 88302 317328
rect 87616 316169 87644 317319
rect 87602 316160 87658 316169
rect 87602 316095 87658 316104
rect 86866 313984 86922 313993
rect 86866 313919 86922 313928
rect 86774 304328 86830 304337
rect 86774 304263 86830 304272
rect 86224 301572 86276 301578
rect 86224 301514 86276 301520
rect 84568 292596 84620 292602
rect 84568 292538 84620 292544
rect 84580 283506 84608 292538
rect 85854 287192 85910 287201
rect 85854 287127 85910 287136
rect 84660 286136 84712 286142
rect 84660 286078 84712 286084
rect 84672 285569 84700 286078
rect 84658 285560 84714 285569
rect 84658 285495 84714 285504
rect 85868 283506 85896 287127
rect 86086 283756 86138 283762
rect 86086 283698 86138 283704
rect 84212 283478 84456 283506
rect 84580 283478 85008 283506
rect 85560 283478 85896 283506
rect 86098 283492 86126 283698
rect 86236 283506 86264 301514
rect 86788 287201 86816 304263
rect 86774 287192 86830 287201
rect 86774 287127 86830 287136
rect 86880 283762 86908 313919
rect 87512 285728 87564 285734
rect 87512 285670 87564 285676
rect 86868 283756 86920 283762
rect 86868 283698 86920 283704
rect 86880 283665 86908 283698
rect 86866 283656 86922 283665
rect 86866 283591 86922 283600
rect 87524 283506 87552 285670
rect 87616 284986 87644 316095
rect 88246 308544 88302 308553
rect 88246 308479 88302 308488
rect 88260 292574 88288 308479
rect 88996 305658 89024 324906
rect 89536 315308 89588 315314
rect 89536 315250 89588 315256
rect 88984 305652 89036 305658
rect 88984 305594 89036 305600
rect 89548 297226 89576 315250
rect 88432 297220 88484 297226
rect 88432 297162 88484 297168
rect 89536 297220 89588 297226
rect 89536 297162 89588 297168
rect 88168 292546 88288 292574
rect 87604 284980 87656 284986
rect 87604 284922 87656 284928
rect 88168 284374 88196 292546
rect 88156 284368 88208 284374
rect 88156 284310 88208 284316
rect 88168 283506 88196 284310
rect 86236 283478 86664 283506
rect 87216 283478 87552 283506
rect 87768 283478 88196 283506
rect 88444 283506 88472 297162
rect 89548 296750 89576 297162
rect 89536 296744 89588 296750
rect 89536 296686 89588 296692
rect 89640 292574 89668 385727
rect 89732 311273 89760 390374
rect 91296 384305 91324 390374
rect 91388 390374 91632 390402
rect 91282 384296 91338 384305
rect 91282 384231 91338 384240
rect 91284 383376 91336 383382
rect 91284 383318 91336 383324
rect 90362 329896 90418 329905
rect 90362 329831 90418 329840
rect 89718 311264 89774 311273
rect 89718 311199 89774 311208
rect 89548 292546 89668 292574
rect 89548 291242 89576 292546
rect 89536 291236 89588 291242
rect 89536 291178 89588 291184
rect 88982 287736 89038 287745
rect 88982 287671 89038 287680
rect 88444 283478 88872 283506
rect 88996 283422 89024 287671
rect 89548 283506 89576 291178
rect 90270 286104 90326 286113
rect 90270 286039 90326 286048
rect 89424 283478 89576 283506
rect 89810 283520 89866 283529
rect 90284 283506 90312 286039
rect 90376 285734 90404 329831
rect 91006 312488 91062 312497
rect 91006 312423 91062 312432
rect 91020 286113 91048 312423
rect 91192 305652 91244 305658
rect 91192 305594 91244 305600
rect 91006 286104 91062 286113
rect 91006 286039 91062 286048
rect 90364 285728 90416 285734
rect 90364 285670 90416 285676
rect 90824 285728 90876 285734
rect 90824 285670 90876 285676
rect 90836 283506 90864 285670
rect 91100 284436 91152 284442
rect 91100 284378 91152 284384
rect 91112 283778 91140 284378
rect 89866 283478 90312 283506
rect 90528 283478 90864 283506
rect 91066 283750 91140 283778
rect 91066 283492 91094 283750
rect 91204 283506 91232 305594
rect 91296 285569 91324 383318
rect 91388 307737 91416 390374
rect 93964 390402 93992 390934
rect 94976 390918 95128 390934
rect 104254 390960 104310 390969
rect 104144 390918 104254 390946
rect 99654 390895 99710 390904
rect 105266 390960 105322 390969
rect 104310 390918 104572 390946
rect 104254 390895 104310 390904
rect 96986 390416 97042 390425
rect 92074 390374 92368 390402
rect 93104 390374 93440 390402
rect 93840 390374 93992 390402
rect 92018 390351 92074 390360
rect 92032 387802 92060 390351
rect 93412 387802 93440 390374
rect 92020 387796 92072 387802
rect 92020 387738 92072 387744
rect 93400 387796 93452 387802
rect 93400 387738 93452 387744
rect 93860 387048 93912 387054
rect 93860 386990 93912 386996
rect 93766 382936 93822 382945
rect 93766 382871 93822 382880
rect 92478 311944 92534 311953
rect 92478 311879 92534 311888
rect 91374 307728 91430 307737
rect 91374 307663 91430 307672
rect 92492 287842 92520 311879
rect 93780 293962 93808 382871
rect 93872 362234 93900 386990
rect 93964 377466 93992 390374
rect 94148 390374 94392 390402
rect 95252 390374 95864 390402
rect 96600 390374 96936 390402
rect 94148 387054 94176 390374
rect 94136 387048 94188 387054
rect 94136 386990 94188 386996
rect 93952 377460 94004 377466
rect 93952 377402 94004 377408
rect 93860 362228 93912 362234
rect 93860 362170 93912 362176
rect 95146 313984 95202 313993
rect 95146 313919 95202 313928
rect 94502 311128 94558 311137
rect 94502 311063 94558 311072
rect 92572 293956 92624 293962
rect 92572 293898 92624 293904
rect 93768 293956 93820 293962
rect 93768 293898 93820 293904
rect 92480 287836 92532 287842
rect 92480 287778 92532 287784
rect 91282 285560 91338 285569
rect 91282 285495 91338 285504
rect 92584 283506 92612 293898
rect 92940 287836 92992 287842
rect 92940 287778 92992 287784
rect 92952 283506 92980 287778
rect 93950 285696 94006 285705
rect 93950 285631 94006 285640
rect 93964 283506 93992 285631
rect 91204 283478 91632 283506
rect 92584 283478 92736 283506
rect 92952 283478 93288 283506
rect 93840 283478 93992 283506
rect 94042 283520 94098 283529
rect 89810 283455 89866 283464
rect 94516 283506 94544 311063
rect 94098 283478 94544 283506
rect 94686 283520 94742 283529
rect 94042 283455 94098 283464
rect 95160 283506 95188 313919
rect 95252 288561 95280 390374
rect 96908 384334 96936 390374
rect 97042 390374 97488 390402
rect 96986 390351 97042 390360
rect 96896 384328 96948 384334
rect 96896 384270 96948 384276
rect 97460 382974 97488 390374
rect 97552 390374 97888 390402
rect 98624 390374 98960 390402
rect 97552 387841 97580 390374
rect 98932 389230 98960 390374
rect 99346 390130 99374 390388
rect 99300 390102 99374 390130
rect 98920 389224 98972 389230
rect 99300 389201 99328 390102
rect 98920 389166 98972 389172
rect 99286 389192 99342 389201
rect 99668 389174 99696 390895
rect 103794 390824 103850 390833
rect 103592 390782 103794 390810
rect 103794 390759 103850 390768
rect 100096 390374 100432 390402
rect 99286 389127 99342 389136
rect 99484 389146 99696 389174
rect 97538 387832 97594 387841
rect 97538 387767 97594 387776
rect 97264 382968 97316 382974
rect 97264 382910 97316 382916
rect 97448 382968 97500 382974
rect 97448 382910 97500 382916
rect 97276 369850 97304 382910
rect 99300 382129 99328 389127
rect 99286 382120 99342 382129
rect 99286 382055 99342 382064
rect 99286 370696 99342 370705
rect 99286 370631 99342 370640
rect 97264 369844 97316 369850
rect 97264 369786 97316 369792
rect 96712 327752 96764 327758
rect 96712 327694 96764 327700
rect 95330 307048 95386 307057
rect 95330 306983 95386 306992
rect 95344 306374 95372 306983
rect 95344 306346 95648 306374
rect 95238 288552 95294 288561
rect 95238 288487 95294 288496
rect 95332 286136 95384 286142
rect 95332 286078 95384 286084
rect 94742 283478 95188 283506
rect 94686 283455 94742 283464
rect 88616 283416 88668 283422
rect 88320 283364 88616 283370
rect 88320 283358 88668 283364
rect 88984 283416 89036 283422
rect 88984 283358 89036 283364
rect 88320 283342 88656 283358
rect 83556 283280 83608 283286
rect 70308 283222 70360 283228
rect 70950 283248 71006 283257
rect 70950 283183 71006 283192
rect 71962 283248 72018 283257
rect 71962 283183 72018 283192
rect 73250 283248 73306 283257
rect 73306 283206 73416 283234
rect 83352 283228 83556 283234
rect 83352 283222 83608 283228
rect 84016 283280 84068 283286
rect 84016 283222 84068 283228
rect 83352 283206 83596 283222
rect 73250 283183 73306 283192
rect 83476 283121 83504 283206
rect 88628 283121 88656 283342
rect 95344 283234 95372 286078
rect 95620 283506 95648 306346
rect 96620 304292 96672 304298
rect 96620 304234 96672 304240
rect 96632 283778 96660 304234
rect 96586 283750 96660 283778
rect 95620 283478 96048 283506
rect 96586 283492 96614 283750
rect 96724 283506 96752 327694
rect 97264 309868 97316 309874
rect 97264 309810 97316 309816
rect 97276 286142 97304 309810
rect 99196 308440 99248 308446
rect 99196 308382 99248 308388
rect 99208 292574 99236 308382
rect 99024 292546 99236 292574
rect 98368 291304 98420 291310
rect 98368 291246 98420 291252
rect 97264 286136 97316 286142
rect 97264 286078 97316 286084
rect 97906 284880 97962 284889
rect 97906 284815 97962 284824
rect 97920 283506 97948 284815
rect 98090 284472 98146 284481
rect 98090 284407 98146 284416
rect 96724 283478 97152 283506
rect 97704 283478 97948 283506
rect 98104 283422 98132 284407
rect 98380 283506 98408 291246
rect 98460 284436 98512 284442
rect 98460 284378 98512 284384
rect 98256 283478 98408 283506
rect 98092 283416 98144 283422
rect 98092 283358 98144 283364
rect 98368 283416 98420 283422
rect 98368 283358 98420 283364
rect 95344 283206 95496 283234
rect 83462 283112 83518 283121
rect 83462 283047 83518 283056
rect 88614 283112 88670 283121
rect 92386 283112 92442 283121
rect 92184 283070 92386 283098
rect 88614 283047 88670 283056
rect 92386 283047 92442 283056
rect 69664 283008 69716 283014
rect 95344 282985 95372 283206
rect 69664 282950 69716 282956
rect 95330 282976 95386 282985
rect 95330 282911 95386 282920
rect 69020 282736 69072 282742
rect 69018 282704 69020 282713
rect 69072 282704 69074 282713
rect 68848 282674 68968 282690
rect 68848 282668 68980 282674
rect 68848 282662 68928 282668
rect 69018 282639 69074 282648
rect 68928 282610 68980 282616
rect 68940 281217 68968 282610
rect 68926 281208 68982 281217
rect 68926 281143 68982 281152
rect 68940 280226 68968 281143
rect 68928 280220 68980 280226
rect 68928 280162 68980 280168
rect 98380 277394 98408 283358
rect 98472 282878 98500 284378
rect 99024 283506 99052 292546
rect 99300 292534 99328 370631
rect 99484 315314 99512 389146
rect 100404 387122 100432 390374
rect 100818 390130 100846 390388
rect 100772 390102 100846 390130
rect 101048 390374 101384 390402
rect 102120 390374 102272 390402
rect 100772 389298 100800 390102
rect 100760 389292 100812 389298
rect 100760 389234 100812 389240
rect 100772 388657 100800 389234
rect 100758 388648 100814 388657
rect 100758 388583 100814 388592
rect 100392 387116 100444 387122
rect 100392 387058 100444 387064
rect 101048 373994 101076 390374
rect 102140 387048 102192 387054
rect 102140 386990 102192 386996
rect 101954 385792 102010 385801
rect 101954 385727 102010 385736
rect 100772 373966 101076 373994
rect 100772 358086 100800 373966
rect 100760 358080 100812 358086
rect 100760 358022 100812 358028
rect 99472 315308 99524 315314
rect 99472 315250 99524 315256
rect 101402 304192 101458 304201
rect 101402 304127 101458 304136
rect 99288 292528 99340 292534
rect 99288 292470 99340 292476
rect 99300 291310 99328 292470
rect 99288 291304 99340 291310
rect 99288 291246 99340 291252
rect 100022 289912 100078 289921
rect 100022 289847 100078 289856
rect 99102 284608 99158 284617
rect 99102 284543 99158 284552
rect 98624 283478 99052 283506
rect 98918 283384 98974 283393
rect 98840 283342 98918 283370
rect 98460 282872 98512 282878
rect 98460 282814 98512 282820
rect 98380 277366 98776 277394
rect 98090 267880 98146 267889
rect 98090 267815 98146 267824
rect 98104 267734 98132 267815
rect 98012 267706 98132 267734
rect 98748 267714 98776 277366
rect 98840 269822 98868 283342
rect 98918 283319 98974 283328
rect 98918 282840 98974 282849
rect 98918 282775 98974 282784
rect 98932 282198 98960 282775
rect 98920 282192 98972 282198
rect 98920 282134 98972 282140
rect 99116 279585 99144 284543
rect 99380 284368 99432 284374
rect 99380 284310 99432 284316
rect 99102 279576 99158 279585
rect 99102 279511 99158 279520
rect 99392 278050 99420 284310
rect 99380 278044 99432 278050
rect 99380 277986 99432 277992
rect 99470 270464 99526 270473
rect 99470 270399 99526 270408
rect 98828 269816 98880 269822
rect 98828 269758 98880 269764
rect 99012 268048 99064 268054
rect 99010 268016 99012 268025
rect 99064 268016 99066 268025
rect 99010 267951 99066 267960
rect 98736 267708 98788 267714
rect 69018 244352 69074 244361
rect 69018 244287 69074 244296
rect 69032 242214 69060 244287
rect 69020 242208 69072 242214
rect 69020 242150 69072 242156
rect 95424 241800 95476 241806
rect 69846 241768 69902 241777
rect 70950 241768 71006 241777
rect 70840 241726 70950 241754
rect 69846 241703 69902 241712
rect 90362 241768 90418 241777
rect 70950 241703 71006 241712
rect 89824 241726 90362 241754
rect 68816 241590 68876 241618
rect 68848 241505 68876 241590
rect 69124 241590 69184 241618
rect 69400 241590 69736 241618
rect 68834 241496 68890 241505
rect 68834 241431 68890 241440
rect 68652 240644 68704 240650
rect 68652 240586 68704 240592
rect 68848 240145 68876 241431
rect 69020 240168 69072 240174
rect 68834 240136 68890 240145
rect 69020 240110 69072 240116
rect 68834 240071 68890 240080
rect 68560 237992 68612 237998
rect 68560 237934 68612 237940
rect 67914 236600 67970 236609
rect 67914 236535 67970 236544
rect 69032 193866 69060 240110
rect 69124 233238 69152 241590
rect 69400 240009 69428 241590
rect 69386 240000 69442 240009
rect 69386 239935 69442 239944
rect 69112 233232 69164 233238
rect 69112 233174 69164 233180
rect 69020 193860 69072 193866
rect 69020 193802 69072 193808
rect 69664 180872 69716 180878
rect 69664 180814 69716 180820
rect 67732 156664 67784 156670
rect 67732 156606 67784 156612
rect 68928 156664 68980 156670
rect 68928 156606 68980 156612
rect 67744 127673 67772 156606
rect 68940 156058 68968 156606
rect 68928 156052 68980 156058
rect 68928 155994 68980 156000
rect 69112 140888 69164 140894
rect 69112 140830 69164 140836
rect 68652 140072 68704 140078
rect 68652 140014 68704 140020
rect 67822 136096 67878 136105
rect 67822 136031 67878 136040
rect 67730 127664 67786 127673
rect 67730 127599 67786 127608
rect 67836 118425 67864 136031
rect 68560 134632 68612 134638
rect 68560 134574 68612 134580
rect 68572 128217 68600 134574
rect 68558 128208 68614 128217
rect 68558 128143 68614 128152
rect 67822 118416 67878 118425
rect 67822 118351 67878 118360
rect 68664 113174 68692 140014
rect 69124 134722 69152 140830
rect 69204 137284 69256 137290
rect 69204 137226 69256 137232
rect 69000 134694 69152 134722
rect 69216 134722 69244 137226
rect 69676 134745 69704 180814
rect 69756 151836 69808 151842
rect 69756 151778 69808 151784
rect 69662 134736 69718 134745
rect 69216 134694 69552 134722
rect 69662 134671 69718 134680
rect 69768 134638 69796 151778
rect 69860 142118 69888 241703
rect 82726 241632 82782 241641
rect 69952 241590 70288 241618
rect 71332 241590 71392 241618
rect 71884 241590 71944 241618
rect 72496 241590 72648 241618
rect 69952 240174 69980 241590
rect 71332 241505 71360 241590
rect 71318 241496 71374 241505
rect 71318 241431 71374 241440
rect 69940 240168 69992 240174
rect 69940 240110 69992 240116
rect 71332 240038 71360 241431
rect 70492 240032 70544 240038
rect 70492 239974 70544 239980
rect 71320 240032 71372 240038
rect 71320 239974 71372 239980
rect 70398 146432 70454 146441
rect 70398 146367 70454 146376
rect 69848 142112 69900 142118
rect 69848 142054 69900 142060
rect 69860 140894 69888 142054
rect 69848 140888 69900 140894
rect 69848 140830 69900 140836
rect 70214 138000 70270 138009
rect 70214 137935 70270 137944
rect 70228 134722 70256 137935
rect 70306 134872 70362 134881
rect 70306 134807 70308 134816
rect 70360 134807 70362 134816
rect 70308 134778 70360 134784
rect 70104 134694 70256 134722
rect 70412 134722 70440 146367
rect 70504 139641 70532 239974
rect 71780 239828 71832 239834
rect 71780 239770 71832 239776
rect 71792 218006 71820 239770
rect 71884 236706 71912 241590
rect 72620 239873 72648 241590
rect 72712 241590 73048 241618
rect 73264 241590 73600 241618
rect 73816 241590 74152 241618
rect 74644 241590 74704 241618
rect 74828 241590 75256 241618
rect 75472 241590 75808 241618
rect 76024 241590 76360 241618
rect 76484 241590 76912 241618
rect 77312 241590 77464 241618
rect 77588 241590 78016 241618
rect 78232 241590 78568 241618
rect 78784 241590 79120 241618
rect 79336 241590 79672 241618
rect 80224 241590 80652 241618
rect 80776 241590 80836 241618
rect 72606 239864 72662 239873
rect 72712 239834 72740 241590
rect 73160 240168 73212 240174
rect 73160 240110 73212 240116
rect 72606 239799 72662 239808
rect 72700 239828 72752 239834
rect 72700 239770 72752 239776
rect 71872 236700 71924 236706
rect 71872 236642 71924 236648
rect 71780 218000 71832 218006
rect 71780 217942 71832 217948
rect 73068 218000 73120 218006
rect 73068 217942 73120 217948
rect 72976 158840 73028 158846
rect 72976 158782 73028 158788
rect 72882 145072 72938 145081
rect 72882 145007 72938 145016
rect 72896 144974 72924 145007
rect 71780 144968 71832 144974
rect 71780 144910 71832 144916
rect 72884 144968 72936 144974
rect 72884 144910 72936 144916
rect 71410 141400 71466 141409
rect 71410 141335 71466 141344
rect 70490 139632 70546 139641
rect 70490 139567 70546 139576
rect 71320 139460 71372 139466
rect 71320 139402 71372 139408
rect 71332 134722 71360 139402
rect 70412 134694 70656 134722
rect 71024 134694 71360 134722
rect 71424 134722 71452 141335
rect 71792 134722 71820 144910
rect 72988 137970 73016 158782
rect 72976 137964 73028 137970
rect 72976 137906 73028 137912
rect 72330 137456 72386 137465
rect 72330 137391 72386 137400
rect 72344 134722 72372 137391
rect 73080 135153 73108 217942
rect 73172 138417 73200 240110
rect 73264 227633 73292 241590
rect 73816 240174 73844 241590
rect 74644 241233 74672 241590
rect 74630 241224 74686 241233
rect 74630 241159 74686 241168
rect 73804 240168 73856 240174
rect 73804 240110 73856 240116
rect 74540 240168 74592 240174
rect 74540 240110 74592 240116
rect 73802 240000 73858 240009
rect 73802 239935 73858 239944
rect 73250 227624 73306 227633
rect 73250 227559 73306 227568
rect 73436 185632 73488 185638
rect 73436 185574 73488 185580
rect 73158 138408 73214 138417
rect 73158 138343 73214 138352
rect 73160 137964 73212 137970
rect 73160 137906 73212 137912
rect 73066 135144 73122 135153
rect 73066 135079 73122 135088
rect 73172 134994 73200 137906
rect 73172 134966 73246 134994
rect 71424 134694 71576 134722
rect 71792 134694 72128 134722
rect 72344 134694 72680 134722
rect 73218 134708 73246 134966
rect 73448 134722 73476 185574
rect 73816 142361 73844 239935
rect 74552 229770 74580 240110
rect 74540 229764 74592 229770
rect 74540 229706 74592 229712
rect 74644 158030 74672 241159
rect 74828 238921 74856 241590
rect 75472 240174 75500 241590
rect 75460 240168 75512 240174
rect 75460 240110 75512 240116
rect 76024 240106 76052 241590
rect 76012 240100 76064 240106
rect 76012 240042 76064 240048
rect 75184 239692 75236 239698
rect 75184 239634 75236 239640
rect 74814 238912 74870 238921
rect 74814 238847 74870 238856
rect 74828 235929 74856 238847
rect 75196 238754 75224 239634
rect 76484 238754 76512 241590
rect 76656 240644 76708 240650
rect 76656 240586 76708 240592
rect 76564 240100 76616 240106
rect 76564 240042 76616 240048
rect 75012 238746 75224 238754
rect 75000 238740 75224 238746
rect 75052 238726 75224 238740
rect 75000 238682 75052 238688
rect 74814 235920 74870 235929
rect 74814 235855 74870 235864
rect 75196 163441 75224 238726
rect 76024 238726 76512 238754
rect 76024 238377 76052 238726
rect 76576 238649 76604 240042
rect 76562 238640 76618 238649
rect 76562 238575 76618 238584
rect 76010 238368 76066 238377
rect 76010 238303 76066 238312
rect 75920 167068 75972 167074
rect 75920 167010 75972 167016
rect 75182 163432 75238 163441
rect 75182 163367 75238 163376
rect 74722 162072 74778 162081
rect 74722 162007 74778 162016
rect 74632 158024 74684 158030
rect 74632 157966 74684 157972
rect 73802 142352 73858 142361
rect 73802 142287 73858 142296
rect 73816 139466 73844 142287
rect 73804 139460 73856 139466
rect 73804 139402 73856 139408
rect 74262 137320 74318 137329
rect 74262 137255 74318 137264
rect 74276 134722 74304 137255
rect 74736 134994 74764 162007
rect 75184 155984 75236 155990
rect 75184 155926 75236 155932
rect 75196 151814 75224 155926
rect 75196 151786 75408 151814
rect 74816 151156 74868 151162
rect 74816 151098 74868 151104
rect 73448 134694 73600 134722
rect 74152 134694 74304 134722
rect 74690 134966 74764 134994
rect 74690 134708 74718 134966
rect 74828 134722 74856 151098
rect 75380 134842 75408 151786
rect 75932 141522 75960 167010
rect 76576 158030 76604 238575
rect 76668 165753 76696 240586
rect 77312 239698 77340 241590
rect 77300 239692 77352 239698
rect 77300 239634 77352 239640
rect 76748 237992 76800 237998
rect 76748 237934 76800 237940
rect 76760 167686 76788 237934
rect 77588 233209 77616 241590
rect 78232 240106 78260 241590
rect 78680 240168 78732 240174
rect 78680 240110 78732 240116
rect 78220 240100 78272 240106
rect 78220 240042 78272 240048
rect 78588 237448 78640 237454
rect 78588 237390 78640 237396
rect 77942 236056 77998 236065
rect 77942 235991 77998 236000
rect 77574 233200 77630 233209
rect 77574 233135 77630 233144
rect 77300 204944 77352 204950
rect 77300 204886 77352 204892
rect 76748 167680 76800 167686
rect 76748 167622 76800 167628
rect 76760 167074 76788 167622
rect 76748 167068 76800 167074
rect 76748 167010 76800 167016
rect 76654 165744 76710 165753
rect 76654 165679 76710 165688
rect 76564 158024 76616 158030
rect 76564 157966 76616 157972
rect 76010 142488 76066 142497
rect 76010 142423 76066 142432
rect 76024 142118 76052 142423
rect 76012 142112 76064 142118
rect 76012 142054 76064 142060
rect 75932 141494 76328 141522
rect 76012 141432 76064 141438
rect 76012 141374 76064 141380
rect 75368 134836 75420 134842
rect 75368 134778 75420 134784
rect 75380 134722 75408 134778
rect 74828 134694 75256 134722
rect 75380 134694 75808 134722
rect 69756 134632 69808 134638
rect 69756 134574 69808 134580
rect 76024 134586 76052 141374
rect 76300 134722 76328 141494
rect 76668 136649 76696 165679
rect 76654 136640 76710 136649
rect 76654 136575 76710 136584
rect 77312 134994 77340 204886
rect 77956 142866 77984 235991
rect 78600 210458 78628 237390
rect 78692 230450 78720 240110
rect 78784 237454 78812 241590
rect 79336 240174 79364 241590
rect 79324 240168 79376 240174
rect 79324 240110 79376 240116
rect 79322 238776 79378 238785
rect 79322 238711 79378 238720
rect 78772 237448 78824 237454
rect 78772 237390 78824 237396
rect 78680 230444 78732 230450
rect 78680 230386 78732 230392
rect 78588 210452 78640 210458
rect 78588 210394 78640 210400
rect 77944 142860 77996 142866
rect 77944 142802 77996 142808
rect 78034 138680 78090 138689
rect 78034 138615 78090 138624
rect 77266 134966 77340 134994
rect 76300 134694 76728 134722
rect 77266 134708 77294 134966
rect 78048 134722 78076 138615
rect 78496 137964 78548 137970
rect 78496 137906 78548 137912
rect 78508 134722 78536 137906
rect 79336 137465 79364 238711
rect 80624 237289 80652 241590
rect 80808 238678 80836 241590
rect 80900 241590 81328 241618
rect 81820 241590 81880 241618
rect 82432 241590 82676 241618
rect 80796 238672 80848 238678
rect 80796 238614 80848 238620
rect 80610 237280 80666 237289
rect 80610 237215 80666 237224
rect 79414 236736 79470 236745
rect 79414 236671 79470 236680
rect 79428 139398 79456 236671
rect 80624 236065 80652 237215
rect 80610 236056 80666 236065
rect 80610 235991 80666 236000
rect 80900 235906 80928 241590
rect 81820 241369 81848 241590
rect 81806 241360 81862 241369
rect 81806 241295 81862 241304
rect 81820 240106 81848 241295
rect 80980 240100 81032 240106
rect 80980 240042 81032 240048
rect 81808 240100 81860 240106
rect 81808 240042 81860 240048
rect 80072 235878 80928 235906
rect 80072 231130 80100 235878
rect 80992 234614 81020 240042
rect 82648 239562 82676 241590
rect 82984 241590 83320 241618
rect 83536 241590 83688 241618
rect 82726 241567 82782 241576
rect 82636 239556 82688 239562
rect 82636 239498 82688 239504
rect 80716 234586 81020 234614
rect 80060 231124 80112 231130
rect 80060 231066 80112 231072
rect 79966 141536 80022 141545
rect 79966 141471 80022 141480
rect 79416 139392 79468 139398
rect 79416 139334 79468 139340
rect 79428 137970 79456 139334
rect 79416 137964 79468 137970
rect 79416 137906 79468 137912
rect 79322 137456 79378 137465
rect 79322 137391 79378 137400
rect 79046 136912 79102 136921
rect 79046 136847 79102 136856
rect 79060 134722 79088 136847
rect 79600 136672 79652 136678
rect 79600 136614 79652 136620
rect 79612 134722 79640 136614
rect 79980 134722 80008 141471
rect 80610 141400 80666 141409
rect 80610 141335 80666 141344
rect 80624 134722 80652 141335
rect 80716 140078 80744 234586
rect 82740 174554 82768 241567
rect 83292 235385 83320 241590
rect 83660 239494 83688 241590
rect 83752 241590 84088 241618
rect 84640 241590 84976 241618
rect 83648 239488 83700 239494
rect 83648 239430 83700 239436
rect 83278 235376 83334 235385
rect 83278 235311 83334 235320
rect 83752 234614 83780 241590
rect 84948 238814 84976 241590
rect 85040 241590 85192 241618
rect 85592 241590 85744 241618
rect 85868 241590 86296 241618
rect 86696 241590 86848 241618
rect 87064 241590 87400 241618
rect 87616 241590 87952 241618
rect 88352 241590 88504 241618
rect 89056 241590 89392 241618
rect 89608 241590 89668 241618
rect 84936 238808 84988 238814
rect 84936 238750 84988 238756
rect 85040 234614 85068 241590
rect 85592 240009 85620 241590
rect 85578 240000 85634 240009
rect 85578 239935 85634 239944
rect 85488 238808 85540 238814
rect 85592 238785 85620 239935
rect 85488 238750 85540 238756
rect 85578 238776 85634 238785
rect 82832 234586 83780 234614
rect 84212 234586 85068 234614
rect 82832 217977 82860 234586
rect 84212 227746 84240 234586
rect 85500 231810 85528 238750
rect 85578 238711 85634 238720
rect 85868 234614 85896 241590
rect 86696 240145 86724 241590
rect 86682 240136 86738 240145
rect 86682 240071 86738 240080
rect 86960 237176 87012 237182
rect 86960 237118 87012 237124
rect 85592 234586 85896 234614
rect 85488 231804 85540 231810
rect 85488 231746 85540 231752
rect 84120 227718 84240 227746
rect 85486 227760 85542 227769
rect 82818 217968 82874 217977
rect 82818 217903 82874 217912
rect 84120 206310 84148 227718
rect 85486 227695 85542 227704
rect 84108 206304 84160 206310
rect 84108 206246 84160 206252
rect 85500 177342 85528 227695
rect 85488 177336 85540 177342
rect 85488 177278 85540 177284
rect 85500 176730 85528 177278
rect 84200 176724 84252 176730
rect 84200 176666 84252 176672
rect 85488 176724 85540 176730
rect 85488 176666 85540 176672
rect 82084 174548 82136 174554
rect 82084 174490 82136 174496
rect 82728 174548 82780 174554
rect 82728 174490 82780 174496
rect 81438 152416 81494 152425
rect 81438 152351 81494 152360
rect 81452 151814 81480 152351
rect 81452 151786 82032 151814
rect 80704 140072 80756 140078
rect 80704 140014 80756 140020
rect 81898 136776 81954 136785
rect 81898 136711 81954 136720
rect 81348 136672 81400 136678
rect 81348 136614 81400 136620
rect 81070 136232 81126 136241
rect 81070 136167 81126 136176
rect 81084 134722 81112 136167
rect 81360 134858 81388 136614
rect 81912 134858 81940 136711
rect 77832 134694 78076 134722
rect 78200 134694 78536 134722
rect 78752 134694 79088 134722
rect 79304 134694 79640 134722
rect 79856 134694 80008 134722
rect 80408 134694 80652 134722
rect 80776 134694 81112 134722
rect 81314 134830 81388 134858
rect 81866 134830 81940 134858
rect 81314 134708 81342 134830
rect 81866 134708 81894 134830
rect 82004 134722 82032 151786
rect 82096 136921 82124 174490
rect 82912 165640 82964 165646
rect 82912 165582 82964 165588
rect 82176 164280 82228 164286
rect 82176 164222 82228 164228
rect 82082 136912 82138 136921
rect 82082 136847 82138 136856
rect 82188 136678 82216 164222
rect 82818 151872 82874 151881
rect 82818 151807 82874 151816
rect 82176 136672 82228 136678
rect 82176 136614 82228 136620
rect 82832 134994 82860 151807
rect 82786 134966 82860 134994
rect 82004 134694 82432 134722
rect 82786 134708 82814 134966
rect 82924 134722 82952 165582
rect 84212 151814 84240 176666
rect 85592 171902 85620 234586
rect 86972 207738 87000 237118
rect 87064 233170 87092 241590
rect 87616 237182 87644 241590
rect 87604 237176 87656 237182
rect 87604 237118 87656 237124
rect 88352 234598 88380 241590
rect 88432 239556 88484 239562
rect 88432 239498 88484 239504
rect 88444 239465 88472 239498
rect 88430 239456 88486 239465
rect 88430 239391 88486 239400
rect 89364 235958 89392 241590
rect 89640 239970 89668 241590
rect 89720 240168 89772 240174
rect 89720 240110 89772 240116
rect 89628 239964 89680 239970
rect 89628 239906 89680 239912
rect 89626 239456 89682 239465
rect 89626 239391 89682 239400
rect 89536 236020 89588 236026
rect 89536 235962 89588 235968
rect 89352 235952 89404 235958
rect 89352 235894 89404 235900
rect 88340 234592 88392 234598
rect 88340 234534 88392 234540
rect 87052 233164 87104 233170
rect 87052 233106 87104 233112
rect 88248 233164 88300 233170
rect 88248 233106 88300 233112
rect 88260 229770 88288 233106
rect 87604 229764 87656 229770
rect 87604 229706 87656 229712
rect 88248 229764 88300 229770
rect 88248 229706 88300 229712
rect 86960 207732 87012 207738
rect 86960 207674 87012 207680
rect 86314 175808 86370 175817
rect 86314 175743 86370 175752
rect 86328 175409 86356 175743
rect 86314 175400 86370 175409
rect 86314 175335 86370 175344
rect 86222 172544 86278 172553
rect 86222 172479 86278 172488
rect 85580 171896 85632 171902
rect 85580 171838 85632 171844
rect 84212 151786 84608 151814
rect 83462 142624 83518 142633
rect 83462 142559 83518 142568
rect 83476 134722 83504 142559
rect 84476 140072 84528 140078
rect 84476 140014 84528 140020
rect 84488 134994 84516 140014
rect 84442 134966 84516 134994
rect 82924 134694 83352 134722
rect 83476 134694 83904 134722
rect 84442 134708 84470 134966
rect 84580 134722 84608 151786
rect 85580 144764 85632 144770
rect 85580 144706 85632 144712
rect 85488 136672 85540 136678
rect 85488 136614 85540 136620
rect 85500 134722 85528 136614
rect 84580 134694 85008 134722
rect 85376 134694 85528 134722
rect 85592 134722 85620 144706
rect 86236 136678 86264 172479
rect 86328 151881 86356 175335
rect 87144 161492 87196 161498
rect 87144 161434 87196 161440
rect 86314 151872 86370 151881
rect 86314 151807 86370 151816
rect 86868 149728 86920 149734
rect 86868 149670 86920 149676
rect 86880 146266 86908 149670
rect 86868 146260 86920 146266
rect 86868 146202 86920 146208
rect 86314 145072 86370 145081
rect 86314 145007 86370 145016
rect 86328 140049 86356 145007
rect 86866 144800 86922 144809
rect 86866 144735 86922 144744
rect 86880 140185 86908 144735
rect 86866 140176 86922 140185
rect 86866 140111 86922 140120
rect 86314 140040 86370 140049
rect 86314 139975 86370 139984
rect 86224 136672 86276 136678
rect 86224 136614 86276 136620
rect 86880 134722 86908 140111
rect 87052 137964 87104 137970
rect 87052 137906 87104 137912
rect 87064 137601 87092 137906
rect 87050 137592 87106 137601
rect 87050 137527 87106 137536
rect 87064 136746 87092 137527
rect 87052 136740 87104 136746
rect 87052 136682 87104 136688
rect 87050 135960 87106 135969
rect 87050 135895 87106 135904
rect 87064 134858 87092 135895
rect 85592 134694 85928 134722
rect 86480 134694 86908 134722
rect 87018 134830 87092 134858
rect 87018 134708 87046 134830
rect 87156 134722 87184 161434
rect 87616 148345 87644 229706
rect 89548 182850 89576 235962
rect 89536 182844 89588 182850
rect 89536 182786 89588 182792
rect 88984 175976 89036 175982
rect 88984 175918 89036 175924
rect 88340 173936 88392 173942
rect 88340 173878 88392 173884
rect 87696 168496 87748 168502
rect 87696 168438 87748 168444
rect 87602 148336 87658 148345
rect 87602 148271 87658 148280
rect 87604 146260 87656 146266
rect 87604 146202 87656 146208
rect 87616 134858 87644 146202
rect 87708 137329 87736 168438
rect 87694 137320 87750 137329
rect 87694 137255 87750 137264
rect 87616 134830 87736 134858
rect 87708 134722 87736 134830
rect 88352 134722 88380 173878
rect 88616 154624 88668 154630
rect 88616 154566 88668 154572
rect 88524 142180 88576 142186
rect 88524 142122 88576 142128
rect 88628 142154 88656 154566
rect 88996 144770 89024 175918
rect 89640 146266 89668 239391
rect 89732 233170 89760 240110
rect 89824 236026 89852 241726
rect 95128 241748 95424 241754
rect 95128 241742 95476 241748
rect 95128 241726 95464 241742
rect 90362 241703 90418 241712
rect 90376 241590 90712 241618
rect 91264 241590 91324 241618
rect 90376 240174 90404 241590
rect 90364 240168 90416 240174
rect 90364 240110 90416 240116
rect 91008 239488 91060 239494
rect 91008 239430 91060 239436
rect 91020 238649 91048 239430
rect 91296 239358 91324 241590
rect 91388 241590 91816 241618
rect 92368 241590 92428 241618
rect 91284 239352 91336 239358
rect 91284 239294 91336 239300
rect 91388 238754 91416 241590
rect 92400 240825 92428 241590
rect 92584 241590 92920 241618
rect 92386 240816 92442 240825
rect 92386 240751 92442 240760
rect 91112 238726 91416 238754
rect 91006 238640 91062 238649
rect 91006 238575 91062 238584
rect 90362 236600 90418 236609
rect 90362 236535 90418 236544
rect 89812 236020 89864 236026
rect 89812 235962 89864 235968
rect 89720 233164 89772 233170
rect 89720 233106 89772 233112
rect 90376 195294 90404 236535
rect 90364 195288 90416 195294
rect 90364 195230 90416 195236
rect 91020 180130 91048 238575
rect 91112 238513 91140 238726
rect 91098 238504 91154 238513
rect 91098 238439 91154 238448
rect 91112 237425 91140 238439
rect 91098 237416 91154 237425
rect 91098 237351 91154 237360
rect 92294 236736 92350 236745
rect 92294 236671 92350 236680
rect 91008 180124 91060 180130
rect 91008 180066 91060 180072
rect 91008 171828 91060 171834
rect 91008 171770 91060 171776
rect 89718 167104 89774 167113
rect 89718 167039 89774 167048
rect 89628 146260 89680 146266
rect 89628 146202 89680 146208
rect 88984 144764 89036 144770
rect 88984 144706 89036 144712
rect 88628 142126 89208 142154
rect 88536 138009 88564 142122
rect 89076 140140 89128 140146
rect 89076 140082 89128 140088
rect 88522 138000 88578 138009
rect 88522 137935 88578 137944
rect 89088 134994 89116 140082
rect 89042 134966 89116 134994
rect 87156 134694 87584 134722
rect 87708 134694 87952 134722
rect 88352 134694 88504 134722
rect 89042 134708 89070 134966
rect 89180 134722 89208 142126
rect 89732 134722 89760 167039
rect 90088 144764 90140 144770
rect 90088 144706 90140 144712
rect 90100 134722 90128 144706
rect 91020 136882 91048 171770
rect 92308 160138 92336 236671
rect 92386 236600 92442 236609
rect 92386 236535 92442 236544
rect 91744 160132 91796 160138
rect 91744 160074 91796 160080
rect 92296 160132 92348 160138
rect 92296 160074 92348 160080
rect 91756 151814 91784 160074
rect 92400 158778 92428 236535
rect 92584 218754 92612 241590
rect 93458 241466 93486 241604
rect 94024 241590 94084 241618
rect 93446 241460 93498 241466
rect 93446 241402 93498 241408
rect 93458 241346 93486 241402
rect 93458 241318 93532 241346
rect 93504 240145 93532 241318
rect 94056 240854 94084 241590
rect 94148 241590 94576 241618
rect 95680 241590 95740 241618
rect 94044 240848 94096 240854
rect 94044 240790 94096 240796
rect 93490 240136 93546 240145
rect 94148 240122 94176 241590
rect 93490 240071 93546 240080
rect 93872 240094 94176 240122
rect 93872 238066 93900 240094
rect 95712 240009 95740 241590
rect 95804 241590 96232 241618
rect 96784 241590 97120 241618
rect 95698 240000 95754 240009
rect 95698 239935 95754 239944
rect 93952 239352 94004 239358
rect 93952 239294 94004 239300
rect 93860 238060 93912 238066
rect 93860 238002 93912 238008
rect 93964 236706 93992 239294
rect 95804 238754 95832 241590
rect 97092 240145 97120 241590
rect 97184 241590 97336 241618
rect 97552 241590 97888 241618
rect 97078 240136 97134 240145
rect 97078 240071 97134 240080
rect 95882 240000 95938 240009
rect 97184 239986 97212 241590
rect 95882 239935 95938 239944
rect 96632 239958 97212 239986
rect 95252 238726 95832 238754
rect 93952 236700 94004 236706
rect 93952 236642 94004 236648
rect 92572 218748 92624 218754
rect 92572 218690 92624 218696
rect 95252 213246 95280 238726
rect 95240 213240 95292 213246
rect 95240 213182 95292 213188
rect 93674 176760 93730 176769
rect 93124 176724 93176 176730
rect 93674 176695 93676 176704
rect 93124 176666 93176 176672
rect 93728 176695 93730 176704
rect 93676 176666 93728 176672
rect 92664 168428 92716 168434
rect 92664 168370 92716 168376
rect 92480 162920 92532 162926
rect 92480 162862 92532 162868
rect 91836 158772 91888 158778
rect 91836 158714 91888 158720
rect 92388 158772 92440 158778
rect 92388 158714 92440 158720
rect 91296 151786 91784 151814
rect 91100 140820 91152 140826
rect 91100 140762 91152 140768
rect 91112 137290 91140 140762
rect 91100 137284 91152 137290
rect 91100 137226 91152 137232
rect 91008 136876 91060 136882
rect 91008 136818 91060 136824
rect 91192 136604 91244 136610
rect 91192 136546 91244 136552
rect 91204 135318 91232 136546
rect 91296 135386 91324 151786
rect 91848 142154 91876 158714
rect 91756 142126 91876 142154
rect 91756 136610 91784 142126
rect 91836 136876 91888 136882
rect 91836 136818 91888 136824
rect 91744 136604 91796 136610
rect 91744 136546 91796 136552
rect 91284 135380 91336 135386
rect 91284 135322 91336 135328
rect 91192 135312 91244 135318
rect 91192 135254 91244 135260
rect 89180 134694 89608 134722
rect 89732 134694 89976 134722
rect 90100 134694 90528 134722
rect 91204 134586 91232 135254
rect 91296 134722 91324 135322
rect 91848 134722 91876 136818
rect 92492 134994 92520 162862
rect 92492 134966 92566 134994
rect 91296 134694 91632 134722
rect 91848 134694 92184 134722
rect 92538 134708 92566 134966
rect 92676 134722 92704 168370
rect 92754 157448 92810 157457
rect 92754 157383 92810 157392
rect 92768 142154 92796 157383
rect 93136 144770 93164 176666
rect 93860 153944 93912 153950
rect 93860 153886 93912 153892
rect 93124 144764 93176 144770
rect 93124 144706 93176 144712
rect 92768 142126 93256 142154
rect 93228 134722 93256 142126
rect 93766 138272 93822 138281
rect 93766 138207 93822 138216
rect 92676 134694 93104 134722
rect 93228 134694 93656 134722
rect 93780 134638 93808 138207
rect 93872 138106 93900 153886
rect 95424 146940 95476 146946
rect 95424 146882 95476 146888
rect 95240 146260 95292 146266
rect 95240 146202 95292 146208
rect 93950 145616 94006 145625
rect 93950 145551 94006 145560
rect 93860 138100 93912 138106
rect 93860 138042 93912 138048
rect 93964 134722 93992 145551
rect 94686 138136 94742 138145
rect 94320 138100 94372 138106
rect 94686 138071 94742 138080
rect 94320 138042 94372 138048
rect 94332 134722 94360 138042
rect 93964 134694 94208 134722
rect 94332 134694 94576 134722
rect 76024 134558 76176 134586
rect 91080 134558 91232 134586
rect 93768 134632 93820 134638
rect 93768 134574 93820 134580
rect 94700 131889 94728 138071
rect 95146 136776 95202 136785
rect 95146 136711 95202 136720
rect 95160 133890 95188 136711
rect 95148 133884 95200 133890
rect 95148 133826 95200 133832
rect 94686 131880 94742 131889
rect 94686 131815 94742 131824
rect 67468 113146 67588 113174
rect 67652 113146 68140 113174
rect 68664 113146 68968 113174
rect 67454 100192 67510 100201
rect 67454 100127 67510 100136
rect 67362 98016 67418 98025
rect 67284 97974 67362 98002
rect 66812 95192 66864 95198
rect 66812 95134 66864 95140
rect 66824 95033 66852 95134
rect 66810 95024 66866 95033
rect 66810 94959 66866 94968
rect 67180 93832 67232 93838
rect 67180 93774 67232 93780
rect 67192 93401 67220 93774
rect 67178 93392 67234 93401
rect 67178 93327 67234 93336
rect 67284 89622 67312 97974
rect 67362 97951 67418 97960
rect 67362 97200 67418 97209
rect 67362 97135 67418 97144
rect 67376 92478 67404 97135
rect 67468 93922 67496 100127
rect 67560 97209 67588 113146
rect 67546 97200 67602 97209
rect 67546 97135 67602 97144
rect 67546 95840 67602 95849
rect 67546 95775 67602 95784
rect 67560 94058 67588 95775
rect 67560 94030 67772 94058
rect 67468 93894 67588 93922
rect 67456 93832 67508 93838
rect 67456 93774 67508 93780
rect 67364 92472 67416 92478
rect 67364 92414 67416 92420
rect 67272 89616 67324 89622
rect 67272 89558 67324 89564
rect 67468 88330 67496 93774
rect 67456 88324 67508 88330
rect 67456 88266 67508 88272
rect 66166 78568 66222 78577
rect 66166 78503 66222 78512
rect 65524 77240 65576 77246
rect 65524 77182 65576 77188
rect 64788 73160 64840 73166
rect 64788 73102 64840 73108
rect 67560 70378 67588 93894
rect 67744 93838 67772 94030
rect 68112 93854 68140 113146
rect 67732 93832 67784 93838
rect 68112 93826 68416 93854
rect 67732 93774 67784 93780
rect 68388 92834 68416 93826
rect 68388 92806 68816 92834
rect 68388 84194 68416 92806
rect 68558 92712 68614 92721
rect 68558 92647 68614 92656
rect 68572 86737 68600 92647
rect 68940 88262 68968 113146
rect 94778 98560 94834 98569
rect 94778 98495 94834 98504
rect 69018 92576 69074 92585
rect 69170 92562 69198 92820
rect 69722 92585 69750 92820
rect 70274 92698 70302 92820
rect 70274 92670 70348 92698
rect 69708 92576 69764 92585
rect 69170 92534 69244 92562
rect 69018 92511 69074 92520
rect 68928 88256 68980 88262
rect 68928 88198 68980 88204
rect 68558 86728 68614 86737
rect 68558 86663 68614 86672
rect 67744 84166 68416 84194
rect 69032 84194 69060 92511
rect 69032 84166 69152 84194
rect 67640 75200 67692 75206
rect 67640 75142 67692 75148
rect 67548 70372 67600 70378
rect 67548 70314 67600 70320
rect 65524 66904 65576 66910
rect 65524 66846 65576 66852
rect 61752 32428 61804 32434
rect 61752 32370 61804 32376
rect 63500 17264 63552 17270
rect 63500 17206 63552 17212
rect 63512 16574 63540 17206
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 59372 16546 59676 16574
rect 60752 16546 60872 16574
rect 63512 16546 64368 16574
rect 52472 6886 52592 6914
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 51368 480 51396 3402
rect 52564 480 52592 6886
rect 53300 490 53328 16546
rect 53576 598 53788 626
rect 53576 490 53604 598
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 462 53604 490
rect 53760 480 53788 598
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 56796 490 56824 16546
rect 58440 10328 58492 10334
rect 58440 10270 58492 10276
rect 57072 598 57284 626
rect 57072 490 57100 598
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 462 57100 490
rect 57256 480 57284 598
rect 58452 480 58480 10270
rect 59648 480 59676 16546
rect 60844 480 60872 16546
rect 61568 13116 61620 13122
rect 61568 13058 61620 13064
rect 61580 490 61608 13058
rect 63224 4140 63276 4146
rect 63224 4082 63276 4088
rect 61856 598 62068 626
rect 61856 490 61884 598
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 462 61884 490
rect 62040 480 62068 598
rect 63236 480 63264 4082
rect 64340 480 64368 16546
rect 65536 6914 65564 66846
rect 66258 55856 66314 55865
rect 66258 55791 66314 55800
rect 66272 16574 66300 55791
rect 67652 16574 67680 75142
rect 67744 63510 67772 84166
rect 69018 82104 69074 82113
rect 69018 82039 69074 82048
rect 67732 63504 67784 63510
rect 67732 63446 67784 63452
rect 66272 16546 66760 16574
rect 67652 16546 67956 16574
rect 65444 6886 65564 6914
rect 65444 4146 65472 6886
rect 65524 4820 65576 4826
rect 65524 4762 65576 4768
rect 65432 4140 65484 4146
rect 65432 4082 65484 4088
rect 65536 480 65564 4762
rect 66732 480 66760 16546
rect 67928 480 67956 16546
rect 69032 3534 69060 82039
rect 69124 60722 69152 84166
rect 69216 81326 69244 92534
rect 69708 92511 69764 92520
rect 70320 91050 70348 92670
rect 70826 92562 70854 92820
rect 71194 92721 71222 92820
rect 71180 92712 71236 92721
rect 71746 92698 71774 92820
rect 71746 92670 71820 92698
rect 71180 92647 71236 92656
rect 70504 92534 70854 92562
rect 70308 91044 70360 91050
rect 70308 90986 70360 90992
rect 70320 89758 70348 90986
rect 70308 89752 70360 89758
rect 70308 89694 70360 89700
rect 69204 81320 69256 81326
rect 69204 81262 69256 81268
rect 70398 73808 70454 73817
rect 70398 73743 70454 73752
rect 69112 60716 69164 60722
rect 69112 60658 69164 60664
rect 69112 25560 69164 25566
rect 69112 25502 69164 25508
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 69124 480 69152 25502
rect 70412 16574 70440 73743
rect 70504 59294 70532 92534
rect 71792 88233 71820 92670
rect 72298 92562 72326 92820
rect 72850 92721 72878 92820
rect 72836 92712 72892 92721
rect 73402 92698 73430 92820
rect 73770 92698 73798 92820
rect 72836 92647 72892 92656
rect 73356 92670 73430 92698
rect 73724 92670 73798 92698
rect 74322 92698 74350 92820
rect 74874 92698 74902 92820
rect 74322 92670 74396 92698
rect 71884 92534 72326 92562
rect 71778 88224 71834 88233
rect 71778 88159 71834 88168
rect 71884 66230 71912 92534
rect 73356 92449 73384 92670
rect 73342 92440 73398 92449
rect 73342 92375 73398 92384
rect 73724 92313 73752 92670
rect 73710 92304 73766 92313
rect 73710 92239 73766 92248
rect 74368 90953 74396 92670
rect 74828 92670 74902 92698
rect 74828 92177 74856 92670
rect 75426 92562 75454 92820
rect 75794 92562 75822 92820
rect 76346 92698 76374 92820
rect 76346 92670 76420 92698
rect 74920 92534 75454 92562
rect 75564 92534 75822 92562
rect 74814 92168 74870 92177
rect 74814 92103 74870 92112
rect 74354 90944 74410 90953
rect 74354 90879 74410 90888
rect 73804 89752 73856 89758
rect 73804 89694 73856 89700
rect 72606 88224 72662 88233
rect 72606 88159 72662 88168
rect 72620 86873 72648 88159
rect 72606 86864 72662 86873
rect 72606 86799 72662 86808
rect 71872 66224 71924 66230
rect 71872 66166 71924 66172
rect 73816 61946 73844 89694
rect 74920 88482 74948 92534
rect 74552 88454 74948 88482
rect 74552 84114 74580 88454
rect 75564 84194 75592 92534
rect 76392 86601 76420 92670
rect 76898 92562 76926 92820
rect 77450 92562 77478 92820
rect 76576 92534 76926 92562
rect 77312 92534 77478 92562
rect 78002 92562 78030 92820
rect 78370 92562 78398 92820
rect 78922 92562 78950 92820
rect 79474 92562 79502 92820
rect 78002 92534 78076 92562
rect 78370 92534 78444 92562
rect 78922 92534 78996 92562
rect 76378 86592 76434 86601
rect 76378 86527 76434 86536
rect 76576 84194 76604 92534
rect 74644 84166 75592 84194
rect 75932 84166 76604 84194
rect 74540 84108 74592 84114
rect 74540 84050 74592 84056
rect 74538 72448 74594 72457
rect 74538 72383 74594 72392
rect 73804 61940 73856 61946
rect 73804 61882 73856 61888
rect 70492 59288 70544 59294
rect 70492 59230 70544 59236
rect 71780 54528 71832 54534
rect 71780 54470 71832 54476
rect 71792 16574 71820 54470
rect 73160 36576 73212 36582
rect 73160 36518 73212 36524
rect 73172 16574 73200 36518
rect 74552 16574 74580 72383
rect 74644 56574 74672 84166
rect 75932 82754 75960 84166
rect 77312 82822 77340 92534
rect 78048 88097 78076 92534
rect 78034 88088 78090 88097
rect 78034 88023 78090 88032
rect 78416 85542 78444 92534
rect 78968 91050 78996 92534
rect 79428 92534 79502 92562
rect 80026 92562 80054 92820
rect 80578 92562 80606 92820
rect 80946 92562 80974 92820
rect 80026 92534 80100 92562
rect 80578 92534 80652 92562
rect 79428 92410 79456 92534
rect 79416 92404 79468 92410
rect 79416 92346 79468 92352
rect 78956 91044 79008 91050
rect 78956 90986 79008 90992
rect 78404 85536 78456 85542
rect 78404 85478 78456 85484
rect 77300 82816 77352 82822
rect 77300 82758 77352 82764
rect 75920 82748 75972 82754
rect 75920 82690 75972 82696
rect 79322 79384 79378 79393
rect 79322 79319 79378 79328
rect 74632 56568 74684 56574
rect 74632 56510 74684 56516
rect 78680 46232 78732 46238
rect 78680 46174 78732 46180
rect 75920 42084 75972 42090
rect 75920 42026 75972 42032
rect 75932 16574 75960 42026
rect 77300 18624 77352 18630
rect 77300 18566 77352 18572
rect 77312 16574 77340 18566
rect 78692 16574 78720 46174
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 75932 16546 76236 16574
rect 77312 16546 78168 16574
rect 78692 16546 79272 16574
rect 70308 3528 70360 3534
rect 70308 3470 70360 3476
rect 70320 480 70348 3470
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 73356 490 73384 16546
rect 73632 598 73844 626
rect 73632 490 73660 598
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 462 73660 490
rect 73816 480 73844 598
rect 75012 480 75040 16546
rect 75184 11756 75236 11762
rect 75184 11698 75236 11704
rect 75196 3466 75224 11698
rect 75184 3460 75236 3466
rect 75184 3402 75236 3408
rect 76208 480 76236 16546
rect 77392 3528 77444 3534
rect 77392 3470 77444 3476
rect 77404 480 77432 3470
rect 78140 490 78168 16546
rect 78416 598 78628 626
rect 78416 490 78444 598
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 462 78444 490
rect 78600 480 78628 598
rect 79244 490 79272 16546
rect 79336 3534 79364 79319
rect 80072 64802 80100 92534
rect 80624 92410 80652 92534
rect 80716 92534 80974 92562
rect 81498 92562 81526 92820
rect 82050 92562 82078 92820
rect 82602 92562 82630 92820
rect 82970 92698 82998 92820
rect 82970 92670 83044 92698
rect 81498 92534 81572 92562
rect 82050 92534 82124 92562
rect 82602 92534 82676 92562
rect 80612 92404 80664 92410
rect 80612 92346 80664 92352
rect 80716 88262 80744 92534
rect 81544 89457 81572 92534
rect 81530 89448 81586 89457
rect 81530 89383 81586 89392
rect 80704 88256 80756 88262
rect 82096 88233 82124 92534
rect 82648 91225 82676 92534
rect 82634 91216 82690 91225
rect 82634 91151 82690 91160
rect 83016 89729 83044 92670
rect 83522 92562 83550 92820
rect 83292 92534 83550 92562
rect 84074 92562 84102 92820
rect 84626 92698 84654 92820
rect 84626 92670 84700 92698
rect 84074 92534 84148 92562
rect 83002 89720 83058 89729
rect 83002 89655 83058 89664
rect 80704 88198 80756 88204
rect 82082 88224 82138 88233
rect 80716 76566 80744 88198
rect 82082 88159 82138 88168
rect 83292 84194 83320 92534
rect 83462 91216 83518 91225
rect 83462 91151 83518 91160
rect 82832 84166 83320 84194
rect 82832 78674 82860 84166
rect 82820 78668 82872 78674
rect 82820 78610 82872 78616
rect 80704 76560 80756 76566
rect 80704 76502 80756 76508
rect 80060 64796 80112 64802
rect 80060 64738 80112 64744
rect 83476 60654 83504 91151
rect 84120 87961 84148 92534
rect 84672 89593 84700 92670
rect 85178 92562 85206 92820
rect 85546 92562 85574 92820
rect 86098 92698 86126 92820
rect 86098 92670 86172 92698
rect 85178 92534 85252 92562
rect 85546 92534 85712 92562
rect 85224 89758 85252 92534
rect 85212 89752 85264 89758
rect 85212 89694 85264 89700
rect 84658 89584 84714 89593
rect 84658 89519 84714 89528
rect 84842 89584 84898 89593
rect 84842 89519 84898 89528
rect 84106 87952 84162 87961
rect 84106 87887 84162 87896
rect 83464 60648 83516 60654
rect 83464 60590 83516 60596
rect 84856 59362 84884 89519
rect 85580 77988 85632 77994
rect 85580 77930 85632 77936
rect 84844 59356 84896 59362
rect 84844 59298 84896 59304
rect 84200 38004 84252 38010
rect 84200 37946 84252 37952
rect 82820 35216 82872 35222
rect 82820 35158 82872 35164
rect 81440 24132 81492 24138
rect 81440 24074 81492 24080
rect 81452 16574 81480 24074
rect 82832 16574 82860 35158
rect 84212 16574 84240 37946
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 84212 16546 84516 16574
rect 79324 3528 79376 3534
rect 79324 3470 79376 3476
rect 80888 3460 80940 3466
rect 80888 3402 80940 3408
rect 79520 598 79732 626
rect 79520 490 79548 598
rect 78558 -960 78670 480
rect 79244 462 79548 490
rect 79704 480 79732 598
rect 80900 480 80928 3402
rect 81636 490 81664 16546
rect 81912 598 82124 626
rect 81912 490 81940 598
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 462 81940 490
rect 82096 480 82124 598
rect 83292 480 83320 16546
rect 84488 480 84516 16546
rect 85592 3534 85620 77930
rect 85684 74526 85712 92534
rect 86144 88262 86172 92670
rect 86650 92562 86678 92820
rect 87202 92698 87230 92820
rect 87202 92670 87276 92698
rect 86328 92534 86678 92562
rect 86132 88256 86184 88262
rect 86132 88198 86184 88204
rect 86328 84194 86356 92534
rect 87248 89593 87276 92670
rect 87570 92562 87598 92820
rect 88122 92562 88150 92820
rect 88674 92750 88702 92820
rect 88662 92744 88714 92750
rect 88662 92686 88714 92692
rect 89226 92562 89254 92820
rect 87340 92534 87598 92562
rect 87800 92534 88150 92562
rect 88352 92534 89254 92562
rect 89778 92562 89806 92820
rect 90146 92682 90174 92820
rect 90134 92676 90186 92682
rect 90134 92618 90186 92624
rect 90698 92562 90726 92820
rect 91008 92676 91060 92682
rect 91008 92618 91060 92624
rect 89778 92534 89852 92562
rect 87234 89584 87290 89593
rect 87234 89519 87290 89528
rect 87340 88482 87368 92534
rect 85776 84166 86356 84194
rect 86972 88454 87368 88482
rect 85776 81394 85804 84166
rect 85764 81388 85816 81394
rect 85764 81330 85816 81336
rect 85672 74520 85724 74526
rect 85672 74462 85724 74468
rect 86972 62014 87000 88454
rect 87800 84194 87828 92534
rect 87064 84166 87828 84194
rect 88352 84182 88380 92534
rect 89824 86970 89852 92534
rect 89916 92534 90726 92562
rect 89812 86964 89864 86970
rect 89812 86906 89864 86912
rect 88340 84176 88392 84182
rect 87064 64870 87092 84166
rect 88340 84118 88392 84124
rect 89916 82793 89944 92534
rect 91020 92449 91048 92618
rect 91250 92562 91278 92820
rect 91802 92698 91830 92820
rect 91802 92670 91876 92698
rect 91250 92534 91324 92562
rect 91006 92440 91062 92449
rect 91006 92375 91062 92384
rect 90362 83464 90418 83473
rect 90362 83399 90418 83408
rect 89902 82784 89958 82793
rect 89902 82719 89958 82728
rect 88340 68332 88392 68338
rect 88340 68274 88392 68280
rect 87052 64864 87104 64870
rect 87052 64806 87104 64812
rect 86960 62008 87012 62014
rect 86960 61950 87012 61956
rect 86960 53100 87012 53106
rect 86960 53042 87012 53048
rect 85670 26888 85726 26897
rect 85670 26823 85726 26832
rect 85580 3528 85632 3534
rect 85580 3470 85632 3476
rect 85684 480 85712 26823
rect 86972 16574 87000 53042
rect 88352 16574 88380 68274
rect 89720 21412 89772 21418
rect 89720 21354 89772 21360
rect 89732 16574 89760 21354
rect 90376 20670 90404 83399
rect 91020 57934 91048 92375
rect 91296 85377 91324 92534
rect 91848 92449 91876 92670
rect 92354 92562 92382 92820
rect 92722 92562 92750 92820
rect 93274 92562 93302 92820
rect 93826 92614 93854 92820
rect 94392 92806 94728 92834
rect 93814 92608 93866 92614
rect 92354 92534 92428 92562
rect 92722 92534 92796 92562
rect 93274 92534 93348 92562
rect 93814 92550 93866 92556
rect 94504 92608 94556 92614
rect 94504 92550 94556 92556
rect 91834 92440 91890 92449
rect 91834 92375 91890 92384
rect 92400 92041 92428 92534
rect 92768 92313 92796 92534
rect 92754 92304 92810 92313
rect 92754 92239 92810 92248
rect 92386 92032 92442 92041
rect 92386 91967 92442 91976
rect 93124 89752 93176 89758
rect 93124 89694 93176 89700
rect 91282 85368 91338 85377
rect 91282 85303 91338 85312
rect 93136 71738 93164 89694
rect 93320 86902 93348 92534
rect 93308 86896 93360 86902
rect 93308 86838 93360 86844
rect 93124 71732 93176 71738
rect 93124 71674 93176 71680
rect 92478 71088 92534 71097
rect 92478 71023 92534 71032
rect 91008 57928 91060 57934
rect 91008 57870 91060 57876
rect 90364 20664 90416 20670
rect 90364 20606 90416 20612
rect 92492 16574 92520 71023
rect 93858 68232 93914 68241
rect 93858 68167 93914 68176
rect 93872 16574 93900 68167
rect 94516 67561 94544 92550
rect 94700 92546 94728 92806
rect 94688 92540 94740 92546
rect 94688 92482 94740 92488
rect 94792 89978 94820 98495
rect 94872 94512 94924 94518
rect 94872 94454 94924 94460
rect 94884 92682 94912 94454
rect 94872 92676 94924 92682
rect 94872 92618 94924 92624
rect 94700 89950 94820 89978
rect 94700 89622 94728 89950
rect 94778 89856 94834 89865
rect 94778 89791 94834 89800
rect 94688 89616 94740 89622
rect 94688 89558 94740 89564
rect 94792 82754 94820 89791
rect 95252 89457 95280 146202
rect 95436 127673 95464 146882
rect 95422 127664 95478 127673
rect 95422 127599 95478 127608
rect 95330 120320 95386 120329
rect 95330 120255 95386 120264
rect 95238 89448 95294 89457
rect 95238 89383 95294 89392
rect 94780 82748 94832 82754
rect 94780 82690 94832 82696
rect 95148 82748 95200 82754
rect 95148 82690 95200 82696
rect 95160 77217 95188 82690
rect 95146 77208 95202 77217
rect 95146 77143 95202 77152
rect 95344 71670 95372 120255
rect 95896 92614 95924 239935
rect 96632 206378 96660 239958
rect 97552 238754 97580 241590
rect 96908 238726 97580 238754
rect 96908 234666 96936 238726
rect 96896 234660 96948 234666
rect 96896 234602 96948 234608
rect 97356 234660 97408 234666
rect 97356 234602 97408 234608
rect 97908 234660 97960 234666
rect 97908 234602 97960 234608
rect 97264 233912 97316 233918
rect 97264 233854 97316 233860
rect 96620 206372 96672 206378
rect 96620 206314 96672 206320
rect 95974 139496 96030 139505
rect 95974 139431 96030 139440
rect 95988 126449 96016 139431
rect 96618 130928 96674 130937
rect 96618 130863 96674 130872
rect 95974 126440 96030 126449
rect 95974 126375 96030 126384
rect 96068 120352 96120 120358
rect 96066 120320 96068 120329
rect 96120 120320 96122 120329
rect 96066 120255 96122 120264
rect 95976 94580 96028 94586
rect 95976 94522 96028 94528
rect 95884 92608 95936 92614
rect 95884 92550 95936 92556
rect 95988 86601 96016 94522
rect 95974 86592 96030 86601
rect 95974 86527 96030 86536
rect 96632 83473 96660 130863
rect 97172 126268 97224 126274
rect 97172 126210 97224 126216
rect 97184 123321 97212 126210
rect 97170 123312 97226 123321
rect 97170 123247 97226 123256
rect 97080 121372 97132 121378
rect 97080 121314 97132 121320
rect 97092 120873 97120 121314
rect 97078 120864 97134 120873
rect 97078 120799 97134 120808
rect 97276 114073 97304 233854
rect 97368 209166 97396 234602
rect 97356 209160 97408 209166
rect 97356 209102 97408 209108
rect 97920 160750 97948 234602
rect 97908 160744 97960 160750
rect 97908 160686 97960 160692
rect 97920 160206 97948 160686
rect 97356 160200 97408 160206
rect 97356 160142 97408 160148
rect 97908 160200 97960 160206
rect 97908 160142 97960 160148
rect 97368 122505 97396 160142
rect 98012 157418 98040 267706
rect 98736 267650 98788 267656
rect 99288 262200 99340 262206
rect 99288 262142 99340 262148
rect 99300 261497 99328 262142
rect 99286 261488 99342 261497
rect 99286 261423 99342 261432
rect 98090 260944 98146 260953
rect 98090 260879 98146 260888
rect 98104 233918 98132 260879
rect 98642 258496 98698 258505
rect 98642 258431 98698 258440
rect 98552 243568 98604 243574
rect 98552 243510 98604 243516
rect 98182 242584 98238 242593
rect 98182 242519 98238 242528
rect 98196 242214 98224 242519
rect 98564 242298 98592 243510
rect 98440 242270 98592 242298
rect 98184 242208 98236 242214
rect 98184 242150 98236 242156
rect 98564 240038 98592 242270
rect 98552 240032 98604 240038
rect 98552 239974 98604 239980
rect 98092 233912 98144 233918
rect 98092 233854 98144 233860
rect 98092 202836 98144 202842
rect 98092 202778 98144 202784
rect 98104 202230 98132 202778
rect 98092 202224 98144 202230
rect 98092 202166 98144 202172
rect 98000 157412 98052 157418
rect 98000 157354 98052 157360
rect 97448 146328 97500 146334
rect 97448 146270 97500 146276
rect 97460 129062 97488 146270
rect 97538 144800 97594 144809
rect 97538 144735 97594 144744
rect 97552 131481 97580 144735
rect 97908 135244 97960 135250
rect 97908 135186 97960 135192
rect 97920 133929 97948 135186
rect 97906 133920 97962 133929
rect 97906 133855 97962 133864
rect 97908 132456 97960 132462
rect 97908 132398 97960 132404
rect 97920 132297 97948 132398
rect 97906 132288 97962 132297
rect 97906 132223 97962 132232
rect 97538 131472 97594 131481
rect 97538 131407 97594 131416
rect 97722 130928 97778 130937
rect 97722 130863 97778 130872
rect 97540 130620 97592 130626
rect 97540 130562 97592 130568
rect 97552 130121 97580 130562
rect 97736 130422 97764 130863
rect 97724 130416 97776 130422
rect 97724 130358 97776 130364
rect 97538 130112 97594 130121
rect 97538 130047 97594 130056
rect 97908 129736 97960 129742
rect 97908 129678 97960 129684
rect 97448 129056 97500 129062
rect 97448 128998 97500 129004
rect 97920 128489 97948 129678
rect 97906 128480 97962 128489
rect 97906 128415 97962 128424
rect 97632 128308 97684 128314
rect 97632 128250 97684 128256
rect 97644 127129 97672 128250
rect 97630 127120 97686 127129
rect 97630 127055 97686 127064
rect 97908 126880 97960 126886
rect 97908 126822 97960 126828
rect 97920 126313 97948 126822
rect 97906 126304 97962 126313
rect 97906 126239 97962 126248
rect 97908 125588 97960 125594
rect 97908 125530 97960 125536
rect 97814 125488 97870 125497
rect 97814 125423 97870 125432
rect 97828 124846 97856 125423
rect 97816 124840 97868 124846
rect 97816 124782 97868 124788
rect 97920 124681 97948 125530
rect 97906 124672 97962 124681
rect 97906 124607 97962 124616
rect 97908 124160 97960 124166
rect 97906 124128 97908 124137
rect 97960 124128 97962 124137
rect 97906 124063 97962 124072
rect 97908 122800 97960 122806
rect 97908 122742 97960 122748
rect 97354 122496 97410 122505
rect 97354 122431 97410 122440
rect 97920 121689 97948 122742
rect 97906 121680 97962 121689
rect 97906 121615 97962 121624
rect 97908 120080 97960 120086
rect 97908 120022 97960 120028
rect 97920 119513 97948 120022
rect 97906 119504 97962 119513
rect 97906 119439 97962 119448
rect 97906 118688 97962 118697
rect 97906 118623 97908 118632
rect 97960 118623 97962 118632
rect 97908 118594 97960 118600
rect 97356 117292 97408 117298
rect 97356 117234 97408 117240
rect 97368 116521 97396 117234
rect 97908 117224 97960 117230
rect 97908 117166 97960 117172
rect 97920 117065 97948 117166
rect 97906 117056 97962 117065
rect 97906 116991 97962 117000
rect 97354 116512 97410 116521
rect 97354 116447 97410 116456
rect 97816 115932 97868 115938
rect 97816 115874 97868 115880
rect 97828 114889 97856 115874
rect 97906 115696 97962 115705
rect 97906 115631 97962 115640
rect 97814 114880 97870 114889
rect 97814 114815 97870 114824
rect 97920 114578 97948 115631
rect 97908 114572 97960 114578
rect 97908 114514 97960 114520
rect 97262 114064 97318 114073
rect 97262 113999 97318 114008
rect 96712 111920 96764 111926
rect 96710 111888 96712 111897
rect 96764 111888 96766 111897
rect 96710 111823 96766 111832
rect 96804 111172 96856 111178
rect 96804 111114 96856 111120
rect 96816 111081 96844 111114
rect 96802 111072 96858 111081
rect 96802 111007 96858 111016
rect 96712 97028 96764 97034
rect 96712 96970 96764 96976
rect 96724 96665 96752 96970
rect 96710 96656 96766 96665
rect 96710 96591 96766 96600
rect 96618 83464 96674 83473
rect 96618 83399 96674 83408
rect 95332 71664 95384 71670
rect 95332 71606 95384 71612
rect 97276 67590 97304 113999
rect 97538 113520 97594 113529
rect 97538 113455 97594 113464
rect 97552 113218 97580 113455
rect 97540 113212 97592 113218
rect 97540 113154 97592 113160
rect 97906 112704 97962 112713
rect 97906 112639 97962 112648
rect 97354 111888 97410 111897
rect 97920 111858 97948 112639
rect 97354 111823 97410 111832
rect 97908 111852 97960 111858
rect 97368 92857 97396 111823
rect 97908 111794 97960 111800
rect 97816 110424 97868 110430
rect 97816 110366 97868 110372
rect 97828 110265 97856 110366
rect 97908 110356 97960 110362
rect 97908 110298 97960 110304
rect 97814 110256 97870 110265
rect 97814 110191 97870 110200
rect 97920 109721 97948 110298
rect 97906 109712 97962 109721
rect 97906 109647 97962 109656
rect 97908 108316 97960 108322
rect 97908 108258 97960 108264
rect 97920 108089 97948 108258
rect 97906 108080 97962 108089
rect 97906 108015 97962 108024
rect 97908 107636 97960 107642
rect 97908 107578 97960 107584
rect 97920 107273 97948 107578
rect 97906 107264 97962 107273
rect 97906 107199 97962 107208
rect 97906 106720 97962 106729
rect 97906 106655 97962 106664
rect 97920 106554 97948 106655
rect 97908 106548 97960 106554
rect 97908 106490 97960 106496
rect 97906 104272 97962 104281
rect 97906 104207 97908 104216
rect 97960 104207 97962 104216
rect 97908 104178 97960 104184
rect 98104 103514 98132 202166
rect 98656 111926 98684 258431
rect 99378 249248 99434 249257
rect 99378 249183 99434 249192
rect 98736 216640 98788 216646
rect 98736 216582 98788 216588
rect 98644 111920 98696 111926
rect 98644 111862 98696 111868
rect 98642 103592 98698 103601
rect 98642 103527 98698 103536
rect 97908 103488 97960 103494
rect 97906 103456 97908 103465
rect 98012 103486 98132 103514
rect 97960 103456 97962 103465
rect 97906 103391 97962 103400
rect 97908 103080 97960 103086
rect 97908 103022 97960 103028
rect 97920 102921 97948 103022
rect 97906 102912 97962 102921
rect 97906 102847 97962 102856
rect 97908 102128 97960 102134
rect 97906 102096 97908 102105
rect 97960 102096 97962 102105
rect 97906 102031 97962 102040
rect 97906 101280 97962 101289
rect 98012 101266 98040 103486
rect 97962 101238 98040 101266
rect 97906 101215 97962 101224
rect 97538 100464 97594 100473
rect 97538 100399 97594 100408
rect 97552 99414 97580 100399
rect 97908 100020 97960 100026
rect 97908 99962 97960 99968
rect 97920 99657 97948 99962
rect 97906 99648 97962 99657
rect 97906 99583 97962 99592
rect 97540 99408 97592 99414
rect 97540 99350 97592 99356
rect 97540 98660 97592 98666
rect 97540 98602 97592 98608
rect 97552 94489 97580 98602
rect 97906 98288 97962 98297
rect 97906 98223 97962 98232
rect 97920 98054 97948 98223
rect 97908 98048 97960 98054
rect 97908 97990 97960 97996
rect 97906 95296 97962 95305
rect 97906 95231 97908 95240
rect 97960 95231 97962 95240
rect 97908 95202 97960 95208
rect 97538 94480 97594 94489
rect 97538 94415 97594 94424
rect 97908 93832 97960 93838
rect 97908 93774 97960 93780
rect 97920 93673 97948 93774
rect 97906 93664 97962 93673
rect 97906 93599 97962 93608
rect 97354 92848 97410 92857
rect 97354 92783 97410 92792
rect 97264 67584 97316 67590
rect 94502 67552 94558 67561
rect 97264 67526 97316 67532
rect 94502 67487 94558 67496
rect 97276 64874 97304 67526
rect 97276 64846 97396 64874
rect 97264 51740 97316 51746
rect 97264 51682 97316 51688
rect 95240 19984 95292 19990
rect 95240 19926 95292 19932
rect 95252 16574 95280 19926
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 92492 16546 92796 16574
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 86868 3528 86920 3534
rect 86868 3470 86920 3476
rect 86880 480 86908 3470
rect 87524 490 87552 16546
rect 87800 598 88012 626
rect 87800 490 87828 598
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 462 87828 490
rect 87984 480 88012 598
rect 89180 480 89208 16546
rect 89916 490 89944 16546
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 90192 598 90404 626
rect 90192 490 90220 598
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 462 90220 490
rect 90376 480 90404 598
rect 91572 480 91600 3470
rect 92768 480 92796 16546
rect 93124 14476 93176 14482
rect 93124 14418 93176 14424
rect 93136 3466 93164 14418
rect 93124 3460 93176 3466
rect 93124 3402 93176 3408
rect 93952 2100 94004 2106
rect 93952 2042 94004 2048
rect 93964 480 93992 2042
rect 94700 490 94728 16546
rect 94976 598 95188 626
rect 94976 490 95004 598
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 462 95004 490
rect 95160 480 95188 598
rect 95804 490 95832 16546
rect 97276 7614 97304 51682
rect 97368 50386 97396 64846
rect 97356 50380 97408 50386
rect 97356 50322 97408 50328
rect 98182 15872 98238 15881
rect 98182 15807 98238 15816
rect 97448 7676 97500 7682
rect 97448 7618 97500 7624
rect 97264 7608 97316 7614
rect 97264 7550 97316 7556
rect 96080 598 96292 626
rect 96080 490 96108 598
rect 95118 -960 95230 480
rect 95804 462 96108 490
rect 96264 480 96292 598
rect 97460 480 97488 7618
rect 98196 490 98224 15807
rect 98656 3534 98684 103527
rect 98748 97034 98776 216582
rect 98826 214568 98882 214577
rect 98826 214503 98882 214512
rect 98840 202842 98868 214503
rect 98828 202836 98880 202842
rect 98828 202778 98880 202784
rect 98828 157412 98880 157418
rect 98828 157354 98880 157360
rect 98840 120358 98868 157354
rect 98828 120352 98880 120358
rect 98828 120294 98880 120300
rect 98828 108384 98880 108390
rect 98828 108326 98880 108332
rect 98736 97028 98788 97034
rect 98736 96970 98788 96976
rect 98840 87961 98868 108326
rect 99392 103086 99420 249183
rect 99484 234666 99512 270399
rect 100036 268394 100064 289847
rect 100206 283112 100262 283121
rect 100206 283047 100262 283056
rect 100220 277370 100248 283047
rect 100758 281888 100814 281897
rect 100758 281823 100814 281832
rect 100772 281586 100800 281823
rect 100760 281580 100812 281586
rect 100760 281522 100812 281528
rect 100852 281512 100904 281518
rect 100852 281454 100904 281460
rect 100864 280265 100892 281454
rect 100850 280256 100906 280265
rect 100850 280191 100906 280200
rect 100760 280152 100812 280158
rect 100760 280094 100812 280100
rect 100772 279449 100800 280094
rect 100758 279440 100814 279449
rect 100758 279375 100814 279384
rect 101416 278633 101444 304127
rect 101494 282704 101550 282713
rect 101494 282639 101550 282648
rect 101402 278624 101458 278633
rect 101402 278559 101458 278568
rect 100208 277364 100260 277370
rect 100208 277306 100260 277312
rect 100758 276176 100814 276185
rect 100758 276111 100814 276120
rect 100772 276078 100800 276111
rect 100760 276072 100812 276078
rect 100760 276014 100812 276020
rect 100758 275360 100814 275369
rect 100758 275295 100814 275304
rect 100944 275324 100996 275330
rect 100772 274718 100800 275295
rect 100944 275266 100996 275272
rect 100760 274712 100812 274718
rect 100760 274654 100812 274660
rect 100852 274644 100904 274650
rect 100852 274586 100904 274592
rect 100864 273737 100892 274586
rect 100956 274553 100984 275266
rect 100942 274544 100998 274553
rect 100942 274479 100998 274488
rect 100850 273728 100906 273737
rect 100850 273663 100906 273672
rect 100852 273216 100904 273222
rect 100852 273158 100904 273164
rect 100758 272912 100814 272921
rect 100758 272847 100814 272856
rect 100772 272542 100800 272847
rect 100760 272536 100812 272542
rect 100760 272478 100812 272484
rect 100864 272105 100892 273158
rect 101508 272513 101536 282639
rect 101968 277001 101996 385727
rect 102048 381608 102100 381614
rect 102048 381550 102100 381556
rect 101954 276992 102010 277001
rect 101954 276927 102010 276936
rect 101494 272504 101550 272513
rect 101494 272439 101550 272448
rect 100850 272096 100906 272105
rect 100850 272031 100906 272040
rect 101218 271280 101274 271289
rect 100760 271244 100812 271250
rect 101218 271215 101274 271224
rect 100760 271186 100812 271192
rect 100772 270473 100800 271186
rect 101232 271182 101260 271215
rect 102060 271182 102088 381550
rect 102152 354686 102180 386990
rect 102244 355978 102272 390374
rect 102520 390374 102856 390402
rect 102520 387054 102548 390374
rect 102508 387048 102560 387054
rect 102508 386990 102560 386996
rect 104162 385656 104218 385665
rect 104162 385591 104218 385600
rect 103426 382936 103482 382945
rect 103426 382871 103482 382880
rect 102232 355972 102284 355978
rect 102232 355914 102284 355920
rect 103336 355972 103388 355978
rect 103336 355914 103388 355920
rect 102140 354680 102192 354686
rect 102140 354622 102192 354628
rect 102138 287192 102194 287201
rect 102138 287127 102194 287136
rect 101220 271176 101272 271182
rect 101220 271118 101272 271124
rect 102048 271176 102100 271182
rect 102048 271118 102100 271124
rect 100758 270464 100814 270473
rect 100758 270399 100814 270408
rect 100760 269136 100812 269142
rect 100760 269078 100812 269084
rect 100772 268841 100800 269078
rect 100758 268832 100814 268841
rect 100758 268767 100814 268776
rect 100024 268388 100076 268394
rect 100024 268330 100076 268336
rect 100758 267200 100814 267209
rect 100758 267135 100814 267144
rect 100772 267102 100800 267135
rect 100760 267096 100812 267102
rect 100760 267038 100812 267044
rect 100758 266384 100814 266393
rect 100758 266319 100814 266328
rect 100772 265674 100800 266319
rect 100760 265668 100812 265674
rect 100760 265610 100812 265616
rect 100942 264752 100998 264761
rect 100942 264687 100998 264696
rect 100758 263936 100814 263945
rect 100758 263871 100814 263880
rect 100772 263634 100800 263871
rect 100760 263628 100812 263634
rect 100760 263570 100812 263576
rect 100668 263560 100720 263566
rect 100668 263502 100720 263508
rect 100680 262313 100708 263502
rect 100666 262304 100722 262313
rect 100666 262239 100722 262248
rect 100574 258088 100630 258097
rect 100574 258023 100630 258032
rect 99472 234660 99524 234666
rect 99472 234602 99524 234608
rect 100588 146334 100616 258023
rect 100024 146328 100076 146334
rect 100024 146270 100076 146276
rect 100576 146328 100628 146334
rect 100576 146270 100628 146276
rect 99472 117360 99524 117366
rect 99472 117302 99524 117308
rect 99484 115938 99512 117302
rect 99472 115932 99524 115938
rect 99472 115874 99524 115880
rect 100036 111178 100064 146270
rect 100680 117366 100708 262239
rect 100850 260672 100906 260681
rect 100850 260607 100906 260616
rect 100758 259856 100814 259865
rect 100758 259791 100814 259800
rect 100772 259554 100800 259791
rect 100760 259548 100812 259554
rect 100760 259490 100812 259496
rect 100864 259486 100892 260607
rect 100956 260137 100984 264687
rect 100942 260128 100998 260137
rect 100942 260063 100998 260072
rect 100852 259480 100904 259486
rect 100852 259422 100904 259428
rect 100758 259040 100814 259049
rect 100758 258975 100814 258984
rect 100772 258738 100800 258975
rect 100760 258732 100812 258738
rect 100760 258674 100812 258680
rect 101678 258224 101734 258233
rect 101678 258159 101734 258168
rect 101692 258058 101720 258159
rect 101680 258052 101732 258058
rect 101680 257994 101732 258000
rect 102046 257408 102102 257417
rect 102046 257343 102048 257352
rect 102100 257343 102102 257352
rect 102048 257314 102100 257320
rect 100758 256592 100814 256601
rect 100758 256527 100814 256536
rect 100772 255338 100800 256527
rect 100852 256012 100904 256018
rect 100852 255954 100904 255960
rect 100864 255785 100892 255954
rect 100850 255776 100906 255785
rect 100850 255711 100906 255720
rect 100760 255332 100812 255338
rect 100760 255274 100812 255280
rect 100758 254144 100814 254153
rect 100758 254079 100814 254088
rect 100772 254046 100800 254079
rect 100760 254040 100812 254046
rect 100760 253982 100812 253988
rect 100758 250880 100814 250889
rect 100758 250815 100814 250824
rect 100772 250510 100800 250815
rect 100760 250504 100812 250510
rect 100760 250446 100812 250452
rect 100864 250322 100892 255711
rect 101588 252544 101640 252550
rect 100942 252512 100998 252521
rect 101588 252486 101640 252492
rect 100942 252447 100998 252456
rect 100956 251161 100984 252447
rect 100942 251152 100998 251161
rect 100942 251087 100998 251096
rect 100772 250294 100892 250322
rect 100772 237425 100800 250294
rect 101494 250064 101550 250073
rect 101494 249999 101550 250008
rect 100852 249076 100904 249082
rect 100852 249018 100904 249024
rect 100864 248441 100892 249018
rect 100850 248432 100906 248441
rect 100850 248367 100906 248376
rect 101036 246356 101088 246362
rect 101036 246298 101088 246304
rect 101404 246356 101456 246362
rect 101404 246298 101456 246304
rect 101048 245993 101076 246298
rect 101034 245984 101090 245993
rect 101034 245919 101090 245928
rect 100944 245608 100996 245614
rect 100944 245550 100996 245556
rect 100852 245200 100904 245206
rect 100850 245168 100852 245177
rect 100904 245168 100906 245177
rect 100850 245103 100906 245112
rect 100956 244361 100984 245550
rect 100942 244352 100998 244361
rect 100942 244287 100998 244296
rect 100850 243536 100906 243545
rect 100850 243471 100852 243480
rect 100904 243471 100906 243480
rect 100852 243442 100904 243448
rect 100850 242720 100906 242729
rect 100850 242655 100906 242664
rect 100864 242282 100892 242655
rect 100852 242276 100904 242282
rect 100852 242218 100904 242224
rect 100758 237416 100814 237425
rect 100758 237351 100814 237360
rect 100760 124840 100812 124846
rect 100758 124808 100760 124817
rect 100812 124808 100814 124817
rect 100758 124743 100814 124752
rect 100668 117360 100720 117366
rect 100668 117302 100720 117308
rect 100024 111172 100076 111178
rect 100024 111114 100076 111120
rect 100116 111104 100168 111110
rect 100116 111046 100168 111052
rect 99380 103080 99432 103086
rect 99380 103022 99432 103028
rect 99392 102814 99420 103022
rect 99380 102808 99432 102814
rect 99380 102750 99432 102756
rect 100022 102232 100078 102241
rect 100022 102167 100078 102176
rect 98918 99104 98974 99113
rect 98918 99039 98974 99048
rect 98826 87952 98882 87961
rect 98826 87887 98882 87896
rect 98932 84153 98960 99039
rect 99012 96688 99064 96694
rect 99012 96630 99064 96636
rect 99024 92410 99052 96630
rect 99012 92404 99064 92410
rect 99012 92346 99064 92352
rect 100036 88330 100064 102167
rect 100128 89690 100156 111046
rect 101312 104848 101364 104854
rect 101312 104790 101364 104796
rect 101324 103494 101352 104790
rect 101312 103488 101364 103494
rect 101312 103430 101364 103436
rect 101416 100026 101444 246298
rect 101508 104854 101536 249999
rect 101600 246809 101628 252486
rect 101586 246800 101642 246809
rect 101586 246735 101642 246744
rect 101586 148336 101642 148345
rect 101586 148271 101642 148280
rect 101600 124234 101628 148271
rect 101588 124228 101640 124234
rect 101588 124170 101640 124176
rect 101496 104848 101548 104854
rect 101496 104790 101548 104796
rect 101404 100020 101456 100026
rect 101404 99962 101456 99968
rect 101404 97300 101456 97306
rect 101404 97242 101456 97248
rect 100116 89684 100168 89690
rect 100116 89626 100168 89632
rect 100024 88324 100076 88330
rect 100024 88266 100076 88272
rect 101416 85241 101444 97242
rect 101402 85232 101458 85241
rect 101402 85167 101458 85176
rect 98918 84144 98974 84153
rect 101600 84114 101628 124170
rect 102060 111926 102088 257314
rect 102152 152425 102180 287127
rect 103348 253978 103376 355914
rect 103440 281518 103468 382871
rect 103428 281512 103480 281518
rect 103428 281454 103480 281460
rect 102968 253972 103020 253978
rect 102968 253914 103020 253920
rect 103336 253972 103388 253978
rect 103336 253914 103388 253920
rect 102876 253224 102928 253230
rect 102876 253166 102928 253172
rect 102784 243500 102836 243506
rect 102784 243442 102836 243448
rect 102796 220794 102824 243442
rect 102888 241505 102916 253166
rect 102980 241806 103008 253914
rect 103612 242276 103664 242282
rect 103612 242218 103664 242224
rect 102968 241800 103020 241806
rect 102968 241742 103020 241748
rect 102874 241496 102930 241505
rect 102874 241431 102930 241440
rect 103520 229764 103572 229770
rect 103520 229706 103572 229712
rect 102784 220788 102836 220794
rect 102784 220730 102836 220736
rect 102138 152416 102194 152425
rect 102138 152351 102194 152360
rect 102874 151872 102930 151881
rect 102874 151807 102930 151816
rect 102782 147928 102838 147937
rect 102782 147863 102838 147872
rect 102140 144220 102192 144226
rect 102140 144162 102192 144168
rect 102048 111920 102100 111926
rect 102048 111862 102100 111868
rect 102060 110430 102088 111862
rect 102048 110424 102100 110430
rect 102048 110366 102100 110372
rect 101680 106548 101732 106554
rect 101680 106490 101732 106496
rect 101692 93129 101720 106490
rect 101678 93120 101734 93129
rect 101678 93055 101734 93064
rect 98918 84079 98974 84088
rect 101588 84108 101640 84114
rect 101588 84050 101640 84056
rect 100024 76560 100076 76566
rect 100024 76502 100076 76508
rect 100036 66162 100064 76502
rect 100024 66156 100076 66162
rect 100024 66098 100076 66104
rect 100760 50380 100812 50386
rect 100760 50322 100812 50328
rect 100772 16574 100800 50322
rect 100772 16546 101076 16574
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99840 3460 99892 3466
rect 99840 3402 99892 3408
rect 98472 598 98684 626
rect 98472 490 98500 598
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 462 98500 490
rect 98656 480 98684 598
rect 99852 480 99880 3402
rect 101048 480 101076 16546
rect 102152 3534 102180 144162
rect 102230 124808 102286 124817
rect 102230 124743 102286 124752
rect 102244 77246 102272 124743
rect 102796 117881 102824 147863
rect 102888 130626 102916 151807
rect 102876 130620 102928 130626
rect 102876 130562 102928 130568
rect 102782 117872 102838 117881
rect 102782 117807 102838 117816
rect 102322 93256 102378 93265
rect 102322 93191 102378 93200
rect 102336 86737 102364 93191
rect 103532 88330 103560 229706
rect 103624 216646 103652 242218
rect 104176 233209 104204 385591
rect 104544 383654 104572 390918
rect 105910 390960 105966 390969
rect 105322 390918 105768 390946
rect 105266 390895 105322 390904
rect 104866 390130 104894 390388
rect 104866 390102 104940 390130
rect 104544 383626 104848 383654
rect 104820 370569 104848 383626
rect 104912 378826 104940 390102
rect 105740 389065 105768 390918
rect 111982 390960 112038 390969
rect 107292 390934 107344 390940
rect 105910 390895 105966 390904
rect 105726 389056 105782 389065
rect 105726 388991 105782 389000
rect 105924 383654 105952 390895
rect 107304 390402 107332 390934
rect 111872 390918 111982 390946
rect 112732 390930 112760 391274
rect 112902 391096 112958 391105
rect 112902 391031 112958 391040
rect 111982 390895 112038 390904
rect 112720 390924 112772 390930
rect 112720 390866 112772 390872
rect 112916 390833 112944 391031
rect 112902 390824 112958 390833
rect 112902 390759 112958 390768
rect 106338 390130 106366 390388
rect 106292 390102 106366 390130
rect 106752 390374 107088 390402
rect 107304 390374 107792 390402
rect 106094 389056 106150 389065
rect 106094 388991 106150 389000
rect 105924 383626 106044 383654
rect 104900 378820 104952 378826
rect 104900 378762 104952 378768
rect 104806 370560 104862 370569
rect 104806 370495 104862 370504
rect 104256 320884 104308 320890
rect 104256 320826 104308 320832
rect 104268 268054 104296 320826
rect 104440 313336 104492 313342
rect 104440 313278 104492 313284
rect 104348 312656 104400 312662
rect 104348 312598 104400 312604
rect 104256 268048 104308 268054
rect 104256 267990 104308 267996
rect 104360 262206 104388 312598
rect 104452 305658 104480 313278
rect 104440 305652 104492 305658
rect 104440 305594 104492 305600
rect 105542 302424 105598 302433
rect 105542 302359 105598 302368
rect 104438 285832 104494 285841
rect 104438 285767 104494 285776
rect 104452 264246 104480 285767
rect 104440 264240 104492 264246
rect 104440 264182 104492 264188
rect 104348 262200 104400 262206
rect 104348 262142 104400 262148
rect 104808 261996 104860 262002
rect 104808 261938 104860 261944
rect 104254 253328 104310 253337
rect 104254 253263 104310 253272
rect 104162 233200 104218 233209
rect 104162 233135 104218 233144
rect 104268 223553 104296 253263
rect 104820 252550 104848 261938
rect 104808 252544 104860 252550
rect 104808 252486 104860 252492
rect 105556 240009 105584 302359
rect 106016 278769 106044 383626
rect 106108 382265 106136 388991
rect 106094 382256 106150 382265
rect 106094 382191 106150 382200
rect 106094 378720 106150 378729
rect 106094 378655 106150 378664
rect 106002 278760 106058 278769
rect 106002 278695 106058 278704
rect 106108 267102 106136 378655
rect 106186 320648 106242 320657
rect 106186 320583 106242 320592
rect 106200 320210 106228 320583
rect 106188 320204 106240 320210
rect 106188 320146 106240 320152
rect 106096 267096 106148 267102
rect 106096 267038 106148 267044
rect 106108 266393 106136 267038
rect 106188 266416 106240 266422
rect 106094 266384 106150 266393
rect 106188 266358 106240 266364
rect 106094 266319 106150 266328
rect 105636 264988 105688 264994
rect 105636 264930 105688 264936
rect 105648 245206 105676 264930
rect 106096 251184 106148 251190
rect 106096 251126 106148 251132
rect 106108 250510 106136 251126
rect 106096 250504 106148 250510
rect 106096 250446 106148 250452
rect 105636 245200 105688 245206
rect 105636 245142 105688 245148
rect 105634 241904 105690 241913
rect 105634 241839 105690 241848
rect 105542 240000 105598 240009
rect 105542 239935 105598 239944
rect 104254 223544 104310 223553
rect 104254 223479 104310 223488
rect 103612 216640 103664 216646
rect 103612 216582 103664 216588
rect 105648 214606 105676 241839
rect 106108 217326 106136 250446
rect 106200 249082 106228 266358
rect 106188 249076 106240 249082
rect 106188 249018 106240 249024
rect 106292 243574 106320 390102
rect 106752 389337 106780 390374
rect 106738 389328 106794 389337
rect 106738 389263 106794 389272
rect 107764 386306 107792 390374
rect 107856 390374 108376 390402
rect 107752 386300 107804 386306
rect 107752 386242 107804 386248
rect 107856 373994 107884 390374
rect 109098 390130 109126 390388
rect 109512 390374 109848 390402
rect 110400 390374 110736 390402
rect 109098 390102 109172 390130
rect 108302 389872 108358 389881
rect 108302 389807 108358 389816
rect 107672 373966 107884 373994
rect 107568 373380 107620 373386
rect 107568 373322 107620 373328
rect 107580 348362 107608 373322
rect 107672 372609 107700 373966
rect 107658 372600 107714 372609
rect 107658 372535 107714 372544
rect 106924 348356 106976 348362
rect 106924 348298 106976 348304
rect 107568 348356 107620 348362
rect 107568 348298 107620 348304
rect 106370 276992 106426 277001
rect 106370 276927 106426 276936
rect 106280 243568 106332 243574
rect 106280 243510 106332 243516
rect 106096 217320 106148 217326
rect 106096 217262 106148 217268
rect 105636 214600 105688 214606
rect 105636 214542 105688 214548
rect 103612 207732 103664 207738
rect 103612 207674 103664 207680
rect 104808 207732 104860 207738
rect 104808 207674 104860 207680
rect 103520 88324 103572 88330
rect 103520 88266 103572 88272
rect 102322 86728 102378 86737
rect 102322 86663 102378 86672
rect 103624 81394 103652 207674
rect 104820 207058 104848 207674
rect 104808 207052 104860 207058
rect 104808 206994 104860 207000
rect 104990 204368 105046 204377
rect 104990 204303 105046 204312
rect 104164 147688 104216 147694
rect 104164 147630 104216 147636
rect 103704 133204 103756 133210
rect 103704 133146 103756 133152
rect 103716 126886 103744 133146
rect 103704 126880 103756 126886
rect 103704 126822 103756 126828
rect 104176 119406 104204 147630
rect 104900 131164 104952 131170
rect 104900 131106 104952 131112
rect 104164 119400 104216 119406
rect 104164 119342 104216 119348
rect 104164 101448 104216 101454
rect 104164 101390 104216 101396
rect 104176 92546 104204 101390
rect 104164 92540 104216 92546
rect 104164 92482 104216 92488
rect 103612 81388 103664 81394
rect 103612 81330 103664 81336
rect 102232 77240 102284 77246
rect 102232 77182 102284 77188
rect 104912 16574 104940 131106
rect 105004 111897 105032 204303
rect 106280 171896 106332 171902
rect 106280 171838 106332 171844
rect 105542 162888 105598 162897
rect 105542 162823 105598 162832
rect 105556 132569 105584 162823
rect 105542 132560 105598 132569
rect 105542 132495 105598 132504
rect 105542 129024 105598 129033
rect 105542 128959 105598 128968
rect 104990 111888 105046 111897
rect 104990 111823 105046 111832
rect 105556 77994 105584 128959
rect 106188 105596 106240 105602
rect 106188 105538 106240 105544
rect 106200 104242 106228 105538
rect 106188 104236 106240 104242
rect 106188 104178 106240 104184
rect 105544 77988 105596 77994
rect 105544 77930 105596 77936
rect 106292 71777 106320 171838
rect 106384 129742 106412 276927
rect 106936 251190 106964 348298
rect 108212 312588 108264 312594
rect 108212 312530 108264 312536
rect 108224 309874 108252 312530
rect 108212 309868 108264 309874
rect 108212 309810 108264 309816
rect 107566 287736 107622 287745
rect 107566 287671 107622 287680
rect 107580 281518 107608 287671
rect 107568 281512 107620 281518
rect 107568 281454 107620 281460
rect 107016 280220 107068 280226
rect 107016 280162 107068 280168
rect 107028 273222 107056 280162
rect 107016 273216 107068 273222
rect 107016 273158 107068 273164
rect 108316 269385 108344 389807
rect 108396 388476 108448 388482
rect 108396 388418 108448 388424
rect 108408 380769 108436 388418
rect 109040 387048 109092 387054
rect 109040 386990 109092 386996
rect 108394 380760 108450 380769
rect 108394 380695 108450 380704
rect 108408 379545 108436 380695
rect 108394 379536 108450 379545
rect 108394 379471 108450 379480
rect 108946 379536 109002 379545
rect 108946 379471 109002 379480
rect 108856 376032 108908 376038
rect 108856 375974 108908 375980
rect 108868 352578 108896 375974
rect 108856 352572 108908 352578
rect 108856 352514 108908 352520
rect 108868 351966 108896 352514
rect 108396 351960 108448 351966
rect 108396 351902 108448 351908
rect 108856 351960 108908 351966
rect 108856 351902 108908 351908
rect 108302 269376 108358 269385
rect 108302 269311 108358 269320
rect 108408 254425 108436 351902
rect 108488 281580 108540 281586
rect 108488 281522 108540 281528
rect 108394 254416 108450 254425
rect 108394 254351 108450 254360
rect 106924 251184 106976 251190
rect 106924 251126 106976 251132
rect 106924 243568 106976 243574
rect 106924 243510 106976 243516
rect 106936 218822 106964 243510
rect 108302 238096 108358 238105
rect 108302 238031 108358 238040
rect 106924 218816 106976 218822
rect 106924 218758 106976 218764
rect 106924 210452 106976 210458
rect 106924 210394 106976 210400
rect 106372 129736 106424 129742
rect 106372 129678 106424 129684
rect 106936 85542 106964 210394
rect 108120 209160 108172 209166
rect 108120 209102 108172 209108
rect 108132 208418 108160 209102
rect 107752 208412 107804 208418
rect 107752 208354 107804 208360
rect 108120 208412 108172 208418
rect 108120 208354 108172 208360
rect 107660 180124 107712 180130
rect 107660 180066 107712 180072
rect 107016 158024 107068 158030
rect 107016 157966 107068 157972
rect 107028 90409 107056 157966
rect 107014 90400 107070 90409
rect 107014 90335 107070 90344
rect 107028 88097 107056 90335
rect 107014 88088 107070 88097
rect 107014 88023 107070 88032
rect 106924 85536 106976 85542
rect 106924 85478 106976 85484
rect 106278 71768 106334 71777
rect 106278 71703 106280 71712
rect 106332 71703 106334 71712
rect 106280 71674 106332 71680
rect 106292 71643 106320 71674
rect 107672 60654 107700 180066
rect 107764 98666 107792 208354
rect 107752 98660 107804 98666
rect 107752 98602 107804 98608
rect 107660 60648 107712 60654
rect 107660 60590 107712 60596
rect 107660 49088 107712 49094
rect 107660 49030 107712 49036
rect 106280 28280 106332 28286
rect 106280 28222 106332 28228
rect 106292 16574 106320 28222
rect 107672 16574 107700 49030
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102232 13184 102284 13190
rect 102232 13126 102284 13132
rect 102140 3528 102192 3534
rect 102140 3470 102192 3476
rect 102244 480 102272 13126
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103348 480 103376 3470
rect 104532 3392 104584 3398
rect 104532 3334 104584 3340
rect 104544 480 104572 3334
rect 105740 480 105768 16546
rect 106476 490 106504 16546
rect 106752 598 106964 626
rect 106752 490 106780 598
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 462 106780 490
rect 106936 480 106964 598
rect 108132 480 108160 16546
rect 108316 3466 108344 238031
rect 108408 236065 108436 254351
rect 108394 236056 108450 236065
rect 108394 235991 108450 236000
rect 108394 233200 108450 233209
rect 108394 233135 108450 233144
rect 108408 90545 108436 233135
rect 108500 227050 108528 281522
rect 108960 230450 108988 379471
rect 109052 361593 109080 386990
rect 109144 380186 109172 390102
rect 109512 387054 109540 390374
rect 110708 387122 110736 390374
rect 110800 390374 111136 390402
rect 111996 390374 112608 390402
rect 110800 389298 110828 390374
rect 110788 389292 110840 389298
rect 110788 389234 110840 389240
rect 110696 387116 110748 387122
rect 110696 387058 110748 387064
rect 109500 387048 109552 387054
rect 109500 386990 109552 386996
rect 109132 380180 109184 380186
rect 109132 380122 109184 380128
rect 110800 373994 110828 389234
rect 111064 387048 111116 387054
rect 111064 386990 111116 386996
rect 111076 383654 111104 386990
rect 111064 383648 111116 383654
rect 111064 383590 111116 383596
rect 111996 373994 112024 390374
rect 110616 373966 110828 373994
rect 111812 373966 112024 373994
rect 110512 362228 110564 362234
rect 110512 362170 110564 362176
rect 109038 361584 109094 361593
rect 109038 361519 109094 361528
rect 109052 360233 109080 361519
rect 109038 360224 109094 360233
rect 109038 360159 109094 360168
rect 109682 360224 109738 360233
rect 109682 360159 109738 360168
rect 109040 305652 109092 305658
rect 109040 305594 109092 305600
rect 109052 305046 109080 305594
rect 109040 305040 109092 305046
rect 109040 304982 109092 304988
rect 109052 296714 109080 304982
rect 109052 296686 109172 296714
rect 109038 236056 109094 236065
rect 109038 235991 109094 236000
rect 108948 230444 109000 230450
rect 108948 230386 109000 230392
rect 108488 227044 108540 227050
rect 108488 226986 108540 226992
rect 109052 108322 109080 235991
rect 109144 204950 109172 296686
rect 109696 264994 109724 360159
rect 109684 264988 109736 264994
rect 109684 264930 109736 264936
rect 110524 235958 110552 362170
rect 110616 262002 110644 373966
rect 111064 368484 111116 368490
rect 111064 368426 111116 368432
rect 110604 261996 110656 262002
rect 110604 261938 110656 261944
rect 111076 258058 111104 368426
rect 111812 362914 111840 373966
rect 111800 362908 111852 362914
rect 111800 362850 111852 362856
rect 112536 362908 112588 362914
rect 112536 362850 112588 362856
rect 112548 266422 112576 362850
rect 112626 280800 112682 280809
rect 112626 280735 112682 280744
rect 112536 266416 112588 266422
rect 112442 266384 112498 266393
rect 112536 266358 112588 266364
rect 112442 266319 112498 266328
rect 111800 261520 111852 261526
rect 111800 261462 111852 261468
rect 111064 258052 111116 258058
rect 111064 257994 111116 258000
rect 111064 254040 111116 254046
rect 111064 253982 111116 253988
rect 110604 240780 110656 240786
rect 110604 240722 110656 240728
rect 110616 238377 110644 240722
rect 110602 238368 110658 238377
rect 110602 238303 110658 238312
rect 110512 235952 110564 235958
rect 110512 235894 110564 235900
rect 110418 235240 110474 235249
rect 110418 235175 110474 235184
rect 109224 206372 109276 206378
rect 109224 206314 109276 206320
rect 109236 205766 109264 206314
rect 109224 205760 109276 205766
rect 109224 205702 109276 205708
rect 109132 204944 109184 204950
rect 109132 204886 109184 204892
rect 109132 127628 109184 127634
rect 109132 127570 109184 127576
rect 109144 126274 109172 127570
rect 109132 126268 109184 126274
rect 109132 126210 109184 126216
rect 109040 108316 109092 108322
rect 109040 108258 109092 108264
rect 109236 93838 109264 205702
rect 109684 108316 109736 108322
rect 109684 108258 109736 108264
rect 109224 93832 109276 93838
rect 109224 93774 109276 93780
rect 108394 90536 108450 90545
rect 108394 90471 108450 90480
rect 108408 82822 108436 90471
rect 108396 82816 108448 82822
rect 108396 82758 108448 82764
rect 109696 81394 109724 108258
rect 109684 81388 109736 81394
rect 109684 81330 109736 81336
rect 109040 76560 109092 76566
rect 109040 76502 109092 76508
rect 109052 16574 109080 76502
rect 109052 16546 109356 16574
rect 108304 3460 108356 3466
rect 108304 3402 108356 3408
rect 109328 480 109356 16546
rect 110432 6914 110460 235175
rect 110524 232665 110552 235894
rect 110510 232656 110566 232665
rect 110510 232591 110566 232600
rect 110512 113824 110564 113830
rect 110512 113766 110564 113772
rect 110524 16574 110552 113766
rect 110616 94586 110644 238303
rect 111076 232529 111104 253982
rect 111062 232520 111118 232529
rect 111062 232455 111118 232464
rect 111064 229764 111116 229770
rect 111064 229706 111116 229712
rect 111076 131170 111104 229706
rect 111156 149116 111208 149122
rect 111156 149058 111208 149064
rect 111064 131164 111116 131170
rect 111064 131106 111116 131112
rect 111168 110430 111196 149058
rect 111156 110424 111208 110430
rect 111156 110366 111208 110372
rect 110604 94580 110656 94586
rect 110604 94522 110656 94528
rect 111812 16574 111840 261462
rect 111892 230444 111944 230450
rect 111892 230386 111944 230392
rect 111904 91050 111932 230386
rect 112456 171154 112484 266319
rect 112640 239465 112668 280735
rect 113100 263566 113128 407050
rect 113192 272542 113220 420815
rect 113284 385801 113312 425983
rect 113836 424969 113864 449783
rect 113822 424960 113878 424969
rect 113822 424895 113878 424904
rect 113362 418976 113418 418985
rect 113362 418911 113418 418920
rect 113270 385792 113326 385801
rect 113270 385727 113326 385736
rect 113376 381614 113404 418911
rect 114480 406473 114508 467842
rect 114650 420064 114706 420073
rect 114650 419999 114706 420008
rect 114558 417888 114614 417897
rect 114558 417823 114614 417832
rect 114466 406464 114522 406473
rect 114466 406399 114522 406408
rect 113454 402384 113510 402393
rect 113454 402319 113510 402328
rect 113468 383722 113496 402319
rect 113456 383716 113508 383722
rect 113456 383658 113508 383664
rect 113364 381608 113416 381614
rect 113364 381550 113416 381556
rect 113468 373994 113496 383658
rect 113284 373966 113496 373994
rect 113284 368490 113312 373966
rect 113272 368484 113324 368490
rect 113272 368426 113324 368432
rect 114468 280220 114520 280226
rect 114468 280162 114520 280168
rect 113180 272536 113232 272542
rect 113180 272478 113232 272484
rect 114480 271153 114508 280162
rect 114572 271250 114600 417823
rect 114664 280226 114692 419999
rect 114756 413953 114784 551278
rect 115202 516760 115258 516769
rect 115202 516695 115258 516704
rect 115216 463593 115244 516695
rect 115202 463584 115258 463593
rect 115202 463519 115258 463528
rect 114834 430128 114890 430137
rect 114834 430063 114890 430072
rect 114742 413944 114798 413953
rect 114742 413879 114798 413888
rect 114756 413642 114784 413879
rect 114744 413636 114796 413642
rect 114744 413578 114796 413584
rect 114848 382945 114876 430063
rect 115216 421977 115244 463519
rect 115756 434716 115808 434722
rect 115756 434658 115808 434664
rect 115768 433401 115796 434658
rect 115754 433392 115810 433401
rect 115754 433327 115810 433336
rect 115848 433288 115900 433294
rect 115848 433230 115900 433236
rect 115860 432313 115888 433230
rect 115846 432304 115902 432313
rect 115846 432239 115902 432248
rect 115572 431928 115624 431934
rect 115572 431870 115624 431876
rect 115584 431225 115612 431870
rect 115570 431216 115626 431225
rect 115570 431151 115626 431160
rect 115756 430568 115808 430574
rect 115756 430510 115808 430516
rect 115768 429321 115796 430510
rect 115754 429312 115810 429321
rect 115754 429247 115810 429256
rect 115848 429140 115900 429146
rect 115848 429082 115900 429088
rect 115860 428233 115888 429082
rect 115846 428224 115902 428233
rect 115846 428159 115902 428168
rect 115848 426420 115900 426426
rect 115848 426362 115900 426368
rect 115860 426057 115888 426362
rect 115846 426048 115902 426057
rect 115846 425983 115902 425992
rect 115848 425060 115900 425066
rect 115848 425002 115900 425008
rect 115860 424153 115888 425002
rect 115846 424144 115902 424153
rect 115846 424079 115902 424088
rect 115848 423632 115900 423638
rect 115848 423574 115900 423580
rect 115860 423065 115888 423574
rect 115846 423056 115902 423065
rect 115846 422991 115902 423000
rect 115202 421968 115258 421977
rect 115202 421903 115258 421912
rect 115848 419416 115900 419422
rect 115848 419358 115900 419364
rect 115860 418985 115888 419358
rect 115846 418976 115902 418985
rect 115846 418911 115902 418920
rect 115848 416832 115900 416838
rect 115846 416800 115848 416809
rect 115900 416800 115902 416809
rect 115846 416735 115902 416744
rect 115846 415712 115902 415721
rect 115846 415647 115902 415656
rect 115860 415478 115888 415647
rect 115848 415472 115900 415478
rect 115848 415414 115900 415420
rect 115846 414896 115902 414905
rect 115846 414831 115902 414840
rect 115860 414730 115888 414831
rect 115848 414724 115900 414730
rect 115848 414666 115900 414672
rect 115756 413976 115808 413982
rect 115756 413918 115808 413924
rect 115768 412729 115796 413918
rect 115754 412720 115810 412729
rect 115754 412655 115810 412664
rect 115020 411936 115072 411942
rect 115020 411878 115072 411884
rect 115032 411641 115060 411878
rect 115018 411632 115074 411641
rect 115018 411567 115074 411576
rect 115572 411256 115624 411262
rect 115572 411198 115624 411204
rect 115584 410553 115612 411198
rect 115570 410544 115626 410553
rect 115570 410479 115626 410488
rect 115848 409828 115900 409834
rect 115848 409770 115900 409776
rect 115860 409737 115888 409770
rect 115846 409728 115902 409737
rect 115846 409663 115902 409672
rect 115846 408640 115902 408649
rect 115846 408575 115902 408584
rect 115860 408542 115888 408575
rect 115848 408536 115900 408542
rect 115848 408478 115900 408484
rect 115202 406464 115258 406473
rect 115202 406399 115258 406408
rect 115112 396568 115164 396574
rect 115112 396510 115164 396516
rect 115124 396409 115152 396510
rect 115110 396400 115166 396409
rect 115110 396335 115166 396344
rect 114834 382936 114890 382945
rect 114834 382871 114890 382880
rect 115216 321706 115244 406399
rect 115848 405680 115900 405686
rect 115846 405648 115848 405657
rect 115900 405648 115902 405657
rect 115846 405583 115902 405592
rect 115846 404560 115902 404569
rect 115846 404495 115902 404504
rect 115860 404394 115888 404495
rect 115848 404388 115900 404394
rect 115848 404330 115900 404336
rect 115846 403472 115902 403481
rect 115846 403407 115902 403416
rect 115860 403034 115888 403407
rect 115848 403028 115900 403034
rect 115848 402970 115900 402976
rect 115754 401296 115810 401305
rect 115754 401231 115810 401240
rect 115572 400716 115624 400722
rect 115572 400658 115624 400664
rect 115584 400489 115612 400658
rect 115768 400586 115796 401231
rect 115756 400580 115808 400586
rect 115756 400522 115808 400528
rect 115570 400480 115626 400489
rect 115570 400415 115626 400424
rect 115846 399392 115902 399401
rect 115846 399327 115902 399336
rect 115860 398954 115888 399327
rect 115848 398948 115900 398954
rect 115848 398890 115900 398896
rect 115848 398336 115900 398342
rect 115846 398304 115848 398313
rect 116032 398336 116084 398342
rect 115900 398304 115902 398313
rect 116032 398278 116084 398284
rect 115846 398239 115902 398248
rect 115570 397216 115626 397225
rect 115570 397151 115626 397160
rect 115584 396098 115612 397151
rect 115572 396092 115624 396098
rect 115572 396034 115624 396040
rect 115846 395312 115902 395321
rect 115846 395247 115902 395256
rect 115860 394806 115888 395247
rect 115848 394800 115900 394806
rect 115848 394742 115900 394748
rect 115848 394664 115900 394670
rect 115848 394606 115900 394612
rect 115860 394233 115888 394606
rect 115846 394224 115902 394233
rect 115846 394159 115902 394168
rect 115846 393136 115902 393145
rect 115902 393094 115980 393122
rect 115846 393071 115902 393080
rect 115952 392358 115980 393094
rect 115940 392352 115992 392358
rect 115940 392294 115992 392300
rect 115846 392048 115902 392057
rect 115846 391983 115848 391992
rect 115900 391983 115902 391992
rect 115848 391954 115900 391960
rect 115952 373386 115980 392294
rect 116044 376038 116072 398278
rect 116136 385665 116164 553959
rect 116596 538218 116624 575486
rect 119356 538898 119384 582655
rect 122116 551342 122144 583714
rect 122208 563718 122236 585142
rect 123484 582480 123536 582486
rect 123484 582422 123536 582428
rect 122196 563712 122248 563718
rect 122196 563654 122248 563660
rect 122748 563712 122800 563718
rect 122748 563654 122800 563660
rect 122104 551336 122156 551342
rect 122104 551278 122156 551284
rect 119344 538892 119396 538898
rect 119344 538834 119396 538840
rect 116584 538212 116636 538218
rect 116584 538154 116636 538160
rect 118700 523728 118752 523734
rect 118700 523670 118752 523676
rect 116584 469872 116636 469878
rect 116584 469814 116636 469820
rect 116596 449857 116624 469814
rect 118606 456920 118662 456929
rect 118606 456855 118662 456864
rect 116582 449848 116638 449857
rect 116582 449783 116638 449792
rect 118620 436801 118648 456855
rect 118606 436792 118662 436801
rect 118606 436727 118662 436736
rect 118712 423638 118740 523670
rect 119342 452840 119398 452849
rect 119342 452775 119398 452784
rect 119356 438161 119384 452775
rect 119342 438152 119398 438161
rect 119342 438087 119398 438096
rect 118790 436792 118846 436801
rect 118790 436727 118846 436736
rect 118700 423632 118752 423638
rect 118700 423574 118752 423580
rect 118700 417240 118752 417246
rect 118700 417182 118752 417188
rect 118712 416838 118740 417182
rect 118700 416832 118752 416838
rect 118700 416774 118752 416780
rect 117320 413636 117372 413642
rect 117320 413578 117372 413584
rect 116584 401668 116636 401674
rect 116584 401610 116636 401616
rect 116596 391338 116624 401610
rect 117228 393984 117280 393990
rect 117228 393926 117280 393932
rect 117240 392358 117268 393926
rect 117228 392352 117280 392358
rect 117228 392294 117280 392300
rect 116584 391332 116636 391338
rect 116584 391274 116636 391280
rect 116122 385656 116178 385665
rect 116122 385591 116178 385600
rect 116584 384328 116636 384334
rect 116584 384270 116636 384276
rect 116032 376032 116084 376038
rect 116032 375974 116084 375980
rect 115940 373380 115992 373386
rect 115940 373322 115992 373328
rect 115204 321700 115256 321706
rect 115204 321642 115256 321648
rect 115216 312662 115244 321642
rect 115204 312656 115256 312662
rect 115204 312598 115256 312604
rect 115938 301472 115994 301481
rect 115938 301407 115994 301416
rect 115388 296744 115440 296750
rect 115388 296686 115440 296692
rect 114652 280220 114704 280226
rect 114652 280162 114704 280168
rect 114560 271244 114612 271250
rect 114560 271186 114612 271192
rect 114466 271144 114522 271153
rect 114466 271079 114522 271088
rect 115296 268388 115348 268394
rect 115296 268330 115348 268336
rect 113824 263628 113876 263634
rect 113824 263570 113876 263576
rect 113088 263560 113140 263566
rect 113088 263502 113140 263508
rect 113836 244905 113864 263570
rect 113914 247616 113970 247625
rect 113914 247551 113970 247560
rect 113822 244896 113878 244905
rect 113822 244831 113878 244840
rect 112626 239456 112682 239465
rect 112626 239391 112682 239400
rect 113180 238060 113232 238066
rect 113180 238002 113232 238008
rect 112444 171148 112496 171154
rect 112444 171090 112496 171096
rect 112456 120086 112484 171090
rect 112444 120080 112496 120086
rect 112444 120022 112496 120028
rect 112444 108316 112496 108322
rect 112444 108258 112496 108264
rect 111892 91044 111944 91050
rect 111892 90986 111944 90992
rect 111904 88262 111932 90986
rect 111892 88256 111944 88262
rect 111892 88198 111944 88204
rect 112456 79966 112484 108258
rect 113192 92313 113220 238002
rect 113928 237289 113956 247551
rect 113914 237280 113970 237289
rect 113914 237215 113970 237224
rect 115202 235376 115258 235385
rect 115202 235311 115258 235320
rect 114652 231124 114704 231130
rect 114652 231066 114704 231072
rect 113272 206304 113324 206310
rect 113272 206246 113324 206252
rect 113916 206304 113968 206310
rect 113916 206246 113968 206252
rect 113284 108390 113312 206246
rect 113928 205698 113956 206246
rect 113916 205692 113968 205698
rect 113916 205634 113968 205640
rect 114560 129124 114612 129130
rect 114560 129066 114612 129072
rect 113272 108384 113324 108390
rect 113272 108326 113324 108332
rect 113178 92304 113234 92313
rect 113178 92239 113234 92248
rect 112444 79960 112496 79966
rect 112444 79902 112496 79908
rect 113180 37936 113232 37942
rect 113180 37878 113232 37884
rect 113192 16574 113220 37878
rect 114572 16574 114600 129066
rect 114664 96694 114692 231066
rect 114652 96688 114704 96694
rect 114652 96630 114704 96636
rect 115216 88233 115244 235311
rect 115308 169794 115336 268330
rect 115400 231169 115428 296686
rect 115480 269136 115532 269142
rect 115480 269078 115532 269084
rect 115492 235958 115520 269078
rect 115480 235952 115532 235958
rect 115480 235894 115532 235900
rect 115386 231160 115442 231169
rect 115386 231095 115442 231104
rect 115296 169788 115348 169794
rect 115296 169730 115348 169736
rect 115308 138689 115336 169730
rect 115294 138680 115350 138689
rect 115294 138615 115350 138624
rect 115848 96688 115900 96694
rect 115848 96630 115900 96636
rect 115860 95946 115888 96630
rect 115848 95940 115900 95946
rect 115848 95882 115900 95888
rect 115202 88224 115258 88233
rect 115202 88159 115258 88168
rect 115952 16574 115980 301407
rect 116596 233170 116624 384270
rect 117332 378729 117360 413578
rect 118712 389881 118740 416774
rect 118698 389872 118754 389881
rect 118698 389807 118754 389816
rect 117962 387152 118018 387161
rect 117962 387087 118018 387096
rect 117318 378720 117374 378729
rect 117318 378655 117374 378664
rect 117976 372638 118004 387087
rect 118700 382968 118752 382974
rect 118700 382910 118752 382916
rect 117964 372632 118016 372638
rect 117964 372574 118016 372580
rect 116768 339584 116820 339590
rect 116768 339526 116820 339532
rect 116676 236700 116728 236706
rect 116676 236642 116728 236648
rect 116584 233164 116636 233170
rect 116584 233106 116636 233112
rect 116030 232656 116086 232665
rect 116030 232591 116086 232600
rect 116044 62014 116072 232591
rect 116688 86970 116716 236642
rect 116780 234569 116808 339526
rect 117976 235385 118004 372574
rect 118056 285728 118108 285734
rect 118056 285670 118108 285676
rect 118068 267034 118096 285670
rect 118056 267028 118108 267034
rect 118056 266970 118108 266976
rect 118712 236706 118740 382910
rect 118804 305658 118832 436727
rect 119344 427100 119396 427106
rect 119344 427042 119396 427048
rect 119356 417246 119384 427042
rect 119344 417240 119396 417246
rect 119344 417182 119396 417188
rect 120080 416084 120132 416090
rect 120080 416026 120132 416032
rect 120092 415478 120120 416026
rect 120080 415472 120132 415478
rect 120080 415414 120132 415420
rect 122196 415472 122248 415478
rect 122196 415414 122248 415420
rect 119988 403640 120040 403646
rect 119988 403582 120040 403588
rect 118884 400920 118936 400926
rect 118884 400862 118936 400868
rect 118896 398342 118924 400862
rect 120000 400722 120028 403582
rect 119988 400716 120040 400722
rect 119988 400658 120040 400664
rect 118884 398336 118936 398342
rect 118884 398278 118936 398284
rect 118884 398200 118936 398206
rect 118884 398142 118936 398148
rect 118896 396574 118924 398142
rect 118884 396568 118936 396574
rect 118884 396510 118936 396516
rect 120092 380905 120120 415414
rect 122208 411262 122236 415414
rect 122760 414730 122788 563654
rect 123496 541754 123524 582422
rect 123484 541748 123536 541754
rect 123484 541690 123536 541696
rect 122840 525088 122892 525094
rect 122840 525030 122892 525036
rect 122748 414724 122800 414730
rect 122748 414666 122800 414672
rect 122852 411942 122880 525030
rect 124232 426426 124260 589290
rect 125600 588668 125652 588674
rect 125600 588610 125652 588616
rect 124864 431248 124916 431254
rect 124864 431190 124916 431196
rect 124220 426420 124272 426426
rect 124220 426362 124272 426368
rect 122840 411936 122892 411942
rect 122840 411878 122892 411884
rect 123484 411936 123536 411942
rect 123484 411878 123536 411884
rect 122196 411256 122248 411262
rect 122196 411198 122248 411204
rect 121460 409896 121512 409902
rect 121460 409838 121512 409844
rect 121472 405686 121500 409838
rect 121460 405680 121512 405686
rect 121460 405622 121512 405628
rect 122196 400580 122248 400586
rect 122196 400522 122248 400528
rect 122104 396092 122156 396098
rect 122104 396034 122156 396040
rect 120078 380896 120134 380905
rect 120078 380831 120134 380840
rect 120724 377460 120776 377466
rect 120724 377402 120776 377408
rect 118792 305652 118844 305658
rect 118792 305594 118844 305600
rect 119344 305652 119396 305658
rect 119344 305594 119396 305600
rect 118884 278044 118936 278050
rect 118884 277986 118936 277992
rect 118700 236700 118752 236706
rect 118700 236642 118752 236648
rect 117962 235376 118018 235385
rect 117962 235311 118018 235320
rect 116766 234560 116822 234569
rect 116766 234495 116822 234504
rect 117412 213240 117464 213246
rect 117412 213182 117464 213188
rect 117424 212566 117452 213182
rect 117412 212560 117464 212566
rect 117412 212502 117464 212508
rect 117318 206272 117374 206281
rect 117318 206207 117374 206216
rect 116676 86964 116728 86970
rect 116676 86906 116728 86912
rect 116032 62008 116084 62014
rect 116032 61950 116084 61956
rect 117332 16574 117360 206207
rect 117424 101454 117452 212502
rect 118792 185632 118844 185638
rect 118792 185574 118844 185580
rect 117412 101448 117464 101454
rect 117412 101390 117464 101396
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 117332 16546 117636 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 112364 490 112392 16546
rect 112640 598 112852 626
rect 112640 490 112668 598
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 462 112668 490
rect 112824 480 112852 598
rect 114020 480 114048 16546
rect 114756 490 114784 16546
rect 115032 598 115244 626
rect 115032 490 115060 598
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 462 115060 490
rect 115216 480 115244 598
rect 116412 480 116440 16546
rect 117608 480 117636 16546
rect 118804 480 118832 185574
rect 118896 140078 118924 277986
rect 118976 236292 119028 236298
rect 118976 236234 119028 236240
rect 118884 140072 118936 140078
rect 118884 140014 118936 140020
rect 118896 139466 118924 140014
rect 118884 139460 118936 139466
rect 118884 139402 118936 139408
rect 118988 16574 119016 236234
rect 119356 229770 119384 305594
rect 120736 234598 120764 377402
rect 122116 376689 122144 396034
rect 122102 376680 122158 376689
rect 122102 376615 122158 376624
rect 122104 345160 122156 345166
rect 122104 345102 122156 345108
rect 121460 302932 121512 302938
rect 121460 302874 121512 302880
rect 120816 268388 120868 268394
rect 120816 268330 120868 268336
rect 120724 234592 120776 234598
rect 120724 234534 120776 234540
rect 119344 229764 119396 229770
rect 119344 229706 119396 229712
rect 119342 228304 119398 228313
rect 119342 228239 119398 228248
rect 119356 215966 119384 228239
rect 120172 217320 120224 217326
rect 120172 217262 120224 217268
rect 119344 215960 119396 215966
rect 119344 215902 119396 215908
rect 120078 185600 120134 185609
rect 120078 185535 120134 185544
rect 120092 74526 120120 185535
rect 120184 105602 120212 217262
rect 120828 186998 120856 268330
rect 120816 186992 120868 186998
rect 120816 186934 120868 186940
rect 120724 142860 120776 142866
rect 120724 142802 120776 142808
rect 120736 140146 120764 142802
rect 120724 140140 120776 140146
rect 120724 140082 120776 140088
rect 120172 105596 120224 105602
rect 120172 105538 120224 105544
rect 120724 100768 120776 100774
rect 120724 100710 120776 100716
rect 120736 84017 120764 100710
rect 120722 84008 120778 84017
rect 120722 83943 120778 83952
rect 120080 74520 120132 74526
rect 120080 74462 120132 74468
rect 120080 29708 120132 29714
rect 120080 29650 120132 29656
rect 120092 16574 120120 29650
rect 121472 16574 121500 302874
rect 121552 291236 121604 291242
rect 121552 291178 121604 291184
rect 121564 175982 121592 291178
rect 122116 251161 122144 345102
rect 122208 307154 122236 400522
rect 123496 378729 123524 411878
rect 123574 409184 123630 409193
rect 123574 409119 123630 409128
rect 123588 389201 123616 409119
rect 123668 400240 123720 400246
rect 123668 400182 123720 400188
rect 123574 389192 123630 389201
rect 123574 389127 123630 389136
rect 123576 387864 123628 387870
rect 123576 387806 123628 387812
rect 123482 378720 123538 378729
rect 123482 378655 123538 378664
rect 123588 364274 123616 387806
rect 123680 379409 123708 400182
rect 123666 379400 123722 379409
rect 123666 379335 123722 379344
rect 123576 364268 123628 364274
rect 123576 364210 123628 364216
rect 122840 358080 122892 358086
rect 122840 358022 122892 358028
rect 123760 358080 123812 358086
rect 123760 358022 123812 358028
rect 122196 307148 122248 307154
rect 122196 307090 122248 307096
rect 122102 251152 122158 251161
rect 122102 251087 122158 251096
rect 122196 250504 122248 250510
rect 122196 250446 122248 250452
rect 122208 235929 122236 250446
rect 122852 238066 122880 358022
rect 123772 357474 123800 358022
rect 123760 357468 123812 357474
rect 123760 357410 123812 357416
rect 124876 342582 124904 431190
rect 125612 387870 125640 588610
rect 130476 582412 130528 582418
rect 130476 582354 130528 582360
rect 130384 567860 130436 567866
rect 130384 567802 130436 567808
rect 130396 567254 130424 567802
rect 130384 567248 130436 567254
rect 130384 567190 130436 567196
rect 129004 532024 129056 532030
rect 129004 531966 129056 531972
rect 127624 494760 127676 494766
rect 127624 494702 127676 494708
rect 126244 478168 126296 478174
rect 126244 478110 126296 478116
rect 126256 431934 126284 478110
rect 126244 431928 126296 431934
rect 126244 431870 126296 431876
rect 126244 416832 126296 416838
rect 126244 416774 126296 416780
rect 125692 414724 125744 414730
rect 125692 414666 125744 414672
rect 125600 387864 125652 387870
rect 125600 387806 125652 387812
rect 124864 342576 124916 342582
rect 124864 342518 124916 342524
rect 125508 342576 125560 342582
rect 125508 342518 125560 342524
rect 125520 342310 125548 342518
rect 125508 342304 125560 342310
rect 125508 342246 125560 342252
rect 124864 313336 124916 313342
rect 124864 313278 124916 313284
rect 123576 304360 123628 304366
rect 123576 304302 123628 304308
rect 122932 297424 122984 297430
rect 122932 297366 122984 297372
rect 122944 293962 122972 297366
rect 122932 293956 122984 293962
rect 122932 293898 122984 293904
rect 123484 279472 123536 279478
rect 123484 279414 123536 279420
rect 122840 238060 122892 238066
rect 122840 238002 122892 238008
rect 122194 235920 122250 235929
rect 122194 235855 122250 235864
rect 122932 234592 122984 234598
rect 122932 234534 122984 234540
rect 122196 233164 122248 233170
rect 122196 233106 122248 233112
rect 122104 182912 122156 182918
rect 122104 182854 122156 182860
rect 121552 175976 121604 175982
rect 121552 175918 121604 175924
rect 122116 38010 122144 182854
rect 122208 89690 122236 233106
rect 122840 180124 122892 180130
rect 122840 180066 122892 180072
rect 122196 89684 122248 89690
rect 122196 89626 122248 89632
rect 122208 84182 122236 89626
rect 122196 84176 122248 84182
rect 122196 84118 122248 84124
rect 122104 38004 122156 38010
rect 122104 37946 122156 37952
rect 122852 16574 122880 180066
rect 122944 89593 122972 234534
rect 123496 231130 123524 279414
rect 123484 231124 123536 231130
rect 123484 231066 123536 231072
rect 123484 193860 123536 193866
rect 123484 193802 123536 193808
rect 122930 89584 122986 89593
rect 122930 89519 122986 89528
rect 123496 66910 123524 193802
rect 123588 192545 123616 304302
rect 124218 237960 124274 237969
rect 124218 237895 124274 237904
rect 123574 192536 123630 192545
rect 123574 192471 123630 192480
rect 123484 66904 123536 66910
rect 123484 66846 123536 66852
rect 124232 16574 124260 237895
rect 124312 182844 124364 182850
rect 124312 182786 124364 182792
rect 124324 94518 124352 182786
rect 124876 149734 124904 313278
rect 124954 309768 125010 309777
rect 124954 309703 125010 309712
rect 124968 236298 124996 309703
rect 125520 308446 125548 342246
rect 125704 320890 125732 414666
rect 126256 409834 126284 416774
rect 127636 413982 127664 494702
rect 127624 413976 127676 413982
rect 127624 413918 127676 413924
rect 126244 409828 126296 409834
rect 126244 409770 126296 409776
rect 129016 398886 129044 531966
rect 129096 451308 129148 451314
rect 129096 451250 129148 451256
rect 129004 398880 129056 398886
rect 129004 398822 129056 398828
rect 129016 383625 129044 398822
rect 129002 383616 129058 383625
rect 129002 383551 129058 383560
rect 129004 380180 129056 380186
rect 129004 380122 129056 380128
rect 129016 356726 129044 380122
rect 129004 356720 129056 356726
rect 129004 356662 129056 356668
rect 129002 337376 129058 337385
rect 129002 337311 129058 337320
rect 126242 336016 126298 336025
rect 126242 335951 126298 335960
rect 125692 320884 125744 320890
rect 125692 320826 125744 320832
rect 125508 308440 125560 308446
rect 125508 308382 125560 308388
rect 125046 291816 125102 291825
rect 125046 291751 125102 291760
rect 125060 243574 125088 291751
rect 125600 253972 125652 253978
rect 125600 253914 125652 253920
rect 125048 243568 125100 243574
rect 125048 243510 125100 243516
rect 124956 236292 125008 236298
rect 124956 236234 125008 236240
rect 124954 153232 125010 153241
rect 124954 153167 125010 153176
rect 124864 149728 124916 149734
rect 124864 149670 124916 149676
rect 124968 124137 124996 153167
rect 124954 124128 125010 124137
rect 124954 124063 125010 124072
rect 124312 94512 124364 94518
rect 124312 94454 124364 94460
rect 125612 89842 125640 253914
rect 125520 89814 125640 89842
rect 125520 86902 125548 89814
rect 124864 86896 124916 86902
rect 124864 86838 124916 86844
rect 125508 86896 125560 86902
rect 125508 86838 125560 86844
rect 124876 69018 124904 86838
rect 124864 69012 124916 69018
rect 124864 68954 124916 68960
rect 126256 49094 126284 335951
rect 127624 330540 127676 330546
rect 127624 330482 127676 330488
rect 126888 321564 126940 321570
rect 126888 321506 126940 321512
rect 126900 320890 126928 321506
rect 126888 320884 126940 320890
rect 126888 320826 126940 320832
rect 126336 311228 126388 311234
rect 126336 311170 126388 311176
rect 126348 79393 126376 311170
rect 126426 296168 126482 296177
rect 126426 296103 126482 296112
rect 126440 257378 126468 296103
rect 126428 257372 126480 257378
rect 126428 257314 126480 257320
rect 126888 254584 126940 254590
rect 126888 254526 126940 254532
rect 126900 253978 126928 254526
rect 126888 253972 126940 253978
rect 126888 253914 126940 253920
rect 126980 240848 127032 240854
rect 126980 240790 127032 240796
rect 126992 240174 127020 240790
rect 126980 240168 127032 240174
rect 126980 240110 127032 240116
rect 126992 95849 127020 240110
rect 127636 119377 127664 330482
rect 128268 284368 128320 284374
rect 128268 284310 128320 284316
rect 128280 252550 128308 284310
rect 128268 252544 128320 252550
rect 128268 252486 128320 252492
rect 129016 129033 129044 337311
rect 129108 313954 129136 451250
rect 129740 385008 129792 385014
rect 129740 384950 129792 384956
rect 129752 384334 129780 384950
rect 129740 384328 129792 384334
rect 129740 384270 129792 384276
rect 129740 369844 129792 369850
rect 129740 369786 129792 369792
rect 129752 369238 129780 369786
rect 130396 369238 130424 567190
rect 130488 534070 130516 582354
rect 130476 534064 130528 534070
rect 130476 534006 130528 534012
rect 130936 534064 130988 534070
rect 130936 534006 130988 534012
rect 130948 385014 130976 534006
rect 131028 525156 131080 525162
rect 131028 525098 131080 525104
rect 130936 385008 130988 385014
rect 130936 384950 130988 384956
rect 129740 369232 129792 369238
rect 129740 369174 129792 369180
rect 130384 369232 130436 369238
rect 130384 369174 130436 369180
rect 130382 325000 130438 325009
rect 130382 324935 130438 324944
rect 129186 317520 129242 317529
rect 129186 317455 129242 317464
rect 129096 313948 129148 313954
rect 129096 313890 129148 313896
rect 129108 313342 129136 313890
rect 129096 313336 129148 313342
rect 129096 313278 129148 313284
rect 129200 301578 129228 317455
rect 129188 301572 129240 301578
rect 129188 301514 129240 301520
rect 129188 300212 129240 300218
rect 129188 300154 129240 300160
rect 129096 276072 129148 276078
rect 129096 276014 129148 276020
rect 129108 198694 129136 276014
rect 129200 261526 129228 300154
rect 129188 261520 129240 261526
rect 129188 261462 129240 261468
rect 129740 252544 129792 252550
rect 129740 252486 129792 252492
rect 129188 249076 129240 249082
rect 129188 249018 129240 249024
rect 129096 198688 129148 198694
rect 129096 198630 129148 198636
rect 129096 195288 129148 195294
rect 129096 195230 129148 195236
rect 129002 129024 129058 129033
rect 129002 128959 129058 128968
rect 127622 119368 127678 119377
rect 127622 119303 127678 119312
rect 127622 118008 127678 118017
rect 127622 117943 127678 117952
rect 126978 95840 127034 95849
rect 126978 95775 127034 95784
rect 126334 79384 126390 79393
rect 126334 79319 126390 79328
rect 127636 68241 127664 117943
rect 127622 68232 127678 68241
rect 127622 68167 127678 68176
rect 126244 49088 126296 49094
rect 126244 49030 126296 49036
rect 125600 32428 125652 32434
rect 125600 32370 125652 32376
rect 125612 16574 125640 32370
rect 129108 16574 129136 195230
rect 129200 102134 129228 249018
rect 129188 102128 129240 102134
rect 129188 102070 129240 102076
rect 129200 101454 129228 102070
rect 129188 101448 129240 101454
rect 129188 101390 129240 101396
rect 129752 99498 129780 252486
rect 129660 99470 129780 99498
rect 129660 99414 129688 99470
rect 129648 99408 129700 99414
rect 129648 99350 129700 99356
rect 129660 73098 129688 99350
rect 129648 73092 129700 73098
rect 129648 73034 129700 73040
rect 118988 16546 119936 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 125612 16546 125916 16574
rect 129108 16546 129412 16574
rect 119908 480 119936 16546
rect 120644 490 120672 16546
rect 120920 598 121132 626
rect 120920 490 120948 598
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 462 120948 490
rect 121104 480 121132 598
rect 122300 480 122328 16546
rect 123036 490 123064 16546
rect 123312 598 123524 626
rect 123312 490 123340 598
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 462 123340 490
rect 123496 480 123524 598
rect 124692 480 124720 16546
rect 125888 480 125916 16546
rect 129384 480 129412 16546
rect 130396 2106 130424 324935
rect 130474 322960 130530 322969
rect 130474 322895 130530 322904
rect 130488 280158 130516 322895
rect 130476 280152 130528 280158
rect 130476 280094 130528 280100
rect 130474 276720 130530 276729
rect 130474 276655 130530 276664
rect 130488 29646 130516 276655
rect 131040 253910 131068 525098
rect 132408 492720 132460 492726
rect 132408 492662 132460 492668
rect 131764 447840 131816 447846
rect 131764 447782 131816 447788
rect 131776 407114 131804 447782
rect 131764 407108 131816 407114
rect 131764 407050 131816 407056
rect 131120 308440 131172 308446
rect 131120 308382 131172 308388
rect 131028 253904 131080 253910
rect 131028 253846 131080 253852
rect 131132 153950 131160 308382
rect 132420 297430 132448 492662
rect 133708 475250 133736 597518
rect 134524 578264 134576 578270
rect 134524 578206 134576 578212
rect 133786 530632 133842 530641
rect 133786 530567 133842 530576
rect 133144 475244 133196 475250
rect 133144 475186 133196 475192
rect 133696 475244 133748 475250
rect 133696 475186 133748 475192
rect 132500 434036 132552 434042
rect 132500 433978 132552 433984
rect 132408 297424 132460 297430
rect 132408 297366 132460 297372
rect 131764 193928 131816 193934
rect 131764 193870 131816 193876
rect 131120 153944 131172 153950
rect 131120 153886 131172 153892
rect 131776 51746 131804 193870
rect 131856 151904 131908 151910
rect 131856 151846 131908 151852
rect 131868 121446 131896 151846
rect 131856 121440 131908 121446
rect 131856 121382 131908 121388
rect 131764 51740 131816 51746
rect 131764 51682 131816 51688
rect 130476 29640 130528 29646
rect 130476 29582 130528 29588
rect 132512 16574 132540 433978
rect 133156 427106 133184 475186
rect 133708 474774 133736 475186
rect 133696 474768 133748 474774
rect 133696 474710 133748 474716
rect 133236 473408 133288 473414
rect 133236 473350 133288 473356
rect 133248 430574 133276 473350
rect 133236 430568 133288 430574
rect 133236 430510 133288 430516
rect 133144 427100 133196 427106
rect 133144 427042 133196 427048
rect 133142 327856 133198 327865
rect 133142 327791 133198 327800
rect 133156 268394 133184 327791
rect 133696 271176 133748 271182
rect 133696 271118 133748 271124
rect 133708 270502 133736 271118
rect 133696 270496 133748 270502
rect 133696 270438 133748 270444
rect 133144 268388 133196 268394
rect 133144 268330 133196 268336
rect 133142 265024 133198 265033
rect 133142 264959 133198 264968
rect 133156 236609 133184 264959
rect 133142 236600 133198 236609
rect 133142 236535 133198 236544
rect 133144 185700 133196 185706
rect 133144 185642 133196 185648
rect 133156 49026 133184 185642
rect 133708 162042 133736 270438
rect 133800 262138 133828 530567
rect 133788 262132 133840 262138
rect 133788 262074 133840 262080
rect 133236 162036 133288 162042
rect 133236 161978 133288 161984
rect 133696 162036 133748 162042
rect 133696 161978 133748 161984
rect 133248 161566 133276 161978
rect 133236 161560 133288 161566
rect 133236 161502 133288 161508
rect 133248 127634 133276 161502
rect 133236 127628 133288 127634
rect 133236 127570 133288 127576
rect 133144 49020 133196 49026
rect 133144 48962 133196 48968
rect 132512 16546 133000 16574
rect 130384 2100 130436 2106
rect 130384 2042 130436 2048
rect 132972 480 133000 16546
rect 134536 4214 134564 578206
rect 137100 573368 137152 573374
rect 137100 573310 137152 573316
rect 137112 572762 137140 573310
rect 136640 572756 136692 572762
rect 136640 572698 136692 572704
rect 137100 572756 137152 572762
rect 137100 572698 137152 572704
rect 134616 539640 134668 539646
rect 134616 539582 134668 539588
rect 134628 386306 134656 539582
rect 135902 538248 135958 538257
rect 135902 538183 135958 538192
rect 134616 386300 134668 386306
rect 134616 386242 134668 386248
rect 135168 386300 135220 386306
rect 135168 386242 135220 386248
rect 135180 385762 135208 386242
rect 135168 385756 135220 385762
rect 135168 385698 135220 385704
rect 135916 383654 135944 538183
rect 136548 505776 136600 505782
rect 136548 505718 136600 505724
rect 135904 383648 135956 383654
rect 135904 383590 135956 383596
rect 135916 383042 135944 383590
rect 135904 383036 135956 383042
rect 135904 382978 135956 382984
rect 134616 346520 134668 346526
rect 134616 346462 134668 346468
rect 134628 113830 134656 346462
rect 134706 334656 134762 334665
rect 134706 334591 134762 334600
rect 134720 182918 134748 334591
rect 135902 331936 135958 331945
rect 135902 331871 135958 331880
rect 134708 182912 134760 182918
rect 134708 182854 134760 182860
rect 134706 153232 134762 153241
rect 134706 153167 134762 153176
rect 134720 118658 134748 153167
rect 134708 118652 134760 118658
rect 134708 118594 134760 118600
rect 134616 113824 134668 113830
rect 134616 113766 134668 113772
rect 135916 11762 135944 331871
rect 136088 274712 136140 274718
rect 136088 274654 136140 274660
rect 135996 272604 136048 272610
rect 135996 272546 136048 272552
rect 136008 76566 136036 272546
rect 136100 257378 136128 274654
rect 136560 271862 136588 505718
rect 136652 393990 136680 572698
rect 137744 461644 137796 461650
rect 137744 461586 137796 461592
rect 137284 398948 137336 398954
rect 137284 398890 137336 398896
rect 136640 393984 136692 393990
rect 136640 393926 136692 393932
rect 137296 365673 137324 398890
rect 137756 367033 137784 461586
rect 137836 459672 137888 459678
rect 137836 459614 137888 459620
rect 137848 445738 137876 459614
rect 137836 445732 137888 445738
rect 137836 445674 137888 445680
rect 137834 392592 137890 392601
rect 137834 392527 137890 392536
rect 137466 367024 137522 367033
rect 137466 366959 137468 366968
rect 137520 366959 137522 366968
rect 137742 367024 137798 367033
rect 137742 366959 137798 366968
rect 137468 366930 137520 366936
rect 137282 365664 137338 365673
rect 137282 365599 137338 365608
rect 137376 335368 137428 335374
rect 137376 335310 137428 335316
rect 137282 328672 137338 328681
rect 137282 328607 137338 328616
rect 136548 271856 136600 271862
rect 136548 271798 136600 271804
rect 136088 257372 136140 257378
rect 136088 257314 136140 257320
rect 135996 76560 136048 76566
rect 135996 76502 136048 76508
rect 137296 42090 137324 328607
rect 137388 256018 137416 335310
rect 137468 294636 137520 294642
rect 137468 294578 137520 294584
rect 137480 278769 137508 294578
rect 137466 278760 137522 278769
rect 137466 278695 137522 278704
rect 137560 259548 137612 259554
rect 137560 259490 137612 259496
rect 137376 256012 137428 256018
rect 137376 255954 137428 255960
rect 137468 249076 137520 249082
rect 137468 249018 137520 249024
rect 137376 195288 137428 195294
rect 137376 195230 137428 195236
rect 137284 42084 137336 42090
rect 137284 42026 137336 42032
rect 137388 14482 137416 195230
rect 137480 193866 137508 249018
rect 137572 226302 137600 259490
rect 137848 234530 137876 392527
rect 137940 333441 137968 610030
rect 140688 608660 140740 608666
rect 140688 608602 140740 608608
rect 139308 507136 139360 507142
rect 139308 507078 139360 507084
rect 138020 445732 138072 445738
rect 138020 445674 138072 445680
rect 138032 445058 138060 445674
rect 138020 445052 138072 445058
rect 138020 444994 138072 445000
rect 137926 333432 137982 333441
rect 137926 333367 137982 333376
rect 138032 307766 138060 444994
rect 139320 429894 139348 507078
rect 140594 489968 140650 489977
rect 140594 489903 140650 489912
rect 139308 429888 139360 429894
rect 139308 429830 139360 429836
rect 140044 396772 140096 396778
rect 140044 396714 140096 396720
rect 140056 386374 140084 396714
rect 140044 386368 140096 386374
rect 139398 386336 139454 386345
rect 140044 386310 140096 386316
rect 139398 386271 139454 386280
rect 139412 385694 139440 386271
rect 139400 385688 139452 385694
rect 139400 385630 139452 385636
rect 140608 321473 140636 489903
rect 140700 408474 140728 608602
rect 142804 605872 142856 605878
rect 142804 605814 142856 605820
rect 141424 600432 141476 600438
rect 141424 600374 141476 600380
rect 140688 408468 140740 408474
rect 140688 408410 140740 408416
rect 141436 389298 141464 600374
rect 142620 593428 142672 593434
rect 142620 593370 142672 593376
rect 142632 593337 142660 593370
rect 142618 593328 142674 593337
rect 142618 593263 142674 593272
rect 141976 518220 142028 518226
rect 141976 518162 142028 518168
rect 141424 389292 141476 389298
rect 141424 389234 141476 389240
rect 141436 380186 141464 389234
rect 141988 384985 142016 518162
rect 142068 500268 142120 500274
rect 142068 500210 142120 500216
rect 141974 384976 142030 384985
rect 141974 384911 142030 384920
rect 141988 384441 142016 384911
rect 141974 384432 142030 384441
rect 141974 384367 142030 384376
rect 141424 380180 141476 380186
rect 141424 380122 141476 380128
rect 141516 374672 141568 374678
rect 141516 374614 141568 374620
rect 140780 361548 140832 361554
rect 140780 361490 140832 361496
rect 140792 360874 140820 361490
rect 140780 360868 140832 360874
rect 140780 360810 140832 360816
rect 140594 321464 140650 321473
rect 140594 321399 140650 321408
rect 140042 313304 140098 313313
rect 140042 313239 140098 313248
rect 138662 307864 138718 307873
rect 138662 307799 138718 307808
rect 138020 307760 138072 307766
rect 138020 307702 138072 307708
rect 138032 307086 138060 307702
rect 138020 307080 138072 307086
rect 138020 307022 138072 307028
rect 138676 294545 138704 307799
rect 138756 298784 138808 298790
rect 138756 298726 138808 298732
rect 138662 294536 138718 294545
rect 138662 294471 138718 294480
rect 138664 278044 138716 278050
rect 138664 277986 138716 277992
rect 137836 234524 137888 234530
rect 137836 234466 137888 234472
rect 137848 233889 137876 234466
rect 137834 233880 137890 233889
rect 137834 233815 137890 233824
rect 138676 227633 138704 277986
rect 138662 227624 138718 227633
rect 138662 227559 138718 227568
rect 137560 226296 137612 226302
rect 137560 226238 137612 226244
rect 137468 193860 137520 193866
rect 137468 193802 137520 193808
rect 138664 193860 138716 193866
rect 138664 193802 138716 193808
rect 137468 172644 137520 172650
rect 137468 172586 137520 172592
rect 137480 135250 137508 172586
rect 137468 135244 137520 135250
rect 137468 135186 137520 135192
rect 137376 14476 137428 14482
rect 137376 14418 137428 14424
rect 135904 11756 135956 11762
rect 135904 11698 135956 11704
rect 138676 10334 138704 193802
rect 138768 185638 138796 298726
rect 138756 185632 138808 185638
rect 138756 185574 138808 185580
rect 140056 13122 140084 313239
rect 141422 304192 141478 304201
rect 141422 304127 141478 304136
rect 140228 300144 140280 300150
rect 140228 300086 140280 300092
rect 140134 262848 140190 262857
rect 140134 262783 140190 262792
rect 140148 180130 140176 262783
rect 140240 261497 140268 300086
rect 140226 261488 140282 261497
rect 140226 261423 140282 261432
rect 140872 231804 140924 231810
rect 140872 231746 140924 231752
rect 140884 231130 140912 231746
rect 140872 231124 140924 231130
rect 140872 231066 140924 231072
rect 140136 180124 140188 180130
rect 140136 180066 140188 180072
rect 140134 160168 140190 160177
rect 140134 160103 140190 160112
rect 140148 128314 140176 160103
rect 140136 128308 140188 128314
rect 140136 128250 140188 128256
rect 140044 13116 140096 13122
rect 140044 13058 140096 13064
rect 138664 10328 138716 10334
rect 138664 10270 138716 10276
rect 141436 7682 141464 304127
rect 141528 231810 141556 374614
rect 142080 360874 142108 500210
rect 142160 450696 142212 450702
rect 142160 450638 142212 450644
rect 142068 360868 142120 360874
rect 142068 360810 142120 360816
rect 141608 332648 141660 332654
rect 141608 332590 141660 332596
rect 141620 262585 141648 332590
rect 141700 331900 141752 331906
rect 141700 331842 141752 331848
rect 141712 300218 141740 331842
rect 142172 312594 142200 450638
rect 142816 375329 142844 605814
rect 147600 600250 147628 614178
rect 152556 611448 152608 611454
rect 152556 611390 152608 611396
rect 147600 600222 147720 600250
rect 147692 599622 147720 600222
rect 147680 599616 147732 599622
rect 147680 599558 147732 599564
rect 146944 596284 146996 596290
rect 146944 596226 146996 596232
rect 143446 593328 143502 593337
rect 143446 593263 143502 593272
rect 143356 504416 143408 504422
rect 143356 504358 143408 504364
rect 142896 488572 142948 488578
rect 142896 488514 142948 488520
rect 142908 458862 142936 488514
rect 142896 458856 142948 458862
rect 142896 458798 142948 458804
rect 142988 458244 143040 458250
rect 142988 458186 143040 458192
rect 143000 450702 143028 458186
rect 142988 450696 143040 450702
rect 142988 450638 143040 450644
rect 143262 433256 143318 433265
rect 143262 433191 143318 433200
rect 142250 375320 142306 375329
rect 142250 375255 142306 375264
rect 142802 375320 142858 375329
rect 142802 375255 142858 375264
rect 142264 374678 142292 375255
rect 142252 374672 142304 374678
rect 142252 374614 142304 374620
rect 143276 347721 143304 433191
rect 143368 429321 143396 504358
rect 143460 488578 143488 593263
rect 146956 541686 146984 596226
rect 147496 585812 147548 585818
rect 147496 585754 147548 585760
rect 146944 541680 146996 541686
rect 146944 541622 146996 541628
rect 143632 537532 143684 537538
rect 143632 537474 143684 537480
rect 143644 537441 143672 537474
rect 143630 537432 143686 537441
rect 143630 537367 143686 537376
rect 143644 528554 143672 537367
rect 143552 528526 143672 528554
rect 143448 488572 143500 488578
rect 143448 488514 143500 488520
rect 143354 429312 143410 429321
rect 143354 429247 143410 429256
rect 143448 420980 143500 420986
rect 143448 420922 143500 420928
rect 142802 347712 142858 347721
rect 142802 347647 142858 347656
rect 143262 347712 143318 347721
rect 143262 347647 143318 347656
rect 142816 347041 142844 347647
rect 142802 347032 142858 347041
rect 142802 346967 142858 346976
rect 142894 326360 142950 326369
rect 142894 326295 142950 326304
rect 142160 312588 142212 312594
rect 142160 312530 142212 312536
rect 142802 301744 142858 301753
rect 142802 301679 142858 301688
rect 141700 300212 141752 300218
rect 141700 300154 141752 300160
rect 141700 272536 141752 272542
rect 141700 272478 141752 272484
rect 141606 262576 141662 262585
rect 141606 262511 141662 262520
rect 141712 242894 141740 272478
rect 141700 242888 141752 242894
rect 141700 242830 141752 242836
rect 141516 231804 141568 231810
rect 141516 231746 141568 231752
rect 141424 7676 141476 7682
rect 141424 7618 141476 7624
rect 134524 4208 134576 4214
rect 134524 4150 134576 4156
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 136468 480 136496 4150
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140056 480 140084 3470
rect 142816 3466 142844 301679
rect 142908 46238 142936 326295
rect 143460 282849 143488 420922
rect 143552 400926 143580 528526
rect 145562 527776 145618 527785
rect 145562 527711 145618 527720
rect 144828 519580 144880 519586
rect 144828 519522 144880 519528
rect 144736 484424 144788 484430
rect 144736 484366 144788 484372
rect 144184 455524 144236 455530
rect 144184 455466 144236 455472
rect 144196 415410 144224 455466
rect 144184 415404 144236 415410
rect 144184 415346 144236 415352
rect 144642 413944 144698 413953
rect 144642 413879 144698 413888
rect 143540 400920 143592 400926
rect 143540 400862 143592 400868
rect 144184 392624 144236 392630
rect 144184 392566 144236 392572
rect 144196 365634 144224 392566
rect 144184 365628 144236 365634
rect 144184 365570 144236 365576
rect 144182 326496 144238 326505
rect 144182 326431 144238 326440
rect 144196 304366 144224 326431
rect 144274 314800 144330 314809
rect 144274 314735 144330 314744
rect 144288 305658 144316 314735
rect 144276 305652 144328 305658
rect 144276 305594 144328 305600
rect 144184 304360 144236 304366
rect 144184 304302 144236 304308
rect 144184 286340 144236 286346
rect 144184 286282 144236 286288
rect 143446 282840 143502 282849
rect 143446 282775 143502 282784
rect 143460 282169 143488 282775
rect 143446 282160 143502 282169
rect 143446 282095 143502 282104
rect 142986 280528 143042 280537
rect 142986 280463 143042 280472
rect 143000 210526 143028 280463
rect 142988 210520 143040 210526
rect 142988 210462 143040 210468
rect 142986 169824 143042 169833
rect 142986 169759 143042 169768
rect 143000 132462 143028 169759
rect 142988 132456 143040 132462
rect 142988 132398 143040 132404
rect 144196 118017 144224 286282
rect 144656 238649 144684 413879
rect 144748 294642 144776 484366
rect 144840 376553 144868 519522
rect 145576 392601 145604 527711
rect 145656 514072 145708 514078
rect 145656 514014 145708 514020
rect 145668 432614 145696 514014
rect 146944 480276 146996 480282
rect 146944 480218 146996 480224
rect 146206 463720 146262 463729
rect 146206 463655 146262 463664
rect 145656 432608 145708 432614
rect 145656 432550 145708 432556
rect 145668 398138 145696 432550
rect 145656 398132 145708 398138
rect 145656 398074 145708 398080
rect 145562 392592 145618 392601
rect 145562 392527 145618 392536
rect 145656 392012 145708 392018
rect 145656 391954 145708 391960
rect 144826 376544 144882 376553
rect 144826 376479 144882 376488
rect 145668 358766 145696 391954
rect 145656 358760 145708 358766
rect 145656 358702 145708 358708
rect 145564 307080 145616 307086
rect 145564 307022 145616 307028
rect 144828 305040 144880 305046
rect 144828 304982 144880 304988
rect 144736 294636 144788 294642
rect 144736 294578 144788 294584
rect 144642 238640 144698 238649
rect 144642 238575 144698 238584
rect 144656 238105 144684 238575
rect 144642 238096 144698 238105
rect 144642 238031 144698 238040
rect 144182 118008 144238 118017
rect 144182 117943 144238 117952
rect 142896 46232 142948 46238
rect 142896 46174 142948 46180
rect 144840 3534 144868 304982
rect 145576 296177 145604 307022
rect 145654 305688 145710 305697
rect 145654 305623 145710 305632
rect 145562 296168 145618 296177
rect 145562 296103 145618 296112
rect 145576 295361 145604 296103
rect 145562 295352 145618 295361
rect 145562 295287 145618 295296
rect 145562 271280 145618 271289
rect 145562 271215 145618 271224
rect 145576 193934 145604 271215
rect 145564 193928 145616 193934
rect 145564 193870 145616 193876
rect 145564 185020 145616 185026
rect 145564 184962 145616 184968
rect 145576 35222 145604 184962
rect 145668 178702 145696 305623
rect 146220 267714 146248 463655
rect 146956 434722 146984 480218
rect 147036 437504 147088 437510
rect 147036 437446 147088 437452
rect 146944 434716 146996 434722
rect 146944 434658 146996 434664
rect 147048 411942 147076 437446
rect 147036 411936 147088 411942
rect 147036 411878 147088 411884
rect 147508 398206 147536 585754
rect 147586 454064 147642 454073
rect 147586 453999 147642 454008
rect 147496 398200 147548 398206
rect 147496 398142 147548 398148
rect 147496 372632 147548 372638
rect 147496 372574 147548 372580
rect 147508 353258 147536 372574
rect 147496 353252 147548 353258
rect 147496 353194 147548 353200
rect 146944 348492 146996 348498
rect 146944 348434 146996 348440
rect 146208 267708 146260 267714
rect 146208 267650 146260 267656
rect 146220 267102 146248 267650
rect 146208 267096 146260 267102
rect 146208 267038 146260 267044
rect 145656 178696 145708 178702
rect 145656 178638 145708 178644
rect 145654 156088 145710 156097
rect 145654 156023 145710 156032
rect 145668 121378 145696 156023
rect 145656 121372 145708 121378
rect 145656 121314 145708 121320
rect 146956 50386 146984 348434
rect 147128 346452 147180 346458
rect 147128 346394 147180 346400
rect 147140 311166 147168 346394
rect 147218 313984 147274 313993
rect 147218 313919 147274 313928
rect 147128 311160 147180 311166
rect 147128 311102 147180 311108
rect 147034 310720 147090 310729
rect 147034 310655 147090 310664
rect 146944 50380 146996 50386
rect 146944 50322 146996 50328
rect 147048 47598 147076 310655
rect 147232 304298 147260 313919
rect 147220 304292 147272 304298
rect 147220 304234 147272 304240
rect 147126 265568 147182 265577
rect 147126 265503 147182 265512
rect 147140 185706 147168 265503
rect 147128 185700 147180 185706
rect 147128 185642 147180 185648
rect 147036 47592 147088 47598
rect 147036 47534 147088 47540
rect 145564 35216 145616 35222
rect 145564 35158 145616 35164
rect 147600 3534 147628 453999
rect 147692 372638 147720 599558
rect 150164 597644 150216 597650
rect 150164 597586 150216 597592
rect 148968 578264 149020 578270
rect 148968 578206 149020 578212
rect 148324 472116 148376 472122
rect 148324 472058 148376 472064
rect 147772 449200 147824 449206
rect 147772 449142 147824 449148
rect 147784 448662 147812 449142
rect 147772 448656 147824 448662
rect 147772 448598 147824 448604
rect 148336 446486 148364 472058
rect 148876 449200 148928 449206
rect 148876 449142 148928 449148
rect 148324 446480 148376 446486
rect 148324 446422 148376 446428
rect 148324 435396 148376 435402
rect 148324 435338 148376 435344
rect 148336 423638 148364 435338
rect 148324 423632 148376 423638
rect 148324 423574 148376 423580
rect 148888 417450 148916 449142
rect 148876 417444 148928 417450
rect 148876 417386 148928 417392
rect 148324 403028 148376 403034
rect 148324 402970 148376 402976
rect 148336 374678 148364 402970
rect 148980 400217 149008 578206
rect 150176 469878 150204 597586
rect 151728 583024 151780 583030
rect 151728 582966 151780 582972
rect 150256 565140 150308 565146
rect 150256 565082 150308 565088
rect 150164 469872 150216 469878
rect 150164 469814 150216 469820
rect 149704 466540 149756 466546
rect 149704 466482 149756 466488
rect 149060 416152 149112 416158
rect 149060 416094 149112 416100
rect 149072 415478 149100 416094
rect 149060 415472 149112 415478
rect 149060 415414 149112 415420
rect 148966 400208 149022 400217
rect 148966 400143 149022 400152
rect 148980 399498 149008 400143
rect 148968 399492 149020 399498
rect 148968 399434 149020 399440
rect 148416 392692 148468 392698
rect 148416 392634 148468 392640
rect 148428 378146 148456 392634
rect 148416 378140 148468 378146
rect 148416 378082 148468 378088
rect 148324 374672 148376 374678
rect 148324 374614 148376 374620
rect 147680 372632 147732 372638
rect 147680 372574 147732 372580
rect 148506 338872 148562 338881
rect 148506 338807 148562 338816
rect 148416 311908 148468 311914
rect 148416 311850 148468 311856
rect 148324 303680 148376 303686
rect 148324 303622 148376 303628
rect 148336 21418 148364 303622
rect 148428 129130 148456 311850
rect 148520 193866 148548 338807
rect 149716 318073 149744 466482
rect 149796 458312 149848 458318
rect 149796 458254 149848 458260
rect 149808 419490 149836 458254
rect 150268 433294 150296 565082
rect 150440 538892 150492 538898
rect 150440 538834 150492 538840
rect 150452 538286 150480 538834
rect 150440 538280 150492 538286
rect 150440 538222 150492 538228
rect 151636 538280 151688 538286
rect 151636 538222 151688 538228
rect 150346 515400 150402 515409
rect 150346 515335 150402 515344
rect 150256 433288 150308 433294
rect 150256 433230 150308 433236
rect 149796 419484 149848 419490
rect 149796 419426 149848 419432
rect 150256 416152 150308 416158
rect 150256 416094 150308 416100
rect 150268 369753 150296 416094
rect 150254 369744 150310 369753
rect 150254 369679 150310 369688
rect 150360 344350 150388 515335
rect 151648 476241 151676 538222
rect 151082 476232 151138 476241
rect 151082 476167 151138 476176
rect 151634 476232 151690 476241
rect 151634 476167 151690 476176
rect 150532 433288 150584 433294
rect 150532 433230 150584 433236
rect 150348 344344 150400 344350
rect 150348 344286 150400 344292
rect 150438 333432 150494 333441
rect 150438 333367 150494 333376
rect 150452 332625 150480 333367
rect 150438 332616 150494 332625
rect 150438 332551 150494 332560
rect 149794 328536 149850 328545
rect 149794 328471 149850 328480
rect 149702 318064 149758 318073
rect 149702 317999 149758 318008
rect 149716 311250 149744 317999
rect 149808 311370 149836 328471
rect 149980 317552 150032 317558
rect 149980 317494 150032 317500
rect 149796 311364 149848 311370
rect 149796 311306 149848 311312
rect 149716 311222 149836 311250
rect 149702 306640 149758 306649
rect 149702 306575 149758 306584
rect 148600 265668 148652 265674
rect 148600 265610 148652 265616
rect 148612 247722 148640 265610
rect 148600 247716 148652 247722
rect 148600 247658 148652 247664
rect 148508 193860 148560 193866
rect 148508 193802 148560 193808
rect 148600 149796 148652 149802
rect 148600 149738 148652 149744
rect 148508 133272 148560 133278
rect 148508 133214 148560 133220
rect 148416 129124 148468 129130
rect 148416 129066 148468 129072
rect 148324 21412 148376 21418
rect 148324 21354 148376 21360
rect 148520 3602 148548 133214
rect 148612 133210 148640 149738
rect 148600 133204 148652 133210
rect 148600 133146 148652 133152
rect 149716 4826 149744 306575
rect 149808 306374 149836 311222
rect 149992 307766 150020 317494
rect 149980 307760 150032 307766
rect 149980 307702 150032 307708
rect 149808 306346 149928 306374
rect 149794 271144 149850 271153
rect 149794 271079 149850 271088
rect 149808 212430 149836 271079
rect 149900 261526 149928 306346
rect 149888 261520 149940 261526
rect 149888 261462 149940 261468
rect 149796 212424 149848 212430
rect 149796 212366 149848 212372
rect 150452 195294 150480 332551
rect 150544 299441 150572 433230
rect 151096 433226 151124 476167
rect 151266 465760 151322 465769
rect 151266 465695 151322 465704
rect 151174 456104 151230 456113
rect 151174 456039 151230 456048
rect 151084 433220 151136 433226
rect 151084 433162 151136 433168
rect 151188 416090 151216 456039
rect 151280 429146 151308 465695
rect 151268 429140 151320 429146
rect 151268 429082 151320 429088
rect 151636 427100 151688 427106
rect 151636 427042 151688 427048
rect 151176 416084 151228 416090
rect 151176 416026 151228 416032
rect 151176 408536 151228 408542
rect 151176 408478 151228 408484
rect 151084 394800 151136 394806
rect 151084 394742 151136 394748
rect 151096 362234 151124 394742
rect 151188 376718 151216 408478
rect 151176 376712 151228 376718
rect 151176 376654 151228 376660
rect 151084 362228 151136 362234
rect 151084 362170 151136 362176
rect 151084 323672 151136 323678
rect 151084 323614 151136 323620
rect 150530 299432 150586 299441
rect 150530 299367 150586 299376
rect 150544 298761 150572 299367
rect 150530 298752 150586 298761
rect 150530 298687 150586 298696
rect 151096 289134 151124 323614
rect 151648 316810 151676 427042
rect 151740 409193 151768 582966
rect 152462 533352 152518 533361
rect 152462 533287 152518 533296
rect 151726 409184 151782 409193
rect 151726 409119 151782 409128
rect 151636 316804 151688 316810
rect 151636 316746 151688 316752
rect 151176 308440 151228 308446
rect 151176 308382 151228 308388
rect 151084 289128 151136 289134
rect 151084 289070 151136 289076
rect 151082 267064 151138 267073
rect 151082 266999 151138 267008
rect 150440 195288 150492 195294
rect 150440 195230 150492 195236
rect 150440 131776 150492 131782
rect 150440 131718 150492 131724
rect 150452 124166 150480 131718
rect 150440 124160 150492 124166
rect 150440 124102 150492 124108
rect 151096 19990 151124 266999
rect 151188 264217 151216 308382
rect 151360 291848 151412 291854
rect 151360 291790 151412 291796
rect 151268 276072 151320 276078
rect 151268 276014 151320 276020
rect 151174 264208 151230 264217
rect 151174 264143 151230 264152
rect 151174 258768 151230 258777
rect 151174 258703 151230 258712
rect 151188 54534 151216 258703
rect 151280 249150 151308 276014
rect 151372 270502 151400 291790
rect 151360 270496 151412 270502
rect 151360 270438 151412 270444
rect 151268 249144 151320 249150
rect 151268 249086 151320 249092
rect 151268 151904 151320 151910
rect 151268 151846 151320 151852
rect 151280 136241 151308 151846
rect 151360 137284 151412 137290
rect 151360 137226 151412 137232
rect 151266 136232 151322 136241
rect 151266 136167 151322 136176
rect 151372 129742 151400 137226
rect 151360 129736 151412 129742
rect 151360 129678 151412 129684
rect 151176 54528 151228 54534
rect 151176 54470 151228 54476
rect 151084 19984 151136 19990
rect 151084 19926 151136 19932
rect 149704 4820 149756 4826
rect 149704 4762 149756 4768
rect 152476 3670 152504 533287
rect 152568 461650 152596 611390
rect 154488 508564 154540 508570
rect 154488 508506 154540 508512
rect 153108 485104 153160 485110
rect 153108 485046 153160 485052
rect 152556 461644 152608 461650
rect 152556 461586 152608 461592
rect 152922 460184 152978 460193
rect 152922 460119 152978 460128
rect 152936 429146 152964 460119
rect 153016 445052 153068 445058
rect 153016 444994 153068 445000
rect 152924 429140 152976 429146
rect 152924 429082 152976 429088
rect 152924 405680 152976 405686
rect 152924 405622 152976 405628
rect 152936 378049 152964 405622
rect 152922 378040 152978 378049
rect 152922 377975 152978 377984
rect 152936 377369 152964 377975
rect 152922 377360 152978 377369
rect 152922 377295 152978 377304
rect 153028 329798 153056 444994
rect 153120 416090 153148 485046
rect 153934 466576 153990 466585
rect 153934 466511 153990 466520
rect 153844 459604 153896 459610
rect 153844 459546 153896 459552
rect 153856 419422 153884 459546
rect 153948 436801 153976 466511
rect 154396 450560 154448 450566
rect 154396 450502 154448 450508
rect 154408 447846 154436 450502
rect 154396 447840 154448 447846
rect 154396 447782 154448 447788
rect 154028 438932 154080 438938
rect 154028 438874 154080 438880
rect 153934 436792 153990 436801
rect 153934 436727 153990 436736
rect 154040 431254 154068 438874
rect 154028 431248 154080 431254
rect 154028 431190 154080 431196
rect 153844 419416 153896 419422
rect 153844 419358 153896 419364
rect 154394 417480 154450 417489
rect 154394 417415 154450 417424
rect 154408 416838 154436 417415
rect 154396 416832 154448 416838
rect 154396 416774 154448 416780
rect 153108 416084 153160 416090
rect 153108 416026 153160 416032
rect 153016 329792 153068 329798
rect 153016 329734 153068 329740
rect 152556 323604 152608 323610
rect 152556 323546 152608 323552
rect 152568 25566 152596 323546
rect 152646 285696 152702 285705
rect 152646 285631 152702 285640
rect 152660 229770 152688 285631
rect 152648 229764 152700 229770
rect 152648 229706 152700 229712
rect 153120 222154 153148 416026
rect 153844 404456 153896 404462
rect 153844 404398 153896 404404
rect 153856 361554 153884 404398
rect 154408 389881 154436 416774
rect 154500 406434 154528 508506
rect 155222 466576 155278 466585
rect 155222 466511 155278 466520
rect 155236 425066 155264 466511
rect 155316 429888 155368 429894
rect 155316 429830 155368 429836
rect 155224 425060 155276 425066
rect 155224 425002 155276 425008
rect 154488 406428 154540 406434
rect 154488 406370 154540 406376
rect 154500 405686 154528 406370
rect 154488 405680 154540 405686
rect 154488 405622 154540 405628
rect 155328 394670 155356 429830
rect 155604 420918 155632 615470
rect 160744 610020 160796 610026
rect 160744 609962 160796 609968
rect 157984 590708 158036 590714
rect 157984 590650 158036 590656
rect 157248 574116 157300 574122
rect 157248 574058 157300 574064
rect 156604 546576 156656 546582
rect 156604 546518 156656 546524
rect 155776 541748 155828 541754
rect 155776 541690 155828 541696
rect 155788 541006 155816 541690
rect 155776 541000 155828 541006
rect 155776 540942 155828 540948
rect 155684 498840 155736 498846
rect 155684 498782 155736 498788
rect 155696 440230 155724 498782
rect 155684 440224 155736 440230
rect 155684 440166 155736 440172
rect 155696 439521 155724 440166
rect 155682 439512 155738 439521
rect 155682 439447 155738 439456
rect 155788 431934 155816 540942
rect 155776 431928 155828 431934
rect 155776 431870 155828 431876
rect 155868 423632 155920 423638
rect 155868 423574 155920 423580
rect 155592 420912 155644 420918
rect 155592 420854 155644 420860
rect 155604 419665 155632 420854
rect 155590 419656 155646 419665
rect 155590 419591 155646 419600
rect 155776 409896 155828 409902
rect 155776 409838 155828 409844
rect 155316 394664 155368 394670
rect 155316 394606 155368 394612
rect 155682 390960 155738 390969
rect 155682 390895 155738 390904
rect 154488 389904 154540 389910
rect 154394 389872 154450 389881
rect 154488 389846 154540 389852
rect 154394 389807 154450 389816
rect 154500 378865 154528 389846
rect 155224 386504 155276 386510
rect 155224 386446 155276 386452
rect 154486 378856 154542 378865
rect 153936 378820 153988 378826
rect 154486 378791 154542 378800
rect 153936 378762 153988 378768
rect 153948 373386 153976 378762
rect 154500 376650 154528 378791
rect 154488 376644 154540 376650
rect 154488 376586 154540 376592
rect 153936 373380 153988 373386
rect 153936 373322 153988 373328
rect 153844 361548 153896 361554
rect 153844 361490 153896 361496
rect 155236 357377 155264 386446
rect 155696 371210 155724 390895
rect 155788 380225 155816 409838
rect 155774 380216 155830 380225
rect 155774 380151 155830 380160
rect 155684 371204 155736 371210
rect 155684 371146 155736 371152
rect 155222 357368 155278 357377
rect 155222 357303 155278 357312
rect 153844 353320 153896 353326
rect 153844 353262 153896 353268
rect 153856 347721 153884 353262
rect 153842 347712 153898 347721
rect 153842 347647 153898 347656
rect 155224 338768 155276 338774
rect 155224 338710 155276 338716
rect 153198 338056 153254 338065
rect 153198 337991 153254 338000
rect 153212 329118 153240 337991
rect 154026 334792 154082 334801
rect 154026 334727 154082 334736
rect 153200 329112 153252 329118
rect 153200 329054 153252 329060
rect 154040 326398 154068 334727
rect 154028 326392 154080 326398
rect 154028 326334 154080 326340
rect 153936 325032 153988 325038
rect 153936 324974 153988 324980
rect 153842 310448 153898 310457
rect 153842 310383 153898 310392
rect 153856 243574 153884 310383
rect 153948 279478 153976 324974
rect 154026 320784 154082 320793
rect 154026 320719 154082 320728
rect 153936 279472 153988 279478
rect 153936 279414 153988 279420
rect 153934 278080 153990 278089
rect 153934 278015 153990 278024
rect 153844 243568 153896 243574
rect 153844 243510 153896 243516
rect 153108 222148 153160 222154
rect 153108 222090 153160 222096
rect 153120 221474 153148 222090
rect 153108 221468 153160 221474
rect 153108 221410 153160 221416
rect 153844 218748 153896 218754
rect 153844 218690 153896 218696
rect 153856 208321 153884 218690
rect 153842 208312 153898 208321
rect 153842 208247 153898 208256
rect 153842 185600 153898 185609
rect 153842 185535 153898 185544
rect 152648 162988 152700 162994
rect 152648 162930 152700 162936
rect 152660 137873 152688 162930
rect 152646 137864 152702 137873
rect 152646 137799 152702 137808
rect 153856 53106 153884 185535
rect 153948 185026 153976 278015
rect 154040 276729 154068 320719
rect 154026 276720 154082 276729
rect 154026 276655 154082 276664
rect 155236 272610 155264 338710
rect 155316 325712 155368 325718
rect 155316 325654 155368 325660
rect 155224 272604 155276 272610
rect 155224 272546 155276 272552
rect 154026 268424 154082 268433
rect 154026 268359 154082 268368
rect 154040 218754 154068 268359
rect 155222 261488 155278 261497
rect 155222 261423 155278 261432
rect 154028 218748 154080 218754
rect 154028 218690 154080 218696
rect 153936 185020 153988 185026
rect 153936 184962 153988 184968
rect 153934 164384 153990 164393
rect 153934 164319 153990 164328
rect 154028 164348 154080 164354
rect 153948 146946 153976 164319
rect 154028 164290 154080 164296
rect 154040 158030 154068 164290
rect 154028 158024 154080 158030
rect 154028 157966 154080 157972
rect 154028 154692 154080 154698
rect 154028 154634 154080 154640
rect 154040 146946 154068 154634
rect 153936 146940 153988 146946
rect 153936 146882 153988 146888
rect 154028 146940 154080 146946
rect 154028 146882 154080 146888
rect 153934 144936 153990 144945
rect 153934 144871 153990 144880
rect 153948 122806 153976 144871
rect 153936 122800 153988 122806
rect 153936 122742 153988 122748
rect 153936 101448 153988 101454
rect 153936 101390 153988 101396
rect 153948 74458 153976 101390
rect 153936 74452 153988 74458
rect 153936 74394 153988 74400
rect 153844 53100 153896 53106
rect 153844 53042 153896 53048
rect 152556 25560 152608 25566
rect 152556 25502 152608 25508
rect 155236 18630 155264 261423
rect 155328 258738 155356 325654
rect 155880 321638 155908 423574
rect 155958 394768 156014 394777
rect 155958 394703 156014 394712
rect 155972 394670 156000 394703
rect 155960 394664 156012 394670
rect 155960 394606 156012 394612
rect 155972 367062 156000 394606
rect 156616 390969 156644 546518
rect 157154 481808 157210 481817
rect 157154 481743 157210 481752
rect 156602 390960 156658 390969
rect 156602 390895 156658 390904
rect 155960 367056 156012 367062
rect 155960 366998 156012 367004
rect 155972 364334 156000 366998
rect 155972 364306 156092 364334
rect 155868 321632 155920 321638
rect 155868 321574 155920 321580
rect 155408 310548 155460 310554
rect 155408 310490 155460 310496
rect 155420 275330 155448 310490
rect 155960 294704 156012 294710
rect 155960 294646 156012 294652
rect 155972 294030 156000 294646
rect 155960 294024 156012 294030
rect 155960 293966 156012 293972
rect 155500 281580 155552 281586
rect 155500 281522 155552 281528
rect 155408 275324 155460 275330
rect 155408 275266 155460 275272
rect 155512 263566 155540 281522
rect 155500 263560 155552 263566
rect 155500 263502 155552 263508
rect 155406 260128 155462 260137
rect 155406 260063 155462 260072
rect 155316 258732 155368 258738
rect 155316 258674 155368 258680
rect 155314 233200 155370 233209
rect 155314 233135 155370 233144
rect 155328 36582 155356 233135
rect 155420 226953 155448 260063
rect 155406 226944 155462 226953
rect 155406 226879 155462 226888
rect 155406 153776 155462 153785
rect 155406 153711 155462 153720
rect 155420 125594 155448 153711
rect 155972 138009 156000 293966
rect 156064 242185 156092 364306
rect 156604 300824 156656 300830
rect 156604 300766 156656 300772
rect 156616 294710 156644 300766
rect 156604 294704 156656 294710
rect 156604 294646 156656 294652
rect 157168 292534 157196 481743
rect 157260 308446 157288 574058
rect 157996 394738 158024 590650
rect 159364 580304 159416 580310
rect 159364 580246 159416 580252
rect 159376 579698 159404 580246
rect 159364 579692 159416 579698
rect 159364 579634 159416 579640
rect 158812 542428 158864 542434
rect 158812 542370 158864 542376
rect 158444 516792 158496 516798
rect 158444 516734 158496 516740
rect 157984 394732 158036 394738
rect 157984 394674 158036 394680
rect 157340 373312 157392 373318
rect 157340 373254 157392 373260
rect 157352 367062 157380 373254
rect 157996 368393 158024 394674
rect 158456 390697 158484 516734
rect 158626 498808 158682 498817
rect 158626 498743 158682 498752
rect 158534 461544 158590 461553
rect 158534 461479 158590 461488
rect 158442 390688 158498 390697
rect 158442 390623 158498 390632
rect 158456 390590 158484 390623
rect 158444 390584 158496 390590
rect 158444 390526 158496 390532
rect 157982 368384 158038 368393
rect 157982 368319 158038 368328
rect 157340 367056 157392 367062
rect 157340 366998 157392 367004
rect 158444 367056 158496 367062
rect 158444 366998 158496 367004
rect 157340 329792 157392 329798
rect 157340 329734 157392 329740
rect 157352 328506 157380 329734
rect 157340 328500 157392 328506
rect 157340 328442 157392 328448
rect 157248 308440 157300 308446
rect 157248 308382 157300 308388
rect 157156 292528 157208 292534
rect 157156 292470 157208 292476
rect 156696 273284 156748 273290
rect 156696 273226 156748 273232
rect 156602 251968 156658 251977
rect 156602 251903 156658 251912
rect 156050 242176 156106 242185
rect 156050 242111 156106 242120
rect 155958 138000 156014 138009
rect 155958 137935 156014 137944
rect 156418 138000 156474 138009
rect 156418 137935 156474 137944
rect 156432 137329 156460 137935
rect 156418 137320 156474 137329
rect 156418 137255 156474 137264
rect 155408 125588 155460 125594
rect 155408 125530 155460 125536
rect 155868 125588 155920 125594
rect 155868 125530 155920 125536
rect 155880 124234 155908 125530
rect 155868 124228 155920 124234
rect 155868 124170 155920 124176
rect 155880 101454 155908 124170
rect 155868 101448 155920 101454
rect 155868 101390 155920 101396
rect 156616 40730 156644 251903
rect 156708 125594 156736 273226
rect 157352 160721 157380 328442
rect 158456 278050 158484 366998
rect 158548 303521 158576 461479
rect 158640 338745 158668 498743
rect 158720 471300 158772 471306
rect 158720 471242 158772 471248
rect 158732 471209 158760 471242
rect 158718 471200 158774 471209
rect 158718 471135 158774 471144
rect 158720 445732 158772 445738
rect 158720 445674 158772 445680
rect 158732 444446 158760 445674
rect 158720 444440 158772 444446
rect 158720 444382 158772 444388
rect 158626 338736 158682 338745
rect 158626 338671 158682 338680
rect 158534 303512 158590 303521
rect 158534 303447 158590 303456
rect 158732 283014 158760 444382
rect 158824 434858 158852 542370
rect 159376 471209 159404 579634
rect 160756 576842 160784 609962
rect 160834 581088 160890 581097
rect 160834 581023 160890 581032
rect 160744 576836 160796 576842
rect 160744 576778 160796 576784
rect 160100 570648 160152 570654
rect 160100 570590 160152 570596
rect 160112 569974 160140 570590
rect 160100 569968 160152 569974
rect 160100 569910 160152 569916
rect 159916 557592 159968 557598
rect 159916 557534 159968 557540
rect 159362 471200 159418 471209
rect 159362 471135 159418 471144
rect 159364 463752 159416 463758
rect 159364 463694 159416 463700
rect 159376 445738 159404 463694
rect 159364 445732 159416 445738
rect 159364 445674 159416 445680
rect 158812 434852 158864 434858
rect 158812 434794 158864 434800
rect 158824 423638 158852 434794
rect 158812 423632 158864 423638
rect 158812 423574 158864 423580
rect 158812 411936 158864 411942
rect 158812 411878 158864 411884
rect 158824 411330 158852 411878
rect 158812 411324 158864 411330
rect 158812 411266 158864 411272
rect 159364 411324 159416 411330
rect 159364 411266 159416 411272
rect 158812 321632 158864 321638
rect 158812 321574 158864 321580
rect 158824 287774 158852 321574
rect 159376 316742 159404 411266
rect 159928 407794 159956 557534
rect 160008 486464 160060 486470
rect 160008 486406 160060 486412
rect 159916 407788 159968 407794
rect 159916 407730 159968 407736
rect 159364 316736 159416 316742
rect 159364 316678 159416 316684
rect 160020 301617 160048 486406
rect 160112 409902 160140 569910
rect 160848 556850 160876 581023
rect 160836 556844 160888 556850
rect 160836 556786 160888 556792
rect 160192 551336 160244 551342
rect 160192 551278 160244 551284
rect 160204 550662 160232 551278
rect 160192 550656 160244 550662
rect 160192 550598 160244 550604
rect 160744 550656 160796 550662
rect 160744 550598 160796 550604
rect 160100 409896 160152 409902
rect 160100 409838 160152 409844
rect 160100 393304 160152 393310
rect 160100 393246 160152 393252
rect 160112 392630 160140 393246
rect 160100 392624 160152 392630
rect 160100 392566 160152 392572
rect 160756 389842 160784 550598
rect 160836 452668 160888 452674
rect 160836 452610 160888 452616
rect 160100 389836 160152 389842
rect 160100 389778 160152 389784
rect 160744 389836 160796 389842
rect 160744 389778 160796 389784
rect 160112 389230 160140 389778
rect 160100 389224 160152 389230
rect 160100 389166 160152 389172
rect 160742 382936 160798 382945
rect 160742 382871 160798 382880
rect 160756 371142 160784 382871
rect 160744 371136 160796 371142
rect 160744 371078 160796 371084
rect 160756 370326 160784 371078
rect 160100 370320 160152 370326
rect 160100 370262 160152 370268
rect 160744 370320 160796 370326
rect 160744 370262 160796 370268
rect 160006 301608 160062 301617
rect 160006 301543 160062 301552
rect 159548 298852 159600 298858
rect 159548 298794 159600 298800
rect 159456 289128 159508 289134
rect 159456 289070 159508 289076
rect 159468 288454 159496 289070
rect 159456 288448 159508 288454
rect 159456 288390 159508 288396
rect 158812 287768 158864 287774
rect 158812 287710 158864 287716
rect 158720 283008 158772 283014
rect 158720 282950 158772 282956
rect 158732 278798 158760 282950
rect 158720 278792 158772 278798
rect 158720 278734 158772 278740
rect 158444 278044 158496 278050
rect 158444 277986 158496 277992
rect 157982 274816 158038 274825
rect 157982 274751 158038 274760
rect 157338 160712 157394 160721
rect 157338 160647 157394 160656
rect 157352 160313 157380 160647
rect 157338 160304 157394 160313
rect 157338 160239 157394 160248
rect 156696 125588 156748 125594
rect 156696 125530 156748 125536
rect 156604 40724 156656 40730
rect 156604 40666 156656 40672
rect 155316 36576 155368 36582
rect 155316 36518 155368 36524
rect 157996 29714 158024 274751
rect 158628 271788 158680 271794
rect 158628 271730 158680 271736
rect 158074 160304 158130 160313
rect 158074 160239 158130 160248
rect 158088 127634 158116 160239
rect 158076 127628 158128 127634
rect 158076 127570 158128 127576
rect 158640 93906 158668 271730
rect 159362 246256 159418 246265
rect 159362 246191 159418 246200
rect 158720 154692 158772 154698
rect 158720 154634 158772 154640
rect 158732 153882 158760 154634
rect 158720 153876 158772 153882
rect 158720 153818 158772 153824
rect 158628 93900 158680 93906
rect 158628 93842 158680 93848
rect 158640 92177 158668 93842
rect 158626 92168 158682 92177
rect 158626 92103 158682 92112
rect 159376 39370 159404 246191
rect 159468 141438 159496 288390
rect 159560 246362 159588 298794
rect 160112 281489 160140 370262
rect 160744 314764 160796 314770
rect 160744 314706 160796 314712
rect 160282 282976 160338 282985
rect 160282 282911 160338 282920
rect 160098 281480 160154 281489
rect 160098 281415 160154 281424
rect 160112 280809 160140 281415
rect 160098 280800 160154 280809
rect 160098 280735 160154 280744
rect 160192 278792 160244 278798
rect 160192 278734 160244 278740
rect 160100 271856 160152 271862
rect 160100 271798 160152 271804
rect 159640 269816 159692 269822
rect 159640 269758 159692 269764
rect 159652 248414 159680 269758
rect 159652 248386 160048 248414
rect 159548 246356 159600 246362
rect 159548 246298 159600 246304
rect 160020 238746 160048 248386
rect 160008 238740 160060 238746
rect 160008 238682 160060 238688
rect 159548 215960 159600 215966
rect 159548 215902 159600 215908
rect 159560 204270 159588 215902
rect 159548 204264 159600 204270
rect 159548 204206 159600 204212
rect 159560 145081 159588 204206
rect 160020 154698 160048 238682
rect 160008 154692 160060 154698
rect 160008 154634 160060 154640
rect 159546 145072 159602 145081
rect 159546 145007 159602 145016
rect 159456 141432 159508 141438
rect 159456 141374 159508 141380
rect 159456 135992 159508 135998
rect 159456 135934 159508 135940
rect 159364 39364 159416 39370
rect 159364 39306 159416 39312
rect 157984 29708 158036 29714
rect 157984 29650 158036 29656
rect 155224 18624 155276 18630
rect 155224 18566 155276 18572
rect 159468 13190 159496 135934
rect 159560 121378 159588 145007
rect 159548 121372 159600 121378
rect 159548 121314 159600 121320
rect 160112 37942 160140 271798
rect 160204 151842 160232 278734
rect 160296 249082 160324 282911
rect 160756 274650 160784 314706
rect 160848 300830 160876 452610
rect 161400 393310 161428 616830
rect 162124 592068 162176 592074
rect 162124 592010 162176 592016
rect 161480 394732 161532 394738
rect 161480 394674 161532 394680
rect 161388 393304 161440 393310
rect 161388 393246 161440 393252
rect 161492 392698 161520 394674
rect 161480 392692 161532 392698
rect 161480 392634 161532 392640
rect 162136 384305 162164 592010
rect 164056 559564 164108 559570
rect 164056 559506 164108 559512
rect 162216 554804 162268 554810
rect 162216 554746 162268 554752
rect 162228 522986 162256 554746
rect 162308 549908 162360 549914
rect 162308 549850 162360 549856
rect 162320 549302 162348 549850
rect 162308 549296 162360 549302
rect 162308 549238 162360 549244
rect 162216 522980 162268 522986
rect 162216 522922 162268 522928
rect 162228 404394 162256 522922
rect 162320 465050 162348 549238
rect 162676 496120 162728 496126
rect 162676 496062 162728 496068
rect 162308 465044 162360 465050
rect 162308 464986 162360 464992
rect 162216 404388 162268 404394
rect 162216 404330 162268 404336
rect 162584 404388 162636 404394
rect 162584 404330 162636 404336
rect 162596 403646 162624 404330
rect 162584 403640 162636 403646
rect 162584 403582 162636 403588
rect 162582 401704 162638 401713
rect 162582 401639 162638 401648
rect 162216 392012 162268 392018
rect 162216 391954 162268 391960
rect 162122 384296 162178 384305
rect 162122 384231 162178 384240
rect 161294 383752 161350 383761
rect 161294 383687 161350 383696
rect 161308 378146 161336 383687
rect 161388 381540 161440 381546
rect 161388 381482 161440 381488
rect 161296 378140 161348 378146
rect 161296 378082 161348 378088
rect 160836 300824 160888 300830
rect 160836 300766 160888 300772
rect 161400 280838 161428 381482
rect 162228 380866 162256 391954
rect 161480 380860 161532 380866
rect 161480 380802 161532 380808
rect 162216 380860 162268 380866
rect 162216 380802 162268 380808
rect 160836 280832 160888 280838
rect 160836 280774 160888 280780
rect 161388 280832 161440 280838
rect 161388 280774 161440 280780
rect 160744 274644 160796 274650
rect 160744 274586 160796 274592
rect 160848 273290 160876 280774
rect 160836 273284 160888 273290
rect 160836 273226 160888 273232
rect 161492 271794 161520 380802
rect 162122 377360 162178 377369
rect 162122 377295 162178 377304
rect 162136 327185 162164 377295
rect 162596 351218 162624 401639
rect 162688 394738 162716 496062
rect 163964 493332 164016 493338
rect 163964 493274 164016 493280
rect 163502 483712 163558 483721
rect 163502 483647 163558 483656
rect 162768 465044 162820 465050
rect 162768 464986 162820 464992
rect 162780 464370 162808 464986
rect 162768 464364 162820 464370
rect 162768 464306 162820 464312
rect 162768 457496 162820 457502
rect 162768 457438 162820 457444
rect 162676 394732 162728 394738
rect 162676 394674 162728 394680
rect 162584 351212 162636 351218
rect 162584 351154 162636 351160
rect 162122 327176 162178 327185
rect 162122 327111 162178 327120
rect 162136 323678 162164 327111
rect 162124 323672 162176 323678
rect 162124 323614 162176 323620
rect 162124 318844 162176 318850
rect 162124 318786 162176 318792
rect 161940 295996 161992 296002
rect 161940 295938 161992 295944
rect 161952 290494 161980 295938
rect 161940 290488 161992 290494
rect 161940 290430 161992 290436
rect 162136 284889 162164 318786
rect 162216 289876 162268 289882
rect 162216 289818 162268 289824
rect 162122 284880 162178 284889
rect 162122 284815 162178 284824
rect 161480 271788 161532 271794
rect 161480 271730 161532 271736
rect 162124 270496 162176 270502
rect 162124 270438 162176 270444
rect 161480 253904 161532 253910
rect 161480 253846 161532 253852
rect 160284 249076 160336 249082
rect 160284 249018 160336 249024
rect 160744 224256 160796 224262
rect 160744 224198 160796 224204
rect 160756 219434 160784 224198
rect 160744 219428 160796 219434
rect 160744 219370 160796 219376
rect 161388 219428 161440 219434
rect 161388 219370 161440 219376
rect 160192 151836 160244 151842
rect 160192 151778 160244 151784
rect 160744 151836 160796 151842
rect 160744 151778 160796 151784
rect 160190 136096 160246 136105
rect 160190 136031 160246 136040
rect 160204 135930 160232 136031
rect 160192 135924 160244 135930
rect 160192 135866 160244 135872
rect 160756 124166 160784 151778
rect 161400 135930 161428 219370
rect 161388 135924 161440 135930
rect 161388 135866 161440 135872
rect 160836 129056 160888 129062
rect 160836 128998 160888 129004
rect 160744 124160 160796 124166
rect 160744 124102 160796 124108
rect 160744 117360 160796 117366
rect 160744 117302 160796 117308
rect 160756 70310 160784 117302
rect 160848 106282 160876 128998
rect 160836 106276 160888 106282
rect 160836 106218 160888 106224
rect 160744 70304 160796 70310
rect 160744 70246 160796 70252
rect 160100 37936 160152 37942
rect 160100 37878 160152 37884
rect 161492 22778 161520 253846
rect 162136 28286 162164 270438
rect 162228 254590 162256 289818
rect 162780 289814 162808 457438
rect 163516 401713 163544 483647
rect 163502 401704 163558 401713
rect 163502 401639 163558 401648
rect 163976 397458 164004 493274
rect 164068 404326 164096 559506
rect 164056 404320 164108 404326
rect 164056 404262 164108 404268
rect 163504 397452 163556 397458
rect 163504 397394 163556 397400
rect 163964 397452 164016 397458
rect 163964 397394 164016 397400
rect 163516 396098 163544 397394
rect 163504 396092 163556 396098
rect 163504 396034 163556 396040
rect 163516 386510 163544 396034
rect 164056 395004 164108 395010
rect 164056 394946 164108 394952
rect 163596 390584 163648 390590
rect 163596 390526 163648 390532
rect 163504 386504 163556 386510
rect 163504 386446 163556 386452
rect 163504 385756 163556 385762
rect 163504 385698 163556 385704
rect 163516 373998 163544 385698
rect 163504 373992 163556 373998
rect 163504 373934 163556 373940
rect 163504 331288 163556 331294
rect 163504 331230 163556 331236
rect 162768 289808 162820 289814
rect 162768 289750 162820 289756
rect 162780 289134 162808 289750
rect 162768 289128 162820 289134
rect 162768 289070 162820 289076
rect 162768 283620 162820 283626
rect 162768 283562 162820 283568
rect 162780 282946 162808 283562
rect 162768 282940 162820 282946
rect 162768 282882 162820 282888
rect 162780 277394 162808 282882
rect 162688 277366 162808 277394
rect 162216 254584 162268 254590
rect 162216 254526 162268 254532
rect 162688 194546 162716 277366
rect 162768 273284 162820 273290
rect 162768 273226 162820 273232
rect 162676 194540 162728 194546
rect 162676 194482 162728 194488
rect 162780 93265 162808 273226
rect 163516 100774 163544 331230
rect 163608 274650 163636 390526
rect 163964 369164 164016 369170
rect 163964 369106 164016 369112
rect 163976 365634 164004 369106
rect 163964 365628 164016 365634
rect 163964 365570 164016 365576
rect 164068 327049 164096 394946
rect 164054 327040 164110 327049
rect 164054 326975 164110 326984
rect 163780 309868 163832 309874
rect 163780 309810 163832 309816
rect 163686 303512 163742 303521
rect 163686 303447 163742 303456
rect 163596 274644 163648 274650
rect 163596 274586 163648 274592
rect 163608 273290 163636 274586
rect 163596 273284 163648 273290
rect 163596 273226 163648 273232
rect 163700 267734 163728 303447
rect 163792 282878 163820 309810
rect 164160 305697 164188 618258
rect 166264 612876 166316 612882
rect 166264 612818 166316 612824
rect 164884 593428 164936 593434
rect 164884 593370 164936 593376
rect 164332 539640 164384 539646
rect 164332 539582 164384 539588
rect 164344 535362 164372 539582
rect 164332 535356 164384 535362
rect 164332 535298 164384 535304
rect 164896 389910 164924 593370
rect 164974 567896 165030 567905
rect 164974 567831 165030 567840
rect 164988 395010 165016 567831
rect 165068 509924 165120 509930
rect 165068 509866 165120 509872
rect 164976 395004 165028 395010
rect 164976 394946 165028 394952
rect 164884 389904 164936 389910
rect 164884 389846 164936 389852
rect 164884 388612 164936 388618
rect 164884 388554 164936 388560
rect 164896 379506 164924 388554
rect 164884 379500 164936 379506
rect 164884 379442 164936 379448
rect 164330 371920 164386 371929
rect 164330 371855 164386 371864
rect 164146 305688 164202 305697
rect 164146 305623 164202 305632
rect 163780 282872 163832 282878
rect 163780 282814 163832 282820
rect 163608 267706 163728 267734
rect 163608 265674 163636 267706
rect 163596 265668 163648 265674
rect 163596 265610 163648 265616
rect 163504 100768 163556 100774
rect 163504 100710 163556 100716
rect 162766 93256 162822 93265
rect 162766 93191 162822 93200
rect 163608 71097 163636 265610
rect 164240 262132 164292 262138
rect 164240 262074 164292 262080
rect 163780 259480 163832 259486
rect 163780 259422 163832 259428
rect 163688 253292 163740 253298
rect 163688 253234 163740 253240
rect 163700 222902 163728 253234
rect 163792 230450 163820 259422
rect 164146 251968 164202 251977
rect 164146 251903 164202 251912
rect 164160 251870 164188 251903
rect 164148 251864 164200 251870
rect 164148 251806 164200 251812
rect 163780 230444 163832 230450
rect 163780 230386 163832 230392
rect 163688 222896 163740 222902
rect 163688 222838 163740 222844
rect 164148 222896 164200 222902
rect 164148 222838 164200 222844
rect 164160 220833 164188 222838
rect 164146 220824 164202 220833
rect 164146 220759 164202 220768
rect 164160 133113 164188 220759
rect 164146 133104 164202 133113
rect 164146 133039 164202 133048
rect 164148 100768 164200 100774
rect 164148 100710 164200 100716
rect 164160 94489 164188 100710
rect 164146 94480 164202 94489
rect 164146 94415 164202 94424
rect 163594 71088 163650 71097
rect 163594 71023 163650 71032
rect 162124 28280 162176 28286
rect 162124 28222 162176 28228
rect 164252 24138 164280 262074
rect 164344 261497 164372 371855
rect 164896 369782 164924 379442
rect 164884 369776 164936 369782
rect 164884 369718 164936 369724
rect 164330 261488 164386 261497
rect 164330 261423 164386 261432
rect 164896 238678 164924 369718
rect 165080 369170 165108 509866
rect 165526 469296 165582 469305
rect 165526 469231 165582 469240
rect 165068 369164 165120 369170
rect 165068 369106 165120 369112
rect 165540 320793 165568 469231
rect 166276 448594 166304 612818
rect 166368 596174 166396 702442
rect 167644 615596 167696 615602
rect 167644 615538 167696 615544
rect 166368 596146 166488 596174
rect 166356 595468 166408 595474
rect 166356 595410 166408 595416
rect 166368 594862 166396 595410
rect 166356 594856 166408 594862
rect 166356 594798 166408 594804
rect 166460 574802 166488 596146
rect 166632 594856 166684 594862
rect 166632 594798 166684 594804
rect 166448 574796 166500 574802
rect 166448 574738 166500 574744
rect 166356 556844 166408 556850
rect 166356 556786 166408 556792
rect 166368 556238 166396 556786
rect 166356 556232 166408 556238
rect 166356 556174 166408 556180
rect 166368 451217 166396 556174
rect 166460 543046 166488 574738
rect 166448 543040 166500 543046
rect 166448 542982 166500 542988
rect 166354 451208 166410 451217
rect 166354 451143 166410 451152
rect 166368 450537 166396 451143
rect 166354 450528 166410 450537
rect 166354 450463 166410 450472
rect 166448 449948 166500 449954
rect 166448 449890 166500 449896
rect 166264 448588 166316 448594
rect 166264 448530 166316 448536
rect 166276 441614 166304 448530
rect 166460 448526 166488 449890
rect 166448 448520 166500 448526
rect 166448 448462 166500 448468
rect 166276 441586 166396 441614
rect 166368 430574 166396 441586
rect 166356 430568 166408 430574
rect 166356 430510 166408 430516
rect 166356 417444 166408 417450
rect 166356 417386 166408 417392
rect 166368 416838 166396 417386
rect 166356 416832 166408 416838
rect 166356 416774 166408 416780
rect 166356 329860 166408 329866
rect 166356 329802 166408 329808
rect 166368 324970 166396 329802
rect 166356 324964 166408 324970
rect 166356 324906 166408 324912
rect 165526 320784 165582 320793
rect 165526 320719 165582 320728
rect 164976 311160 165028 311166
rect 164976 311102 165028 311108
rect 164988 302258 165016 311102
rect 166460 309806 166488 448462
rect 166644 387870 166672 594798
rect 166816 471300 166868 471306
rect 166816 471242 166868 471248
rect 166724 416832 166776 416838
rect 166724 416774 166776 416780
rect 166632 387864 166684 387870
rect 166632 387806 166684 387812
rect 166736 329866 166764 416774
rect 166724 329860 166776 329866
rect 166724 329802 166776 329808
rect 166448 309800 166500 309806
rect 166448 309742 166500 309748
rect 164976 302252 165028 302258
rect 164976 302194 165028 302200
rect 164884 238672 164936 238678
rect 164884 238614 164936 238620
rect 164896 237318 164924 238614
rect 164884 237312 164936 237318
rect 164884 237254 164936 237260
rect 164988 195294 165016 302194
rect 166262 301744 166318 301753
rect 166262 301679 166318 301688
rect 166276 300898 166304 301679
rect 166264 300892 166316 300898
rect 166264 300834 166316 300840
rect 166460 296714 166488 309742
rect 166276 296686 166488 296714
rect 165528 295384 165580 295390
rect 165528 295326 165580 295332
rect 165540 282826 165568 295326
rect 165540 282798 165660 282826
rect 165528 262064 165580 262070
rect 165528 262006 165580 262012
rect 165540 261497 165568 262006
rect 165526 261488 165582 261497
rect 165526 261423 165582 261432
rect 165528 249620 165580 249626
rect 165528 249562 165580 249568
rect 165540 223582 165568 249562
rect 165632 245614 165660 282798
rect 166276 269074 166304 296686
rect 166828 287745 166856 471242
rect 167656 449954 167684 615538
rect 173808 614168 173860 614174
rect 173808 614110 173860 614116
rect 172428 604580 172480 604586
rect 172428 604522 172480 604528
rect 169024 603220 169076 603226
rect 169024 603162 169076 603168
rect 168288 574796 168340 574802
rect 168288 574738 168340 574744
rect 168196 545148 168248 545154
rect 168196 545090 168248 545096
rect 168104 478236 168156 478242
rect 168104 478178 168156 478184
rect 167644 449948 167696 449954
rect 167644 449890 167696 449896
rect 167000 447092 167052 447098
rect 167000 447034 167052 447040
rect 167012 446418 167040 447034
rect 167000 446412 167052 446418
rect 167000 446354 167052 446360
rect 167000 407788 167052 407794
rect 167000 407730 167052 407736
rect 167012 407182 167040 407730
rect 167000 407176 167052 407182
rect 167000 407118 167052 407124
rect 167012 402974 167040 407118
rect 167012 402946 167132 402974
rect 167000 365696 167052 365702
rect 167000 365638 167052 365644
rect 166906 344312 166962 344321
rect 166906 344247 166962 344256
rect 166814 287736 166870 287745
rect 166814 287671 166870 287680
rect 166814 280120 166870 280129
rect 166814 280055 166870 280064
rect 166828 279449 166856 280055
rect 166814 279440 166870 279449
rect 166814 279375 166870 279384
rect 166264 269068 166316 269074
rect 166264 269010 166316 269016
rect 166264 261520 166316 261526
rect 166264 261462 166316 261468
rect 165620 245608 165672 245614
rect 165620 245550 165672 245556
rect 165632 244934 165660 245550
rect 165620 244928 165672 244934
rect 165620 244870 165672 244876
rect 166276 230489 166304 261462
rect 166828 249121 166856 279375
rect 166814 249112 166870 249121
rect 166814 249047 166870 249056
rect 166356 245676 166408 245682
rect 166356 245618 166408 245624
rect 166368 237386 166396 245618
rect 166920 240038 166948 344247
rect 166908 240032 166960 240038
rect 166908 239974 166960 239980
rect 166356 237380 166408 237386
rect 166356 237322 166408 237328
rect 166262 230480 166318 230489
rect 166262 230415 166318 230424
rect 166368 224942 166396 237322
rect 166814 230480 166870 230489
rect 166814 230415 166870 230424
rect 166356 224936 166408 224942
rect 166356 224878 166408 224884
rect 165528 223576 165580 223582
rect 165528 223518 165580 223524
rect 164976 195288 165028 195294
rect 164976 195230 165028 195236
rect 165540 109002 165568 223518
rect 166828 162081 166856 230415
rect 166908 224936 166960 224942
rect 166908 224878 166960 224884
rect 166814 162072 166870 162081
rect 166814 162007 166870 162016
rect 166264 111920 166316 111926
rect 166264 111862 166316 111868
rect 165528 108996 165580 109002
rect 165528 108938 165580 108944
rect 165540 108322 165568 108938
rect 165528 108316 165580 108322
rect 165528 108258 165580 108264
rect 166276 71738 166304 111862
rect 166920 101522 166948 224878
rect 167012 218006 167040 365638
rect 167104 280129 167132 402946
rect 167644 387864 167696 387870
rect 167644 387806 167696 387812
rect 167656 386073 167684 387806
rect 167642 386064 167698 386073
rect 167642 385999 167698 386008
rect 167656 365702 167684 385999
rect 167644 365696 167696 365702
rect 167644 365638 167696 365644
rect 168116 331809 168144 478178
rect 168208 447098 168236 545090
rect 168196 447092 168248 447098
rect 168196 447034 168248 447040
rect 168194 423736 168250 423745
rect 168194 423671 168250 423680
rect 168102 331800 168158 331809
rect 168102 331735 168158 331744
rect 167644 285728 167696 285734
rect 167644 285670 167696 285676
rect 167090 280120 167146 280129
rect 167090 280055 167146 280064
rect 167000 218000 167052 218006
rect 167000 217942 167052 217948
rect 167656 151094 167684 285670
rect 167736 269068 167788 269074
rect 167736 269010 167788 269016
rect 167748 234598 167776 269010
rect 168208 260817 168236 423671
rect 168300 395350 168328 574738
rect 169036 562358 169064 603162
rect 171046 602032 171102 602041
rect 171046 601967 171102 601976
rect 170404 588600 170456 588606
rect 170404 588542 170456 588548
rect 169668 585880 169720 585886
rect 169668 585822 169720 585828
rect 169576 565208 169628 565214
rect 169576 565150 169628 565156
rect 169024 562352 169076 562358
rect 169024 562294 169076 562300
rect 169484 560312 169536 560318
rect 169484 560254 169536 560260
rect 168840 511964 168892 511970
rect 168840 511906 168892 511912
rect 168852 511290 168880 511906
rect 168840 511284 168892 511290
rect 168840 511226 168892 511232
rect 169496 471306 169524 560254
rect 169588 511290 169616 565150
rect 169576 511284 169628 511290
rect 169576 511226 169628 511232
rect 169574 475552 169630 475561
rect 169574 475487 169630 475496
rect 169484 471300 169536 471306
rect 169484 471242 169536 471248
rect 169484 458856 169536 458862
rect 169484 458798 169536 458804
rect 168288 395344 168340 395350
rect 168288 395286 168340 395292
rect 169496 389162 169524 458798
rect 169024 389156 169076 389162
rect 169024 389098 169076 389104
rect 169484 389156 169536 389162
rect 169484 389098 169536 389104
rect 169036 381546 169064 389098
rect 169024 381540 169076 381546
rect 169024 381482 169076 381488
rect 168380 360868 168432 360874
rect 168380 360810 168432 360816
rect 168392 360126 168420 360810
rect 168380 360120 168432 360126
rect 168380 360062 168432 360068
rect 169484 360120 169536 360126
rect 169484 360062 169536 360068
rect 168380 356720 168432 356726
rect 168380 356662 168432 356668
rect 168392 295390 168420 356662
rect 169022 333296 169078 333305
rect 169022 333231 169078 333240
rect 169036 332722 169064 333231
rect 169024 332716 169076 332722
rect 169024 332658 169076 332664
rect 169496 306610 169524 360062
rect 169484 306604 169536 306610
rect 169484 306546 169536 306552
rect 168472 298104 168524 298110
rect 168472 298046 168524 298052
rect 168484 297401 168512 298046
rect 168470 297392 168526 297401
rect 168470 297327 168526 297336
rect 168380 295384 168432 295390
rect 168380 295326 168432 295332
rect 168380 292664 168432 292670
rect 168380 292606 168432 292612
rect 169116 292664 169168 292670
rect 169116 292606 169168 292612
rect 168392 292534 168420 292606
rect 168380 292528 168432 292534
rect 168380 292470 168432 292476
rect 169024 282192 169076 282198
rect 168378 282160 168434 282169
rect 169024 282134 169076 282140
rect 168378 282095 168434 282104
rect 168194 260808 168250 260817
rect 168194 260743 168250 260752
rect 167828 254040 167880 254046
rect 167828 253982 167880 253988
rect 167840 250510 167868 253982
rect 167828 250504 167880 250510
rect 167828 250446 167880 250452
rect 168392 249626 168420 282095
rect 168470 250472 168526 250481
rect 168470 250407 168526 250416
rect 168380 249620 168432 249626
rect 168380 249562 168432 249568
rect 167736 234592 167788 234598
rect 167736 234534 167788 234540
rect 167644 151088 167696 151094
rect 167644 151030 167696 151036
rect 167656 117978 167684 151030
rect 167748 143614 167776 234534
rect 168484 230353 168512 250407
rect 168470 230344 168526 230353
rect 168470 230279 168526 230288
rect 167736 143608 167788 143614
rect 167736 143550 167788 143556
rect 167748 125594 167776 143550
rect 169036 135998 169064 282134
rect 169128 165714 169156 292606
rect 169588 270502 169616 475487
rect 169680 341465 169708 585822
rect 169760 528556 169812 528562
rect 169760 528498 169812 528504
rect 169772 416158 169800 528498
rect 169760 416152 169812 416158
rect 169760 416094 169812 416100
rect 169760 404320 169812 404326
rect 169760 404262 169812 404268
rect 169772 403034 169800 404262
rect 169760 403028 169812 403034
rect 169760 402970 169812 402976
rect 169772 368422 169800 402970
rect 170416 382129 170444 588542
rect 170494 541104 170550 541113
rect 170494 541039 170550 541048
rect 170508 528562 170536 541039
rect 170496 528556 170548 528562
rect 170496 528498 170548 528504
rect 170496 431248 170548 431254
rect 170496 431190 170548 431196
rect 170402 382120 170458 382129
rect 170402 382055 170458 382064
rect 170416 371142 170444 382055
rect 170404 371136 170456 371142
rect 170404 371078 170456 371084
rect 169760 368416 169812 368422
rect 169760 368358 169812 368364
rect 169772 364334 169800 368358
rect 169772 364306 169892 364334
rect 169666 341456 169722 341465
rect 169666 341391 169722 341400
rect 169668 316804 169720 316810
rect 169668 316746 169720 316752
rect 169680 316062 169708 316746
rect 169668 316056 169720 316062
rect 169668 315998 169720 316004
rect 169680 284170 169708 315998
rect 169668 284164 169720 284170
rect 169668 284106 169720 284112
rect 169576 270496 169628 270502
rect 169576 270438 169628 270444
rect 169206 269104 169262 269113
rect 169206 269039 169262 269048
rect 169220 251161 169248 269039
rect 169758 264888 169814 264897
rect 169758 264823 169814 264832
rect 169576 251184 169628 251190
rect 169206 251152 169262 251161
rect 169206 251087 169262 251096
rect 169574 251152 169576 251161
rect 169628 251152 169630 251161
rect 169574 251087 169630 251096
rect 169666 230344 169722 230353
rect 169666 230279 169722 230288
rect 169680 224913 169708 230279
rect 169666 224904 169722 224913
rect 169666 224839 169722 224848
rect 169116 165708 169168 165714
rect 169116 165650 169168 165656
rect 169128 145625 169156 165650
rect 169298 150648 169354 150657
rect 169298 150583 169354 150592
rect 169114 145616 169170 145625
rect 169114 145551 169170 145560
rect 169206 137320 169262 137329
rect 169206 137255 169262 137264
rect 169024 135992 169076 135998
rect 169024 135934 169076 135940
rect 169220 131102 169248 137255
rect 169208 131096 169260 131102
rect 169208 131038 169260 131044
rect 167736 125588 167788 125594
rect 167736 125530 167788 125536
rect 169220 122834 169248 131038
rect 169312 124817 169340 150583
rect 169298 124808 169354 124817
rect 169298 124743 169354 124752
rect 169220 122806 169616 122834
rect 167644 117972 167696 117978
rect 167644 117914 167696 117920
rect 169024 113212 169076 113218
rect 169024 113154 169076 113160
rect 166908 101516 166960 101522
rect 166908 101458 166960 101464
rect 169036 77246 169064 113154
rect 169116 111920 169168 111926
rect 169116 111862 169168 111868
rect 169128 97306 169156 111862
rect 169116 97300 169168 97306
rect 169116 97242 169168 97248
rect 169024 77240 169076 77246
rect 169024 77182 169076 77188
rect 166264 71732 166316 71738
rect 166264 71674 166316 71680
rect 169588 50386 169616 122806
rect 169680 112470 169708 224839
rect 169668 112464 169720 112470
rect 169668 112406 169720 112412
rect 169680 111926 169708 112406
rect 169668 111920 169720 111926
rect 169668 111862 169720 111868
rect 169772 68338 169800 264823
rect 169864 245682 169892 364306
rect 170508 287026 170536 431190
rect 171060 383489 171088 601967
rect 171784 583772 171836 583778
rect 171784 583714 171836 583720
rect 171796 388618 171824 583714
rect 172336 525088 172388 525094
rect 172336 525030 172388 525036
rect 171876 491972 171928 491978
rect 171876 491914 171928 491920
rect 171888 392018 171916 491914
rect 172348 402974 172376 525030
rect 172440 403646 172468 604522
rect 173164 581052 173216 581058
rect 173164 580994 173216 581000
rect 173176 554033 173204 580994
rect 173716 554872 173768 554878
rect 173716 554814 173768 554820
rect 173256 554056 173308 554062
rect 173162 554024 173218 554033
rect 173256 553998 173308 554004
rect 173162 553959 173218 553968
rect 173164 532024 173216 532030
rect 173164 531966 173216 531972
rect 173176 469305 173204 531966
rect 173268 523705 173296 553998
rect 173254 523696 173310 523705
rect 173254 523631 173310 523640
rect 173622 489152 173678 489161
rect 173622 489087 173678 489096
rect 173162 469296 173218 469305
rect 173162 469231 173218 469240
rect 172518 453928 172574 453937
rect 172518 453863 172574 453872
rect 172532 438161 172560 453863
rect 173164 444372 173216 444378
rect 173164 444314 173216 444320
rect 173176 443086 173204 444314
rect 173164 443080 173216 443086
rect 173164 443022 173216 443028
rect 172518 438152 172574 438161
rect 172518 438087 172574 438096
rect 172428 403640 172480 403646
rect 172428 403582 172480 403588
rect 172072 402946 172376 402974
rect 172072 400926 172100 402946
rect 172060 400920 172112 400926
rect 172060 400862 172112 400868
rect 171876 392012 171928 392018
rect 171876 391954 171928 391960
rect 171968 390652 172020 390658
rect 171968 390594 172020 390600
rect 171784 388612 171836 388618
rect 171784 388554 171836 388560
rect 171046 383480 171102 383489
rect 171046 383415 171102 383424
rect 171876 375352 171928 375358
rect 171876 375294 171928 375300
rect 171140 364336 171192 364342
rect 171140 364278 171192 364284
rect 171046 347032 171102 347041
rect 171046 346967 171102 346976
rect 170496 287020 170548 287026
rect 170496 286962 170548 286968
rect 170508 285734 170536 286962
rect 170496 285728 170548 285734
rect 170496 285670 170548 285676
rect 169944 284164 169996 284170
rect 169944 284106 169996 284112
rect 169852 245676 169904 245682
rect 169852 245618 169904 245624
rect 169956 227798 169984 284106
rect 170312 264988 170364 264994
rect 170312 264930 170364 264936
rect 170324 264897 170352 264930
rect 170310 264888 170366 264897
rect 170310 264823 170366 264832
rect 170770 254280 170826 254289
rect 170770 254215 170826 254224
rect 170784 254046 170812 254215
rect 170772 254040 170824 254046
rect 170772 253982 170824 253988
rect 171060 246265 171088 346967
rect 171046 246256 171102 246265
rect 171046 246191 171102 246200
rect 171152 238762 171180 364278
rect 171782 258904 171838 258913
rect 171782 258839 171838 258848
rect 171060 238734 171180 238762
rect 171060 233238 171088 238734
rect 171048 233232 171100 233238
rect 171048 233174 171100 233180
rect 171060 231810 171088 233174
rect 171048 231804 171100 231810
rect 171048 231746 171100 231752
rect 169944 227792 169996 227798
rect 169944 227734 169996 227740
rect 170496 227792 170548 227798
rect 170496 227734 170548 227740
rect 170404 194540 170456 194546
rect 170404 194482 170456 194488
rect 170416 136610 170444 194482
rect 170508 193866 170536 227734
rect 170496 193860 170548 193866
rect 170496 193802 170548 193808
rect 170404 136604 170456 136610
rect 170404 136546 170456 136552
rect 171060 84182 171088 231746
rect 169852 84176 169904 84182
rect 169852 84118 169904 84124
rect 171048 84176 171100 84182
rect 171048 84118 171100 84124
rect 169864 81326 169892 84118
rect 169852 81320 169904 81326
rect 169852 81262 169904 81268
rect 171796 75206 171824 258839
rect 171888 233209 171916 375294
rect 171980 364342 172008 390594
rect 172072 375358 172100 400862
rect 172428 392012 172480 392018
rect 172428 391954 172480 391960
rect 172440 389094 172468 391954
rect 172428 389088 172480 389094
rect 172428 389030 172480 389036
rect 172060 375352 172112 375358
rect 172060 375294 172112 375300
rect 171968 364336 172020 364342
rect 171968 364278 172020 364284
rect 173176 311166 173204 443022
rect 173256 398200 173308 398206
rect 173256 398142 173308 398148
rect 173268 379409 173296 398142
rect 173636 391270 173664 489087
rect 173728 457502 173756 554814
rect 173716 457496 173768 457502
rect 173716 457438 173768 457444
rect 173820 425746 173848 614110
rect 175186 608696 175242 608705
rect 175186 608631 175242 608640
rect 174544 558952 174596 558958
rect 174544 558894 174596 558900
rect 174556 486470 174584 558894
rect 175004 487824 175056 487830
rect 175004 487766 175056 487772
rect 174544 486464 174596 486470
rect 174544 486406 174596 486412
rect 174544 461032 174596 461038
rect 174544 460974 174596 460980
rect 174556 440298 174584 460974
rect 174544 440292 174596 440298
rect 174544 440234 174596 440240
rect 173808 425740 173860 425746
rect 173808 425682 173860 425688
rect 173820 412634 173848 425682
rect 173728 412606 173848 412634
rect 173624 391264 173676 391270
rect 173624 391206 173676 391212
rect 173636 390658 173664 391206
rect 173624 390652 173676 390658
rect 173624 390594 173676 390600
rect 173530 388920 173586 388929
rect 173530 388855 173586 388864
rect 173544 387705 173572 388855
rect 173530 387696 173586 387705
rect 173530 387631 173586 387640
rect 173254 379400 173310 379409
rect 173254 379335 173310 379344
rect 173254 346488 173310 346497
rect 173254 346423 173310 346432
rect 173164 311160 173216 311166
rect 173164 311102 173216 311108
rect 172520 306604 172572 306610
rect 172520 306546 172572 306552
rect 172058 242176 172114 242185
rect 172058 242111 172114 242120
rect 171874 233200 171930 233209
rect 171874 233135 171930 233144
rect 171888 220114 171916 233135
rect 171876 220108 171928 220114
rect 171876 220050 171928 220056
rect 171888 219434 171916 220050
rect 171888 219406 172008 219434
rect 171876 216708 171928 216714
rect 171876 216650 171928 216656
rect 171888 102241 171916 216650
rect 171980 116521 172008 219406
rect 172072 217938 172100 242111
rect 172532 239465 172560 306546
rect 173268 260166 173296 346423
rect 173728 307766 173756 412606
rect 173806 387696 173862 387705
rect 173806 387631 173862 387640
rect 173716 307760 173768 307766
rect 173716 307702 173768 307708
rect 173348 264240 173400 264246
rect 173348 264182 173400 264188
rect 173256 260160 173308 260166
rect 173256 260102 173308 260108
rect 173268 258074 173296 260102
rect 173176 258046 173296 258074
rect 172518 239456 172574 239465
rect 172518 239391 172574 239400
rect 172060 217932 172112 217938
rect 172060 217874 172112 217880
rect 172072 216714 172100 217874
rect 172060 216708 172112 216714
rect 172060 216650 172112 216656
rect 171966 116512 172022 116521
rect 171966 116447 172022 116456
rect 171874 102232 171930 102241
rect 171874 102167 171930 102176
rect 172426 102232 172482 102241
rect 172426 102167 172482 102176
rect 172440 95849 172468 102167
rect 172426 95840 172482 95849
rect 172426 95775 172482 95784
rect 171784 75200 171836 75206
rect 171784 75142 171836 75148
rect 173176 73817 173204 258046
rect 173360 233073 173388 264182
rect 173820 253230 173848 387631
rect 174268 383036 174320 383042
rect 174268 382978 174320 382984
rect 174280 375358 174308 382978
rect 174268 375352 174320 375358
rect 174268 375294 174320 375300
rect 174556 321609 174584 440234
rect 175016 398206 175044 487766
rect 175096 479596 175148 479602
rect 175096 479538 175148 479544
rect 175004 398200 175056 398206
rect 175004 398142 175056 398148
rect 174634 366344 174690 366353
rect 174634 366279 174690 366288
rect 174542 321600 174598 321609
rect 174542 321535 174598 321544
rect 174544 256692 174596 256698
rect 174544 256634 174596 256640
rect 173808 253224 173860 253230
rect 173808 253166 173860 253172
rect 173808 243228 173860 243234
rect 173808 243170 173860 243176
rect 173346 233064 173402 233073
rect 173346 232999 173402 233008
rect 173360 229094 173388 232999
rect 173360 229066 173756 229094
rect 173728 151814 173756 229066
rect 173820 209778 173848 243170
rect 173808 209772 173860 209778
rect 173808 209714 173860 209720
rect 173820 209098 173848 209714
rect 173808 209092 173860 209098
rect 173808 209034 173860 209040
rect 173268 151786 173756 151814
rect 173268 148073 173296 151786
rect 173254 148064 173310 148073
rect 173254 147999 173310 148008
rect 173268 141545 173296 147999
rect 173254 141536 173310 141545
rect 173254 141471 173310 141480
rect 173256 140072 173308 140078
rect 173256 140014 173308 140020
rect 173268 110362 173296 140014
rect 173256 110356 173308 110362
rect 173256 110298 173308 110304
rect 173820 95305 173848 209034
rect 173806 95296 173862 95305
rect 173806 95231 173862 95240
rect 173162 73808 173218 73817
rect 173162 73743 173218 73752
rect 169760 68332 169812 68338
rect 169760 68274 169812 68280
rect 169576 50380 169628 50386
rect 169576 50322 169628 50328
rect 174556 33794 174584 256634
rect 174648 253298 174676 366279
rect 175108 322289 175136 479538
rect 175200 424386 175228 608631
rect 177304 607232 177356 607238
rect 177304 607174 177356 607180
rect 176568 605940 176620 605946
rect 176568 605882 176620 605888
rect 176016 586560 176068 586566
rect 176016 586502 176068 586508
rect 175924 466472 175976 466478
rect 175924 466414 175976 466420
rect 175188 424380 175240 424386
rect 175188 424322 175240 424328
rect 175094 322280 175150 322289
rect 175094 322215 175150 322224
rect 175186 321600 175242 321609
rect 175186 321535 175242 321544
rect 175200 296002 175228 321535
rect 175936 315353 175964 466414
rect 176028 458862 176056 586502
rect 176108 490612 176160 490618
rect 176108 490554 176160 490560
rect 176016 458856 176068 458862
rect 176016 458798 176068 458804
rect 176120 453801 176148 490554
rect 176106 453792 176162 453801
rect 176106 453727 176162 453736
rect 176476 451376 176528 451382
rect 176476 451318 176528 451324
rect 176014 444272 176070 444281
rect 176014 444207 176070 444216
rect 176028 323678 176056 444207
rect 176108 395344 176160 395350
rect 176108 395286 176160 395292
rect 176120 366994 176148 395286
rect 176108 366988 176160 366994
rect 176108 366930 176160 366936
rect 176016 323672 176068 323678
rect 176014 323640 176016 323649
rect 176068 323640 176070 323649
rect 176014 323575 176070 323584
rect 176028 323549 176056 323575
rect 175922 315344 175978 315353
rect 175922 315279 175978 315288
rect 175280 307760 175332 307766
rect 175280 307702 175332 307708
rect 175188 295996 175240 296002
rect 175188 295938 175240 295944
rect 175188 294636 175240 294642
rect 175188 294578 175240 294584
rect 175200 294030 175228 294578
rect 175188 294024 175240 294030
rect 175188 293966 175240 293972
rect 175200 277394 175228 293966
rect 175292 289785 175320 307702
rect 175278 289776 175334 289785
rect 175278 289711 175334 289720
rect 175292 289105 175320 289711
rect 175278 289096 175334 289105
rect 175278 289031 175334 289040
rect 175936 282946 175964 315279
rect 176488 307154 176516 451318
rect 176580 418810 176608 605882
rect 177316 452577 177344 607174
rect 178774 599584 178830 599593
rect 178774 599519 178830 599528
rect 177948 587172 178000 587178
rect 177948 587114 178000 587120
rect 177856 561740 177908 561746
rect 177856 561682 177908 561688
rect 177396 540252 177448 540258
rect 177396 540194 177448 540200
rect 177408 468489 177436 540194
rect 177394 468480 177450 468489
rect 177394 468415 177450 468424
rect 177578 468480 177634 468489
rect 177578 468415 177634 468424
rect 176658 452568 176714 452577
rect 176658 452503 176714 452512
rect 177302 452568 177358 452577
rect 177302 452503 177358 452512
rect 176672 451897 176700 452503
rect 176658 451888 176714 451897
rect 176658 451823 176714 451832
rect 176672 427786 176700 451823
rect 176660 427780 176712 427786
rect 176660 427722 176712 427728
rect 176672 427106 176700 427722
rect 177302 427136 177358 427145
rect 176660 427100 176712 427106
rect 177302 427071 177358 427080
rect 176660 427042 176712 427048
rect 176568 418804 176620 418810
rect 176568 418746 176620 418752
rect 176658 367024 176714 367033
rect 176658 366959 176714 366968
rect 176752 366988 176804 366994
rect 176016 307148 176068 307154
rect 176016 307090 176068 307096
rect 176476 307148 176528 307154
rect 176476 307090 176528 307096
rect 176028 306406 176056 307090
rect 176016 306400 176068 306406
rect 176016 306342 176068 306348
rect 176028 283626 176056 306342
rect 176106 289776 176162 289785
rect 176106 289711 176162 289720
rect 176016 283620 176068 283626
rect 176016 283562 176068 283568
rect 175924 282940 175976 282946
rect 175924 282882 175976 282888
rect 175924 280696 175976 280702
rect 175924 280638 175976 280644
rect 175108 277366 175228 277394
rect 174636 253292 174688 253298
rect 174636 253234 174688 253240
rect 174728 253224 174780 253230
rect 174728 253166 174780 253172
rect 174740 234161 174768 253166
rect 174726 234152 174782 234161
rect 174726 234087 174782 234096
rect 175108 202230 175136 277366
rect 175186 234560 175242 234569
rect 175186 234495 175242 234504
rect 175200 234161 175228 234495
rect 175186 234152 175242 234161
rect 175186 234087 175242 234096
rect 175096 202224 175148 202230
rect 175096 202166 175148 202172
rect 175200 92449 175228 234087
rect 175936 180878 175964 280638
rect 176120 267073 176148 289711
rect 176568 284980 176620 284986
rect 176568 284922 176620 284928
rect 176106 267064 176162 267073
rect 176106 266999 176162 267008
rect 175924 180872 175976 180878
rect 175924 180814 175976 180820
rect 175936 144294 175964 180814
rect 175924 144288 175976 144294
rect 175924 144230 175976 144236
rect 175924 135924 175976 135930
rect 175924 135866 175976 135872
rect 175936 124098 175964 135866
rect 175924 124092 175976 124098
rect 175924 124034 175976 124040
rect 175186 92440 175242 92449
rect 175186 92375 175242 92384
rect 176580 91050 176608 284922
rect 176672 243234 176700 366959
rect 176752 366930 176804 366936
rect 176764 366382 176792 366930
rect 176752 366376 176804 366382
rect 176752 366318 176804 366324
rect 176764 307222 176792 366318
rect 177316 341562 177344 427071
rect 177592 419665 177620 468415
rect 177578 419656 177634 419665
rect 177578 419591 177634 419600
rect 177868 410582 177896 561682
rect 177960 439550 177988 587114
rect 178684 569220 178736 569226
rect 178684 569162 178736 569168
rect 178408 541680 178460 541686
rect 178408 541622 178460 541628
rect 178420 541006 178448 541622
rect 178408 541000 178460 541006
rect 178408 540942 178460 540948
rect 178696 538150 178724 569162
rect 178788 567866 178816 599519
rect 179236 589348 179288 589354
rect 179236 589290 179288 589296
rect 179052 580440 179104 580446
rect 179052 580382 179104 580388
rect 178776 567860 178828 567866
rect 178776 567802 178828 567808
rect 178684 538144 178736 538150
rect 178684 538086 178736 538092
rect 178684 458312 178736 458318
rect 178684 458254 178736 458260
rect 177948 439544 178000 439550
rect 177948 439486 178000 439492
rect 178040 438184 178092 438190
rect 178040 438126 178092 438132
rect 177948 436824 178000 436830
rect 177948 436766 178000 436772
rect 177856 410576 177908 410582
rect 177856 410518 177908 410524
rect 177488 404388 177540 404394
rect 177488 404330 177540 404336
rect 177396 393372 177448 393378
rect 177396 393314 177448 393320
rect 177408 367033 177436 393314
rect 177500 383654 177528 404330
rect 177488 383648 177540 383654
rect 177488 383590 177540 383596
rect 177394 367024 177450 367033
rect 177394 366959 177450 366968
rect 177304 341556 177356 341562
rect 177304 341498 177356 341504
rect 177578 340912 177634 340921
rect 177578 340847 177634 340856
rect 177592 338881 177620 340847
rect 177578 338872 177634 338881
rect 177578 338807 177634 338816
rect 176752 307216 176804 307222
rect 176752 307158 176804 307164
rect 176752 307080 176804 307086
rect 176752 307022 176804 307028
rect 176764 306513 176792 307022
rect 176750 306504 176806 306513
rect 176750 306439 176806 306448
rect 177856 292596 177908 292602
rect 177856 292538 177908 292544
rect 177868 292126 177896 292538
rect 177856 292120 177908 292126
rect 177856 292062 177908 292068
rect 177396 267096 177448 267102
rect 177396 267038 177448 267044
rect 177302 257408 177358 257417
rect 177302 257343 177358 257352
rect 176660 243228 176712 243234
rect 176660 243170 176712 243176
rect 176568 91044 176620 91050
rect 176568 90986 176620 90992
rect 174544 33788 174596 33794
rect 174544 33730 174596 33736
rect 164240 24132 164292 24138
rect 164240 24074 164292 24080
rect 161480 22772 161532 22778
rect 161480 22714 161532 22720
rect 177316 17270 177344 257343
rect 177408 228993 177436 267038
rect 177394 228984 177450 228993
rect 177394 228919 177450 228928
rect 177408 227769 177436 228919
rect 177394 227760 177450 227769
rect 177394 227695 177450 227704
rect 177394 155408 177450 155417
rect 177394 155343 177450 155352
rect 177408 107642 177436 155343
rect 177486 145752 177542 145761
rect 177486 145687 177542 145696
rect 177500 117230 177528 145687
rect 177868 145042 177896 292062
rect 177960 275330 177988 436766
rect 178052 435305 178080 438126
rect 178038 435296 178094 435305
rect 178038 435231 178094 435240
rect 178040 431928 178092 431934
rect 178040 431870 178092 431876
rect 178052 387569 178080 431870
rect 178038 387560 178094 387569
rect 178038 387495 178094 387504
rect 178052 387025 178080 387495
rect 178038 387016 178094 387025
rect 178038 386951 178094 386960
rect 178038 341456 178094 341465
rect 178038 341391 178094 341400
rect 178052 337929 178080 341391
rect 178038 337920 178094 337929
rect 178038 337855 178094 337864
rect 178052 337482 178080 337855
rect 178040 337476 178092 337482
rect 178040 337418 178092 337424
rect 178038 337376 178094 337385
rect 178038 337311 178094 337320
rect 178052 336870 178080 337311
rect 178130 337240 178186 337249
rect 178130 337175 178186 337184
rect 178040 336864 178092 336870
rect 178040 336806 178092 336812
rect 178144 336802 178172 337175
rect 178132 336796 178184 336802
rect 178132 336738 178184 336744
rect 178590 334656 178646 334665
rect 178590 334591 178646 334600
rect 178604 334082 178632 334591
rect 178592 334076 178644 334082
rect 178592 334018 178644 334024
rect 178696 319433 178724 458254
rect 178868 389224 178920 389230
rect 178868 389166 178920 389172
rect 178774 387560 178830 387569
rect 178774 387495 178830 387504
rect 178788 322153 178816 387495
rect 178880 360126 178908 389166
rect 179064 372570 179092 580382
rect 179144 541680 179196 541686
rect 179144 541622 179196 541628
rect 179156 532710 179184 541622
rect 179144 532704 179196 532710
rect 179144 532646 179196 532652
rect 179248 438190 179276 589290
rect 179340 580310 179368 702918
rect 188344 702908 188396 702914
rect 188344 702850 188396 702856
rect 187608 702772 187660 702778
rect 187608 702714 187660 702720
rect 184296 612808 184348 612814
rect 184296 612750 184348 612756
rect 182824 607300 182876 607306
rect 182824 607242 182876 607248
rect 180706 604616 180762 604625
rect 180706 604551 180762 604560
rect 180064 601792 180116 601798
rect 180064 601734 180116 601740
rect 179328 580304 179380 580310
rect 179328 580246 179380 580252
rect 179420 572008 179472 572014
rect 179420 571950 179472 571956
rect 179432 570654 179460 571950
rect 179420 570648 179472 570654
rect 179420 570590 179472 570596
rect 180076 560998 180104 601734
rect 180524 570648 180576 570654
rect 180524 570590 180576 570596
rect 180064 560992 180116 560998
rect 180064 560934 180116 560940
rect 180064 554804 180116 554810
rect 180064 554746 180116 554752
rect 180076 545086 180104 554746
rect 180064 545080 180116 545086
rect 180064 545022 180116 545028
rect 180536 485790 180564 570590
rect 180616 552152 180668 552158
rect 180616 552094 180668 552100
rect 179420 485784 179472 485790
rect 179420 485726 179472 485732
rect 180524 485784 180576 485790
rect 180524 485726 180576 485732
rect 179432 485110 179460 485726
rect 179420 485104 179472 485110
rect 179420 485046 179472 485052
rect 180430 474192 180486 474201
rect 180430 474127 180486 474136
rect 180064 452736 180116 452742
rect 180064 452678 180116 452684
rect 180076 444378 180104 452678
rect 180064 444372 180116 444378
rect 180064 444314 180116 444320
rect 179236 438184 179288 438190
rect 179236 438126 179288 438132
rect 180444 403617 180472 474127
rect 180524 468580 180576 468586
rect 180524 468522 180576 468528
rect 180430 403608 180486 403617
rect 180430 403543 180486 403552
rect 180156 398200 180208 398206
rect 180156 398142 180208 398148
rect 180168 390969 180196 398142
rect 180536 396778 180564 468522
rect 180628 452742 180656 552094
rect 180616 452736 180668 452742
rect 180616 452678 180668 452684
rect 180614 400208 180670 400217
rect 180614 400143 180670 400152
rect 180524 396772 180576 396778
rect 180524 396714 180576 396720
rect 180628 393417 180656 400143
rect 180614 393408 180670 393417
rect 180614 393343 180670 393352
rect 180720 393314 180748 604551
rect 181812 603152 181864 603158
rect 181812 603094 181864 603100
rect 181444 584452 181496 584458
rect 181444 584394 181496 584400
rect 181456 401674 181484 584394
rect 181536 543040 181588 543046
rect 181536 542982 181588 542988
rect 181548 534041 181576 542982
rect 181534 534032 181590 534041
rect 181534 533967 181590 533976
rect 181548 466546 181576 533967
rect 181536 466540 181588 466546
rect 181536 466482 181588 466488
rect 181444 401668 181496 401674
rect 181444 401610 181496 401616
rect 180628 393286 180748 393314
rect 180154 390960 180210 390969
rect 180154 390895 180210 390904
rect 180062 387560 180118 387569
rect 180062 387495 180118 387504
rect 179052 372564 179104 372570
rect 179052 372506 179104 372512
rect 180076 372502 180104 387495
rect 180168 380769 180196 390895
rect 180628 387569 180656 393286
rect 180706 393136 180762 393145
rect 180706 393071 180762 393080
rect 180614 387560 180670 387569
rect 180614 387495 180670 387504
rect 180720 383761 180748 393071
rect 180706 383752 180762 383761
rect 180706 383687 180762 383696
rect 180706 383616 180762 383625
rect 180706 383551 180762 383560
rect 180154 380760 180210 380769
rect 180154 380695 180210 380704
rect 180720 374105 180748 383551
rect 181456 381750 181484 401610
rect 181536 399492 181588 399498
rect 181536 399434 181588 399440
rect 181548 384985 181576 399434
rect 181534 384976 181590 384985
rect 181534 384911 181590 384920
rect 181824 381993 181852 603094
rect 181996 515432 182048 515438
rect 181996 515374 182048 515380
rect 181902 454744 181958 454753
rect 181902 454679 181958 454688
rect 181916 400217 181944 454679
rect 181902 400208 181958 400217
rect 181902 400143 181958 400152
rect 182008 393961 182036 515374
rect 182088 466540 182140 466546
rect 182088 466482 182140 466488
rect 182100 465730 182128 466482
rect 182088 465724 182140 465730
rect 182088 465666 182140 465672
rect 181994 393952 182050 393961
rect 181994 393887 182050 393896
rect 182836 390833 182864 607242
rect 184204 599072 184256 599078
rect 184204 599014 184256 599020
rect 184216 558890 184244 599014
rect 184308 591326 184336 612750
rect 186962 600672 187018 600681
rect 186962 600607 187018 600616
rect 186226 595504 186282 595513
rect 186226 595439 186282 595448
rect 184296 591320 184348 591326
rect 184296 591262 184348 591268
rect 184848 581120 184900 581126
rect 184848 581062 184900 581068
rect 184204 558884 184256 558890
rect 184204 558826 184256 558832
rect 184204 552084 184256 552090
rect 184204 552026 184256 552032
rect 184216 538218 184244 552026
rect 184756 543788 184808 543794
rect 184756 543730 184808 543736
rect 184664 542360 184716 542366
rect 184664 542302 184716 542308
rect 184204 538212 184256 538218
rect 184676 538214 184704 542302
rect 184768 540258 184796 543730
rect 184756 540252 184808 540258
rect 184756 540194 184808 540200
rect 184676 538186 184796 538214
rect 184204 538154 184256 538160
rect 182914 536072 182970 536081
rect 182914 536007 182970 536016
rect 182928 525162 182956 536007
rect 183376 530664 183428 530670
rect 183376 530606 183428 530612
rect 182916 525156 182968 525162
rect 182916 525098 182968 525104
rect 183388 449954 183416 530606
rect 184664 512644 184716 512650
rect 184664 512586 184716 512592
rect 183466 485072 183522 485081
rect 183466 485007 183522 485016
rect 183376 449948 183428 449954
rect 183376 449890 183428 449896
rect 183374 446584 183430 446593
rect 183374 446519 183430 446528
rect 182916 403640 182968 403646
rect 182916 403582 182968 403588
rect 182822 390824 182878 390833
rect 182822 390759 182878 390768
rect 181994 389192 182050 389201
rect 181994 389127 182050 389136
rect 181810 381984 181866 381993
rect 181810 381919 181866 381928
rect 181444 381744 181496 381750
rect 181444 381686 181496 381692
rect 182008 375193 182036 389127
rect 182088 382220 182140 382226
rect 182088 382162 182140 382168
rect 182100 381750 182128 382162
rect 182088 381744 182140 381750
rect 182088 381686 182140 381692
rect 181994 375184 182050 375193
rect 181994 375119 182050 375128
rect 180706 374096 180762 374105
rect 180706 374031 180762 374040
rect 180706 373960 180762 373969
rect 180706 373895 180762 373904
rect 180064 372496 180116 372502
rect 180064 372438 180116 372444
rect 180076 371822 180104 372438
rect 179420 371816 179472 371822
rect 179420 371758 179472 371764
rect 180064 371816 180116 371822
rect 180064 371758 180116 371764
rect 178868 360120 178920 360126
rect 178868 360062 178920 360068
rect 179326 343088 179382 343097
rect 179326 343023 179382 343032
rect 178868 334008 178920 334014
rect 178868 333950 178920 333956
rect 178774 322144 178830 322153
rect 178774 322079 178830 322088
rect 178682 319424 178738 319433
rect 178682 319359 178738 319368
rect 178696 317490 178724 319359
rect 178684 317484 178736 317490
rect 178684 317426 178736 317432
rect 178696 316034 178724 317426
rect 178696 316006 178816 316034
rect 178592 308508 178644 308514
rect 178592 308450 178644 308456
rect 178604 306374 178632 308450
rect 178604 306346 178724 306374
rect 177948 275324 178000 275330
rect 177948 275266 178000 275272
rect 177946 227760 178002 227769
rect 177946 227695 178002 227704
rect 177960 151162 177988 227695
rect 177948 151156 178000 151162
rect 177948 151098 178000 151104
rect 177856 145036 177908 145042
rect 177856 144978 177908 144984
rect 177868 142154 177896 144978
rect 177592 142126 177896 142154
rect 177592 133890 177620 142126
rect 178696 138718 178724 306346
rect 178788 280702 178816 316006
rect 178880 292126 178908 333950
rect 179340 302297 179368 343023
rect 179326 302288 179382 302297
rect 179326 302223 179382 302232
rect 179326 302152 179382 302161
rect 179326 302087 179382 302096
rect 179340 301510 179368 302087
rect 179328 301504 179380 301510
rect 179328 301446 179380 301452
rect 178868 292120 178920 292126
rect 178868 292062 178920 292068
rect 178960 291916 179012 291922
rect 178960 291858 179012 291864
rect 178776 280696 178828 280702
rect 178776 280638 178828 280644
rect 178972 271289 179000 291858
rect 179326 287736 179382 287745
rect 179326 287671 179382 287680
rect 178958 271280 179014 271289
rect 178958 271215 179014 271224
rect 178776 269136 178828 269142
rect 178776 269078 178828 269084
rect 178788 144226 178816 269078
rect 178868 257372 178920 257378
rect 178868 257314 178920 257320
rect 178880 236745 178908 257314
rect 179340 253230 179368 287671
rect 179328 253224 179380 253230
rect 179328 253166 179380 253172
rect 179432 247625 179460 371758
rect 180064 369232 180116 369238
rect 180064 369174 180116 369180
rect 180076 364342 180104 369174
rect 180720 364449 180748 373895
rect 180706 364440 180762 364449
rect 180706 364375 180762 364384
rect 180064 364336 180116 364342
rect 180064 364278 180116 364284
rect 180616 364336 180668 364342
rect 180616 364278 180668 364284
rect 180706 364304 180762 364313
rect 180628 354770 180656 364278
rect 180706 364239 180762 364248
rect 180720 354929 180748 364239
rect 180706 354920 180762 354929
rect 180706 354855 180762 354864
rect 180628 354742 180748 354770
rect 180614 354648 180670 354657
rect 180614 354583 180670 354592
rect 180628 347041 180656 354583
rect 180614 347032 180670 347041
rect 180614 346967 180670 346976
rect 180614 341456 180670 341465
rect 180614 341391 180670 341400
rect 180062 300112 180118 300121
rect 180062 300047 180118 300056
rect 180076 296041 180104 300047
rect 180062 296032 180118 296041
rect 180062 295967 180118 295976
rect 180156 282940 180208 282946
rect 180156 282882 180208 282888
rect 180062 254008 180118 254017
rect 180062 253943 180118 253952
rect 179418 247616 179474 247625
rect 179418 247551 179474 247560
rect 178866 236736 178922 236745
rect 178866 236671 178922 236680
rect 178868 231124 178920 231130
rect 178868 231066 178920 231072
rect 178880 229090 178908 231066
rect 178868 229084 178920 229090
rect 178868 229026 178920 229032
rect 178880 227798 178908 229026
rect 178868 227792 178920 227798
rect 178868 227734 178920 227740
rect 179328 227792 179380 227798
rect 179328 227734 179380 227740
rect 178866 156224 178922 156233
rect 178866 156159 178922 156168
rect 178776 144220 178828 144226
rect 178776 144162 178828 144168
rect 178684 138712 178736 138718
rect 178684 138654 178736 138660
rect 177580 133884 177632 133890
rect 177580 133826 177632 133832
rect 177488 117224 177540 117230
rect 177488 117166 177540 117172
rect 177396 107636 177448 107642
rect 177396 107578 177448 107584
rect 178696 105602 178724 138654
rect 178880 117298 178908 156159
rect 179236 126268 179288 126274
rect 179236 126210 179288 126216
rect 178868 117292 178920 117298
rect 178868 117234 178920 117240
rect 177396 105596 177448 105602
rect 177396 105538 177448 105544
rect 178684 105596 178736 105602
rect 178684 105538 178736 105544
rect 177408 78606 177436 105538
rect 177488 95260 177540 95266
rect 177488 95202 177540 95208
rect 177500 79966 177528 95202
rect 178038 81424 178094 81433
rect 178038 81359 178094 81368
rect 177488 79960 177540 79966
rect 177488 79902 177540 79908
rect 178052 78674 178080 81359
rect 178040 78668 178092 78674
rect 178040 78610 178092 78616
rect 177396 78600 177448 78606
rect 177396 78542 177448 78548
rect 179248 39370 179276 126210
rect 179340 81433 179368 227734
rect 179326 81424 179382 81433
rect 179326 81359 179382 81368
rect 180076 80753 180104 253943
rect 180168 171834 180196 282882
rect 180628 254017 180656 341391
rect 180614 254008 180670 254017
rect 180614 253943 180670 253952
rect 180340 247716 180392 247722
rect 180340 247658 180392 247664
rect 180246 231296 180302 231305
rect 180246 231231 180302 231240
rect 180260 199345 180288 231231
rect 180352 224233 180380 247658
rect 180720 240786 180748 354742
rect 181904 319116 181956 319122
rect 181904 319058 181956 319064
rect 181444 304292 181496 304298
rect 181444 304234 181496 304240
rect 180708 240780 180760 240786
rect 180708 240722 180760 240728
rect 180720 240258 180748 240722
rect 180720 240230 180932 240258
rect 180904 234161 180932 240230
rect 180890 234152 180946 234161
rect 180890 234087 180946 234096
rect 180338 224224 180394 224233
rect 180338 224159 180394 224168
rect 180246 199336 180302 199345
rect 180246 199271 180302 199280
rect 180156 171828 180208 171834
rect 180156 171770 180208 171776
rect 180156 131844 180208 131850
rect 180156 131786 180208 131792
rect 180168 124166 180196 131786
rect 180156 124160 180208 124166
rect 180156 124102 180208 124108
rect 180062 80744 180118 80753
rect 180062 80679 180118 80688
rect 179236 39364 179288 39370
rect 179236 39306 179288 39312
rect 180168 18630 180196 124102
rect 180260 97986 180288 199271
rect 180800 101516 180852 101522
rect 180800 101458 180852 101464
rect 180248 97980 180300 97986
rect 180248 97922 180300 97928
rect 180812 70378 180840 101458
rect 181456 82113 181484 304234
rect 181916 268394 181944 319058
rect 181904 268388 181956 268394
rect 181904 268330 181956 268336
rect 182008 247761 182036 375119
rect 181994 247752 182050 247761
rect 181994 247687 182050 247696
rect 181536 247104 181588 247110
rect 181536 247046 181588 247052
rect 181548 234530 181576 247046
rect 182100 240106 182128 381686
rect 182836 373969 182864 390759
rect 182822 373960 182878 373969
rect 182822 373895 182878 373904
rect 182928 372502 182956 403582
rect 182916 372496 182968 372502
rect 182916 372438 182968 372444
rect 183284 339448 183336 339454
rect 183284 339390 183336 339396
rect 182824 318096 182876 318102
rect 182824 318038 182876 318044
rect 182180 317552 182232 317558
rect 182180 317494 182232 317500
rect 182192 314022 182220 317494
rect 182180 314016 182232 314022
rect 182180 313958 182232 313964
rect 182836 282198 182864 318038
rect 182916 287564 182968 287570
rect 182916 287506 182968 287512
rect 182824 282192 182876 282198
rect 182824 282134 182876 282140
rect 182928 274650 182956 287506
rect 182916 274644 182968 274650
rect 182916 274586 182968 274592
rect 182916 267028 182968 267034
rect 182916 266970 182968 266976
rect 182824 249076 182876 249082
rect 182824 249018 182876 249024
rect 182088 240100 182140 240106
rect 182088 240042 182140 240048
rect 182100 239970 182128 240042
rect 182088 239964 182140 239970
rect 182088 239906 182140 239912
rect 181536 234524 181588 234530
rect 181536 234466 181588 234472
rect 182086 234152 182142 234161
rect 182086 234087 182142 234096
rect 181994 162208 182050 162217
rect 181994 162143 182050 162152
rect 181534 146568 181590 146577
rect 181534 146503 181590 146512
rect 181548 130422 181576 146503
rect 181536 130416 181588 130422
rect 181536 130358 181588 130364
rect 181904 101516 181956 101522
rect 181904 101458 181956 101464
rect 181916 100774 181944 101458
rect 181904 100768 181956 100774
rect 181904 100710 181956 100716
rect 182008 90982 182036 162143
rect 182100 92410 182128 234087
rect 182836 202162 182864 249018
rect 182928 235890 182956 266970
rect 183296 242865 183324 339390
rect 183388 331906 183416 446519
rect 183376 331900 183428 331906
rect 183376 331842 183428 331848
rect 183480 323610 183508 485007
rect 184202 459912 184258 459921
rect 184202 459847 184258 459856
rect 184216 441726 184244 459847
rect 184204 441720 184256 441726
rect 184204 441662 184256 441668
rect 183560 398064 183612 398070
rect 183560 398006 183612 398012
rect 183572 339590 183600 398006
rect 183560 339584 183612 339590
rect 183560 339526 183612 339532
rect 183468 323604 183520 323610
rect 183468 323546 183520 323552
rect 183466 312488 183522 312497
rect 183466 312423 183522 312432
rect 183376 278044 183428 278050
rect 183376 277986 183428 277992
rect 183388 277438 183416 277986
rect 183376 277432 183428 277438
rect 183376 277374 183428 277380
rect 183388 246362 183416 277374
rect 183480 256698 183508 312423
rect 184216 309233 184244 441662
rect 184676 436830 184704 512586
rect 184768 452441 184796 538186
rect 184754 452432 184810 452441
rect 184754 452367 184810 452376
rect 184756 442944 184808 442950
rect 184756 442886 184808 442892
rect 184768 441658 184796 442886
rect 184756 441652 184808 441658
rect 184756 441594 184808 441600
rect 184664 436824 184716 436830
rect 184664 436766 184716 436772
rect 184296 339584 184348 339590
rect 184296 339526 184348 339532
rect 184308 326398 184336 339526
rect 184296 326392 184348 326398
rect 184296 326334 184348 326340
rect 184202 309224 184258 309233
rect 184202 309159 184258 309168
rect 184216 287706 184244 309159
rect 184662 305280 184718 305289
rect 184662 305215 184718 305224
rect 184204 287700 184256 287706
rect 184204 287642 184256 287648
rect 184296 281648 184348 281654
rect 184296 281590 184348 281596
rect 184204 275324 184256 275330
rect 184204 275266 184256 275272
rect 183468 256692 183520 256698
rect 183468 256634 183520 256640
rect 183376 246356 183428 246362
rect 183376 246298 183428 246304
rect 184216 245002 184244 275266
rect 184308 271862 184336 281590
rect 184676 277370 184704 305215
rect 184768 292602 184796 441594
rect 184860 415342 184888 581062
rect 186136 575612 186188 575618
rect 186136 575554 186188 575560
rect 186044 549364 186096 549370
rect 186044 549306 186096 549312
rect 185676 461372 185728 461378
rect 185676 461314 185728 461320
rect 185584 455524 185636 455530
rect 185584 455466 185636 455472
rect 185596 455394 185624 455466
rect 185584 455388 185636 455394
rect 185584 455330 185636 455336
rect 184940 449948 184992 449954
rect 184940 449890 184992 449896
rect 184952 442950 184980 449890
rect 184940 442944 184992 442950
rect 184940 442886 184992 442892
rect 185584 439544 185636 439550
rect 185584 439486 185636 439492
rect 184848 415336 184900 415342
rect 184848 415278 184900 415284
rect 184848 412684 184900 412690
rect 184848 412626 184900 412632
rect 184860 367033 184888 412626
rect 184938 403608 184994 403617
rect 184938 403543 184994 403552
rect 184846 367024 184902 367033
rect 184846 366959 184902 366968
rect 184860 366353 184888 366959
rect 184846 366344 184902 366353
rect 184846 366279 184902 366288
rect 184848 297424 184900 297430
rect 184848 297366 184900 297372
rect 184756 292596 184808 292602
rect 184756 292538 184808 292544
rect 184664 277364 184716 277370
rect 184664 277306 184716 277312
rect 184676 276146 184704 277306
rect 184664 276140 184716 276146
rect 184664 276082 184716 276088
rect 184296 271856 184348 271862
rect 184296 271798 184348 271804
rect 184388 270700 184440 270706
rect 184388 270642 184440 270648
rect 184296 254040 184348 254046
rect 184296 253982 184348 253988
rect 184204 244996 184256 245002
rect 184204 244938 184256 244944
rect 183282 242856 183338 242865
rect 183282 242791 183338 242800
rect 184202 242720 184258 242729
rect 184202 242655 184258 242664
rect 184216 241641 184244 242655
rect 184202 241632 184258 241641
rect 184202 241567 184258 241576
rect 182916 235884 182968 235890
rect 182916 235826 182968 235832
rect 182928 235074 182956 235826
rect 182916 235068 182968 235074
rect 182916 235010 182968 235016
rect 183468 235068 183520 235074
rect 183468 235010 183520 235016
rect 182824 202156 182876 202162
rect 182824 202098 182876 202104
rect 182916 151972 182968 151978
rect 182916 151914 182968 151920
rect 182178 144800 182234 144809
rect 182178 144735 182234 144744
rect 182192 135969 182220 144735
rect 182178 135960 182234 135969
rect 182178 135895 182234 135904
rect 182822 133104 182878 133113
rect 182822 133039 182878 133048
rect 182836 107642 182864 133039
rect 182928 131782 182956 151914
rect 183480 144809 183508 235010
rect 183466 144800 183522 144809
rect 183466 144735 183522 144744
rect 183480 143721 183508 144735
rect 183466 143712 183522 143721
rect 183466 143647 183522 143656
rect 182916 131776 182968 131782
rect 182916 131718 182968 131724
rect 183468 127628 183520 127634
rect 183468 127570 183520 127576
rect 183480 127022 183508 127570
rect 183468 127016 183520 127022
rect 183468 126958 183520 126964
rect 182824 107636 182876 107642
rect 182824 107578 182876 107584
rect 182824 102808 182876 102814
rect 182824 102750 182876 102756
rect 182088 92404 182140 92410
rect 182088 92346 182140 92352
rect 181996 90976 182048 90982
rect 181996 90918 182048 90924
rect 181442 82104 181498 82113
rect 181442 82039 181498 82048
rect 182836 75886 182864 102750
rect 182824 75880 182876 75886
rect 182824 75822 182876 75828
rect 180800 70372 180852 70378
rect 180800 70314 180852 70320
rect 181444 70372 181496 70378
rect 181444 70314 181496 70320
rect 181456 49026 181484 70314
rect 183480 51746 183508 126958
rect 183468 51740 183520 51746
rect 183468 51682 183520 51688
rect 181444 49020 181496 49026
rect 181444 48962 181496 48968
rect 180156 18624 180208 18630
rect 180156 18566 180208 18572
rect 177304 17264 177356 17270
rect 177304 17206 177356 17212
rect 159456 13184 159508 13190
rect 159456 13126 159508 13132
rect 184216 8974 184244 241567
rect 184308 216578 184336 253982
rect 184400 235249 184428 270642
rect 184754 264208 184810 264217
rect 184754 264143 184756 264152
rect 184808 264143 184810 264152
rect 184756 264114 184808 264120
rect 184860 242894 184888 297366
rect 184848 242888 184900 242894
rect 184848 242830 184900 242836
rect 184952 242729 184980 403543
rect 185596 401878 185624 439486
rect 185688 435402 185716 461314
rect 186056 440910 186084 549306
rect 186148 461378 186176 575554
rect 186136 461372 186188 461378
rect 186136 461314 186188 461320
rect 186148 460970 186176 461314
rect 186136 460964 186188 460970
rect 186136 460906 186188 460912
rect 186240 452577 186268 595439
rect 186976 565146 187004 600607
rect 187056 567248 187108 567254
rect 187056 567190 187108 567196
rect 186964 565140 187016 565146
rect 186964 565082 187016 565088
rect 186964 545760 187016 545766
rect 186964 545702 187016 545708
rect 186320 542428 186372 542434
rect 186320 542370 186372 542376
rect 186332 538354 186360 542370
rect 186320 538348 186372 538354
rect 186320 538290 186372 538296
rect 186976 535430 187004 545702
rect 187068 542366 187096 567190
rect 187620 565214 187648 702714
rect 188250 596864 188306 596873
rect 188250 596799 188306 596808
rect 188264 596329 188292 596799
rect 188250 596320 188306 596329
rect 188250 596255 188306 596264
rect 188264 596222 188292 596255
rect 188252 596216 188304 596222
rect 188252 596158 188304 596164
rect 187608 565208 187660 565214
rect 187608 565150 187660 565156
rect 187700 564460 187752 564466
rect 187700 564402 187752 564408
rect 187712 559570 187740 564402
rect 187700 559564 187752 559570
rect 187700 559506 187752 559512
rect 187516 547936 187568 547942
rect 187516 547878 187568 547884
rect 187056 542360 187108 542366
rect 187056 542302 187108 542308
rect 186964 535424 187016 535430
rect 186964 535366 187016 535372
rect 187528 505850 187556 547878
rect 188356 541686 188384 702850
rect 201512 621042 201540 702986
rect 235184 702914 235212 703520
rect 242808 703180 242860 703186
rect 242808 703122 242860 703128
rect 235172 702908 235224 702914
rect 235172 702850 235224 702856
rect 233240 702840 233292 702846
rect 233240 702782 233292 702788
rect 205640 702704 205692 702710
rect 205640 702646 205692 702652
rect 201500 621036 201552 621042
rect 201500 620978 201552 620984
rect 202144 621036 202196 621042
rect 202144 620978 202196 620984
rect 202156 609346 202184 620978
rect 202144 609340 202196 609346
rect 202144 609282 202196 609288
rect 191654 607880 191710 607889
rect 191654 607815 191710 607824
rect 189722 605976 189778 605985
rect 189722 605911 189778 605920
rect 188434 604480 188490 604489
rect 188434 604415 188490 604424
rect 188448 589966 188476 604415
rect 188436 589960 188488 589966
rect 188436 589902 188488 589908
rect 189736 583030 189764 605911
rect 191196 599004 191248 599010
rect 191196 598946 191248 598952
rect 191010 597952 191066 597961
rect 191010 597887 191066 597896
rect 191024 597650 191052 597887
rect 191012 597644 191064 597650
rect 191012 597586 191064 597592
rect 190368 597576 190420 597582
rect 190368 597518 190420 597524
rect 189724 583024 189776 583030
rect 189724 582966 189776 582972
rect 188436 580304 188488 580310
rect 188436 580246 188488 580252
rect 188448 572694 188476 580246
rect 188988 578332 189040 578338
rect 188988 578274 189040 578280
rect 188436 572688 188488 572694
rect 188436 572630 188488 572636
rect 188528 549296 188580 549302
rect 188528 549238 188580 549244
rect 188436 548548 188488 548554
rect 188436 548490 188488 548496
rect 188344 541680 188396 541686
rect 188344 541622 188396 541628
rect 188448 539345 188476 548490
rect 188540 540598 188568 549238
rect 188528 540592 188580 540598
rect 188528 540534 188580 540540
rect 188434 539336 188490 539345
rect 188434 539271 188490 539280
rect 188344 536104 188396 536110
rect 188344 536046 188396 536052
rect 187606 530768 187662 530777
rect 187606 530703 187662 530712
rect 187620 530602 187648 530703
rect 187608 530596 187660 530602
rect 187608 530538 187660 530544
rect 187516 505844 187568 505850
rect 187516 505786 187568 505792
rect 186964 504484 187016 504490
rect 186964 504426 187016 504432
rect 186226 452568 186282 452577
rect 186226 452503 186282 452512
rect 186318 451480 186374 451489
rect 186318 451415 186374 451424
rect 186228 449948 186280 449954
rect 186228 449890 186280 449896
rect 186044 440904 186096 440910
rect 186044 440846 186096 440852
rect 185676 435396 185728 435402
rect 185676 435338 185728 435344
rect 186136 424380 186188 424386
rect 186136 424322 186188 424328
rect 185584 401872 185636 401878
rect 185584 401814 185636 401820
rect 186044 401056 186096 401062
rect 186044 400998 186096 401004
rect 186056 400246 186084 400998
rect 186044 400240 186096 400246
rect 186044 400182 186096 400188
rect 186056 382129 186084 400182
rect 186042 382120 186098 382129
rect 186042 382055 186098 382064
rect 185032 341556 185084 341562
rect 185032 341498 185084 341504
rect 185044 318102 185072 341498
rect 186148 336054 186176 424322
rect 186136 336048 186188 336054
rect 186136 335990 186188 335996
rect 186240 329118 186268 449890
rect 186332 436762 186360 451415
rect 186320 436756 186372 436762
rect 186320 436698 186372 436704
rect 186320 408468 186372 408474
rect 186320 408410 186372 408416
rect 186332 339454 186360 408410
rect 186976 401062 187004 504426
rect 187514 469840 187570 469849
rect 187514 469775 187570 469784
rect 187056 469260 187108 469266
rect 187056 469202 187108 469208
rect 187068 454102 187096 469202
rect 187056 454096 187108 454102
rect 187056 454038 187108 454044
rect 187146 452432 187202 452441
rect 187146 452367 187202 452376
rect 187160 451489 187188 452367
rect 187146 451480 187202 451489
rect 187146 451415 187202 451424
rect 187056 434716 187108 434722
rect 187056 434658 187108 434664
rect 186964 401056 187016 401062
rect 186964 400998 187016 401004
rect 186778 393952 186834 393961
rect 186778 393887 186834 393896
rect 186412 389836 186464 389842
rect 186412 389778 186464 389784
rect 186424 386374 186452 389778
rect 186792 387734 186820 393887
rect 186780 387728 186832 387734
rect 186780 387670 186832 387676
rect 186412 386368 186464 386374
rect 186412 386310 186464 386316
rect 186962 384296 187018 384305
rect 186962 384231 187018 384240
rect 186410 380352 186466 380361
rect 186410 380287 186466 380296
rect 186424 375329 186452 380287
rect 186976 376553 187004 384231
rect 186962 376544 187018 376553
rect 186962 376479 187018 376488
rect 186410 375320 186466 375329
rect 186410 375255 186466 375264
rect 186412 373380 186464 373386
rect 186412 373322 186464 373328
rect 186424 365702 186452 373322
rect 186412 365696 186464 365702
rect 186412 365638 186464 365644
rect 186320 339448 186372 339454
rect 186320 339390 186372 339396
rect 186228 329112 186280 329118
rect 186228 329054 186280 329060
rect 185676 321700 185728 321706
rect 185676 321642 185728 321648
rect 185032 318096 185084 318102
rect 185032 318038 185084 318044
rect 185582 306504 185638 306513
rect 185582 306439 185638 306448
rect 185596 284986 185624 306439
rect 185688 305658 185716 321642
rect 186226 315344 186282 315353
rect 186226 315279 186282 315288
rect 185676 305652 185728 305658
rect 185676 305594 185728 305600
rect 185676 295996 185728 296002
rect 185676 295938 185728 295944
rect 185584 284980 185636 284986
rect 185584 284922 185636 284928
rect 185584 273284 185636 273290
rect 185584 273226 185636 273232
rect 184938 242720 184994 242729
rect 184938 242655 184994 242664
rect 184386 235240 184442 235249
rect 184386 235175 184442 235184
rect 184296 216572 184348 216578
rect 184296 216514 184348 216520
rect 184308 215694 184336 216514
rect 184296 215688 184348 215694
rect 184296 215630 184348 215636
rect 184848 215688 184900 215694
rect 184848 215630 184900 215636
rect 184478 151056 184534 151065
rect 184478 150991 184534 151000
rect 184294 150512 184350 150521
rect 184294 150447 184350 150456
rect 184308 120086 184336 150447
rect 184492 140078 184520 150991
rect 184480 140072 184532 140078
rect 184480 140014 184532 140020
rect 184754 126304 184810 126313
rect 184754 126239 184810 126248
rect 184768 125769 184796 126239
rect 184754 125760 184810 125769
rect 184754 125695 184810 125704
rect 184296 120080 184348 120086
rect 184296 120022 184348 120028
rect 184296 98116 184348 98122
rect 184296 98058 184348 98064
rect 184308 92478 184336 98058
rect 184296 92472 184348 92478
rect 184296 92414 184348 92420
rect 184768 42090 184796 125695
rect 184860 92177 184888 215630
rect 185596 206281 185624 273226
rect 185688 243506 185716 295938
rect 186240 270706 186268 315279
rect 186228 270700 186280 270706
rect 186228 270642 186280 270648
rect 185766 267064 185822 267073
rect 185766 266999 185822 267008
rect 185780 248414 185808 266999
rect 185780 248386 186268 248414
rect 185676 243500 185728 243506
rect 185676 243442 185728 243448
rect 186240 235929 186268 248386
rect 186320 242820 186372 242826
rect 186320 242762 186372 242768
rect 186332 242282 186360 242762
rect 186320 242276 186372 242282
rect 186320 242218 186372 242224
rect 186226 235920 186282 235929
rect 186226 235855 186282 235864
rect 185582 206272 185638 206281
rect 185582 206207 185638 206216
rect 185766 162072 185822 162081
rect 185766 162007 185822 162016
rect 185780 144129 185808 162007
rect 185766 144120 185822 144129
rect 185766 144055 185822 144064
rect 185582 143576 185638 143585
rect 185582 143511 185638 143520
rect 185596 111790 185624 143511
rect 186136 118652 186188 118658
rect 186136 118594 186188 118600
rect 185584 111784 185636 111790
rect 185584 111726 185636 111732
rect 185584 103556 185636 103562
rect 185584 103498 185636 103504
rect 184846 92168 184902 92177
rect 184846 92103 184902 92112
rect 185596 82822 185624 103498
rect 185676 100020 185728 100026
rect 185676 99962 185728 99968
rect 185688 92313 185716 99962
rect 185674 92304 185730 92313
rect 185674 92239 185730 92248
rect 185584 82816 185636 82822
rect 185584 82758 185636 82764
rect 186148 43450 186176 118594
rect 186240 115666 186268 235855
rect 186976 222193 187004 376479
rect 187068 319122 187096 434658
rect 187528 410446 187556 469775
rect 187620 469266 187648 530538
rect 187608 469260 187660 469266
rect 187608 469202 187660 469208
rect 187620 465769 187648 469202
rect 187698 468072 187754 468081
rect 187698 468007 187754 468016
rect 187606 465760 187662 465769
rect 187606 465695 187662 465704
rect 187712 465050 187740 468007
rect 187790 467936 187846 467945
rect 187790 467871 187846 467880
rect 187700 465044 187752 465050
rect 187700 464986 187752 464992
rect 187804 461689 187832 467871
rect 187790 461680 187846 461689
rect 187790 461615 187846 461624
rect 187698 459640 187754 459649
rect 187698 459575 187754 459584
rect 187712 456113 187740 459575
rect 187698 456104 187754 456113
rect 187698 456039 187754 456048
rect 188356 449206 188384 536046
rect 189000 526454 189028 578274
rect 189722 567488 189778 567497
rect 189722 567423 189778 567432
rect 189736 554062 189764 567423
rect 189724 554056 189776 554062
rect 189724 553998 189776 554004
rect 189814 553480 189870 553489
rect 189814 553415 189870 553424
rect 189078 536208 189134 536217
rect 189078 536143 189134 536152
rect 189092 530641 189120 536143
rect 189078 530632 189134 530641
rect 189078 530567 189134 530576
rect 188988 526448 189040 526454
rect 188988 526390 189040 526396
rect 189724 503056 189776 503062
rect 189724 502998 189776 503004
rect 188436 501696 188488 501702
rect 188436 501638 188488 501644
rect 188448 460193 188476 501638
rect 188434 460184 188490 460193
rect 188434 460119 188490 460128
rect 189080 454164 189132 454170
rect 189080 454106 189132 454112
rect 188434 452704 188490 452713
rect 188434 452639 188490 452648
rect 188344 449200 188396 449206
rect 188344 449142 188396 449148
rect 188448 438841 188476 452639
rect 189092 447134 189120 454106
rect 189000 447106 189120 447134
rect 189000 441614 189028 447106
rect 189000 441586 189120 441614
rect 188434 438832 188490 438841
rect 188434 438767 188490 438776
rect 189092 434722 189120 441586
rect 189080 434716 189132 434722
rect 189080 434658 189132 434664
rect 187700 418804 187752 418810
rect 187700 418746 187752 418752
rect 187516 410440 187568 410446
rect 187516 410382 187568 410388
rect 187148 396772 187200 396778
rect 187148 396714 187200 396720
rect 187160 389298 187188 396714
rect 187148 389292 187200 389298
rect 187148 389234 187200 389240
rect 187712 389201 187740 418746
rect 188344 415336 188396 415342
rect 188344 415278 188396 415284
rect 187698 389192 187754 389201
rect 187698 389127 187754 389136
rect 188356 387802 188384 415278
rect 189080 410440 189132 410446
rect 189080 410382 189132 410388
rect 188434 409184 188490 409193
rect 188434 409119 188490 409128
rect 188344 387796 188396 387802
rect 188344 387738 188396 387744
rect 188448 386209 188476 409119
rect 188896 398132 188948 398138
rect 188896 398074 188948 398080
rect 188526 389872 188582 389881
rect 188526 389807 188582 389816
rect 188434 386200 188490 386209
rect 188434 386135 188490 386144
rect 188540 383625 188568 389807
rect 188620 387116 188672 387122
rect 188620 387058 188672 387064
rect 188526 383616 188582 383625
rect 188526 383551 188582 383560
rect 188632 380866 188660 387058
rect 188802 384432 188858 384441
rect 188802 384367 188858 384376
rect 188620 380860 188672 380866
rect 188620 380802 188672 380808
rect 187700 380180 187752 380186
rect 187700 380122 187752 380128
rect 187712 379438 187740 380122
rect 187700 379432 187752 379438
rect 187700 379374 187752 379380
rect 187698 378720 187754 378729
rect 187698 378655 187754 378664
rect 187712 378049 187740 378655
rect 187698 378040 187754 378049
rect 187698 377975 187754 377984
rect 187698 370560 187754 370569
rect 187698 370495 187754 370504
rect 187712 369850 187740 370495
rect 187700 369844 187752 369850
rect 187700 369786 187752 369792
rect 187608 338836 187660 338842
rect 187608 338778 187660 338784
rect 187516 329112 187568 329118
rect 187516 329054 187568 329060
rect 187056 319116 187108 319122
rect 187056 319058 187108 319064
rect 187056 302252 187108 302258
rect 187056 302194 187108 302200
rect 187068 286346 187096 302194
rect 187056 286340 187108 286346
rect 187056 286282 187108 286288
rect 187054 257272 187110 257281
rect 187054 257207 187110 257216
rect 187068 244633 187096 257207
rect 187528 248878 187556 329054
rect 187516 248872 187568 248878
rect 187516 248814 187568 248820
rect 187054 244624 187110 244633
rect 187054 244559 187110 244568
rect 186962 222184 187018 222193
rect 186962 222119 187018 222128
rect 186976 217977 187004 222119
rect 186962 217968 187018 217977
rect 186962 217903 187018 217912
rect 186976 216753 187004 217903
rect 186318 216744 186374 216753
rect 186318 216679 186374 216688
rect 186962 216744 187018 216753
rect 186962 216679 187018 216688
rect 186228 115660 186280 115666
rect 186228 115602 186280 115608
rect 186332 89729 186360 216679
rect 187068 196654 187096 244559
rect 187620 242282 187648 338778
rect 188816 333305 188844 384367
rect 188908 348498 188936 398074
rect 188988 380860 189040 380866
rect 188988 380802 189040 380808
rect 188896 348492 188948 348498
rect 188896 348434 188948 348440
rect 188894 345672 188950 345681
rect 188894 345607 188950 345616
rect 188802 333296 188858 333305
rect 188802 333231 188858 333240
rect 188344 319456 188396 319462
rect 188344 319398 188396 319404
rect 188356 313993 188384 319398
rect 188342 313984 188398 313993
rect 188342 313919 188398 313928
rect 187698 310584 187754 310593
rect 187698 310519 187754 310528
rect 187712 309777 187740 310519
rect 187698 309768 187754 309777
rect 187698 309703 187754 309712
rect 188342 308000 188398 308009
rect 188342 307935 188398 307944
rect 188356 306377 188384 307935
rect 188342 306368 188398 306377
rect 188342 306303 188398 306312
rect 188342 305144 188398 305153
rect 188342 305079 188398 305088
rect 187698 301200 187754 301209
rect 187698 301135 187754 301144
rect 187712 298790 187740 301135
rect 187700 298784 187752 298790
rect 187700 298726 187752 298732
rect 188356 291922 188384 305079
rect 188712 292596 188764 292602
rect 188712 292538 188764 292544
rect 188344 291916 188396 291922
rect 188344 291858 188396 291864
rect 188724 290086 188752 292538
rect 188712 290080 188764 290086
rect 188712 290022 188764 290028
rect 188908 273290 188936 345607
rect 189000 298858 189028 380802
rect 189092 330449 189120 410382
rect 189736 398138 189764 502998
rect 189828 471889 189856 553415
rect 189814 471880 189870 471889
rect 189814 471815 189870 471824
rect 190380 445058 190408 597518
rect 191102 594960 191158 594969
rect 191102 594895 191158 594904
rect 190550 588160 190606 588169
rect 190550 588095 190606 588104
rect 190460 586560 190512 586566
rect 190458 586528 190460 586537
rect 190512 586528 190514 586537
rect 190458 586463 190514 586472
rect 190564 585886 190592 588095
rect 190552 585880 190604 585886
rect 190552 585822 190604 585828
rect 191010 585168 191066 585177
rect 191010 585103 191066 585112
rect 191024 580446 191052 585103
rect 191012 580440 191064 580446
rect 191012 580382 191064 580388
rect 190918 579048 190974 579057
rect 190918 578983 190974 578992
rect 190932 578338 190960 578983
rect 190920 578332 190972 578338
rect 190920 578274 190972 578280
rect 190826 574560 190882 574569
rect 190826 574495 190882 574504
rect 190840 574122 190868 574495
rect 190828 574116 190880 574122
rect 190828 574058 190880 574064
rect 190828 572688 190880 572694
rect 190828 572630 190880 572636
rect 190840 572257 190868 572630
rect 190826 572248 190882 572257
rect 190826 572183 190882 572192
rect 191116 567905 191144 594895
rect 191208 593337 191236 598946
rect 191668 597281 191696 607815
rect 205548 604580 205600 604586
rect 205548 604522 205600 604528
rect 196714 604480 196770 604489
rect 196714 604415 196770 604424
rect 191746 603664 191802 603673
rect 191746 603599 191802 603608
rect 191654 597272 191710 597281
rect 191654 597207 191710 597216
rect 191378 596320 191434 596329
rect 191378 596255 191380 596264
rect 191432 596255 191434 596264
rect 191380 596226 191432 596232
rect 191286 594008 191342 594017
rect 191286 593943 191342 593952
rect 191300 593434 191328 593943
rect 191288 593428 191340 593434
rect 191288 593370 191340 593376
rect 191194 593328 191250 593337
rect 191194 593263 191250 593272
rect 191378 592104 191434 592113
rect 191378 592039 191380 592048
rect 191432 592039 191434 592048
rect 191380 592010 191432 592016
rect 191286 591288 191342 591297
rect 191286 591223 191342 591232
rect 191300 590714 191328 591223
rect 191288 590708 191340 590714
rect 191288 590650 191340 590656
rect 191378 589384 191434 589393
rect 191378 589319 191380 589328
rect 191432 589319 191434 589328
rect 191380 589290 191432 589296
rect 191668 588606 191696 597207
rect 191656 588600 191708 588606
rect 191656 588542 191708 588548
rect 191760 586129 191788 603599
rect 194138 601896 194194 601905
rect 194138 601831 194194 601840
rect 194152 600953 194180 601831
rect 194138 600944 194194 600953
rect 194138 600879 194194 600888
rect 192574 600808 192630 600817
rect 192574 600743 192630 600752
rect 192484 600364 192536 600370
rect 192484 600306 192536 600312
rect 192496 587178 192524 600306
rect 192588 592686 192616 600743
rect 195428 600364 195480 600370
rect 195428 600306 195480 600312
rect 192666 599448 192722 599457
rect 192666 599383 192722 599392
rect 192680 595474 192708 599383
rect 195440 599148 195468 600306
rect 196728 599148 196756 604415
rect 199108 603220 199160 603226
rect 199108 603162 199160 603168
rect 198554 599448 198610 599457
rect 198554 599383 198610 599392
rect 198568 599148 198596 599383
rect 199120 599148 199148 603162
rect 201130 602032 201186 602041
rect 201130 601967 201186 601976
rect 199842 600672 199898 600681
rect 199842 600607 199898 600616
rect 199856 599148 199884 600607
rect 200396 600432 200448 600438
rect 200396 600374 200448 600380
rect 200408 599148 200436 600374
rect 201144 599148 201172 601967
rect 204810 601896 204866 601905
rect 204810 601831 204866 601840
rect 204258 600808 204314 600817
rect 204258 600743 204314 600752
rect 202418 600672 202474 600681
rect 202418 600607 202474 600616
rect 202432 599148 202460 600607
rect 204272 599162 204300 600743
rect 204442 599176 204498 599185
rect 204272 599148 204442 599162
rect 193404 599140 193456 599146
rect 193126 599108 193182 599117
rect 204286 599134 204442 599148
rect 204824 599148 204852 601831
rect 205560 599148 205588 604522
rect 205652 599593 205680 702646
rect 215300 702636 215352 702642
rect 215300 702578 215352 702584
rect 222844 702636 222896 702642
rect 222844 702578 222896 702584
rect 213184 611448 213236 611454
rect 213184 611390 213236 611396
rect 213092 610088 213144 610094
rect 207662 610056 207718 610065
rect 213092 610030 213144 610036
rect 207662 609991 207718 610000
rect 205732 608660 205784 608666
rect 205732 608602 205784 608608
rect 205638 599584 205694 599593
rect 205638 599519 205694 599528
rect 205744 599162 205772 608602
rect 206834 599584 206890 599593
rect 206834 599519 206890 599528
rect 205744 599134 206126 599162
rect 206848 599148 206876 599519
rect 207676 599162 207704 609991
rect 208398 608832 208454 608841
rect 208398 608767 208454 608776
rect 208412 599162 208440 608767
rect 209410 607336 209466 607345
rect 209410 607271 209466 607280
rect 207676 599134 208150 599162
rect 208412 599134 208702 599162
rect 209424 599148 209452 607271
rect 212540 605940 212592 605946
rect 212540 605882 212592 605888
rect 211252 601724 211304 601730
rect 211252 601666 211304 601672
rect 209962 600808 210018 600817
rect 209962 600743 210018 600752
rect 209976 599148 210004 600743
rect 211264 599148 211292 601666
rect 211804 601656 211856 601662
rect 211804 601598 211856 601604
rect 211816 599148 211844 601598
rect 212448 600364 212500 600370
rect 212448 600306 212500 600312
rect 212460 599457 212488 600306
rect 212446 599448 212502 599457
rect 212446 599383 212502 599392
rect 212552 599148 212580 605882
rect 213104 599298 213132 610030
rect 213196 601662 213224 611390
rect 214380 603152 214432 603158
rect 214380 603094 214432 603100
rect 213184 601656 213236 601662
rect 213184 601598 213236 601604
rect 213104 599270 213408 599298
rect 213274 599176 213330 599185
rect 213118 599134 213274 599162
rect 204442 599111 204498 599120
rect 213380 599162 213408 599270
rect 213380 599134 213854 599162
rect 214392 599148 214420 603094
rect 215312 600409 215340 702578
rect 222856 615494 222884 702578
rect 224224 702568 224276 702574
rect 224224 702510 224276 702516
rect 222856 615466 222976 615494
rect 215944 614236 215996 614242
rect 215944 614178 215996 614184
rect 215956 607170 215984 614178
rect 219348 609272 219400 609278
rect 219348 609214 219400 609220
rect 217692 607300 217744 607306
rect 217692 607242 217744 607248
rect 216956 607232 217008 607238
rect 216956 607174 217008 607180
rect 215944 607164 215996 607170
rect 215944 607106 215996 607112
rect 215298 600400 215354 600409
rect 215298 600335 215354 600344
rect 215956 599162 215984 607106
rect 216402 600400 216458 600409
rect 216402 600335 216458 600344
rect 215694 599134 215984 599162
rect 216416 599148 216444 600335
rect 216968 599148 216996 607174
rect 217704 599148 217732 607242
rect 218796 607232 218848 607238
rect 218796 607174 218848 607180
rect 218242 600400 218298 600409
rect 218242 600335 218298 600344
rect 218256 599148 218284 600335
rect 218808 599148 218836 607174
rect 219360 600409 219388 609214
rect 222106 605976 222162 605985
rect 222106 605911 222162 605920
rect 221372 600840 221424 600846
rect 221372 600782 221424 600788
rect 219346 600400 219402 600409
rect 219346 600335 219402 600344
rect 219532 600364 219584 600370
rect 219532 600306 219584 600312
rect 219544 599148 219572 600306
rect 221384 599148 221412 600782
rect 222120 599148 222148 605911
rect 222948 600545 222976 615466
rect 223028 609340 223080 609346
rect 223028 609282 223080 609288
rect 222934 600536 222990 600545
rect 222934 600471 222990 600480
rect 222660 599480 222712 599486
rect 222660 599422 222712 599428
rect 222672 599162 222700 599422
rect 222948 599162 222976 600471
rect 223040 599486 223068 609282
rect 224236 601662 224264 702510
rect 227718 619712 227774 619721
rect 227718 619647 227774 619656
rect 226340 618316 226392 618322
rect 226340 618258 226392 618264
rect 226352 615494 226380 618258
rect 226352 615466 226656 615494
rect 226430 608696 226486 608705
rect 226430 608631 226486 608640
rect 226338 603120 226394 603129
rect 226338 603055 226394 603064
rect 224224 601656 224276 601662
rect 224224 601598 224276 601604
rect 225236 601656 225288 601662
rect 225236 601598 225288 601604
rect 223028 599480 223080 599486
rect 223028 599422 223080 599428
rect 222672 599148 222884 599162
rect 222686 599134 222884 599148
rect 222948 599134 223422 599162
rect 225248 599148 225276 601598
rect 226352 600846 226380 603055
rect 226340 600840 226392 600846
rect 226340 600782 226392 600788
rect 225786 600400 225842 600409
rect 225786 600335 225842 600344
rect 226340 600364 226392 600370
rect 225800 599148 225828 600335
rect 226340 600306 226392 600312
rect 226352 599457 226380 600306
rect 226338 599448 226394 599457
rect 226338 599383 226394 599392
rect 226444 599162 226472 608631
rect 226628 599162 226656 615466
rect 227732 599162 227760 619647
rect 233252 616010 233280 702782
rect 233240 616004 233292 616010
rect 233240 615946 233292 615952
rect 233884 616004 233936 616010
rect 233884 615946 233936 615952
rect 233252 615602 233280 615946
rect 233240 615596 233292 615602
rect 233240 615538 233292 615544
rect 231860 615528 231912 615534
rect 231912 615476 232360 615494
rect 231860 615470 232360 615476
rect 231872 615466 232360 615470
rect 230110 603256 230166 603265
rect 230110 603191 230166 603200
rect 230124 601905 230152 603191
rect 230110 601896 230166 601905
rect 230032 601854 230110 601882
rect 229100 601792 229152 601798
rect 229100 601734 229152 601740
rect 226444 599134 226550 599162
rect 226628 599134 227102 599162
rect 227732 599134 227838 599162
rect 229112 599148 229140 601734
rect 230032 599162 230060 601854
rect 230110 601831 230166 601840
rect 231766 600536 231822 600545
rect 231766 600471 231822 600480
rect 231780 600370 231808 600471
rect 231768 600364 231820 600370
rect 231768 600306 231820 600312
rect 232228 600364 232280 600370
rect 232228 600306 232280 600312
rect 229678 599134 230060 599162
rect 231214 599176 231270 599185
rect 213274 599111 213330 599120
rect 193404 599082 193456 599088
rect 193126 599043 193182 599052
rect 192668 595468 192720 595474
rect 192668 595410 192720 595416
rect 193034 593464 193090 593473
rect 193034 593399 193090 593408
rect 192576 592680 192628 592686
rect 192576 592622 192628 592628
rect 192484 587172 192536 587178
rect 192484 587114 192536 587120
rect 191746 586120 191802 586129
rect 191746 586055 191802 586064
rect 191760 585818 191788 586055
rect 191748 585812 191800 585818
rect 191748 585754 191800 585760
rect 191746 583944 191802 583953
rect 191746 583879 191802 583888
rect 191760 583778 191788 583879
rect 191748 583772 191800 583778
rect 191748 583714 191800 583720
rect 191286 582720 191342 582729
rect 191286 582655 191342 582664
rect 191194 581768 191250 581777
rect 191194 581703 191250 581712
rect 191208 581126 191236 581703
rect 191196 581120 191248 581126
rect 191196 581062 191248 581068
rect 191300 574802 191328 582655
rect 191746 581224 191802 581233
rect 191746 581159 191802 581168
rect 191760 581058 191788 581159
rect 191748 581052 191800 581058
rect 191748 580994 191800 581000
rect 191562 579728 191618 579737
rect 191562 579663 191618 579672
rect 191576 578921 191604 579663
rect 191562 578912 191618 578921
rect 191562 578847 191618 578856
rect 191654 578368 191710 578377
rect 191654 578303 191710 578312
rect 191668 578270 191696 578303
rect 191656 578264 191708 578270
rect 191656 578206 191708 578212
rect 191748 578196 191800 578202
rect 191748 578138 191800 578144
rect 191760 578105 191788 578138
rect 191746 578096 191802 578105
rect 191746 578031 191802 578040
rect 191654 576192 191710 576201
rect 191654 576127 191710 576136
rect 191668 575618 191696 576127
rect 191746 575648 191802 575657
rect 191656 575612 191708 575618
rect 191746 575583 191802 575592
rect 191656 575554 191708 575560
rect 191760 575550 191788 575583
rect 191748 575544 191800 575550
rect 191748 575486 191800 575492
rect 191288 574796 191340 574802
rect 191288 574738 191340 574744
rect 191746 572792 191802 572801
rect 191746 572727 191748 572736
rect 191800 572727 191802 572736
rect 191748 572698 191800 572704
rect 191746 570888 191802 570897
rect 191746 570823 191802 570832
rect 191760 570654 191788 570823
rect 191748 570648 191800 570654
rect 191748 570590 191800 570596
rect 191746 570072 191802 570081
rect 191746 570007 191802 570016
rect 191760 569974 191788 570007
rect 191748 569968 191800 569974
rect 191748 569910 191800 569916
rect 191102 567896 191158 567905
rect 191102 567831 191158 567840
rect 191380 567248 191432 567254
rect 191378 567216 191380 567225
rect 191432 567216 191434 567225
rect 191378 567151 191434 567160
rect 191748 565208 191800 565214
rect 191286 565176 191342 565185
rect 191748 565150 191800 565156
rect 191286 565111 191342 565120
rect 191300 564466 191328 565111
rect 191760 565049 191788 565150
rect 191746 565040 191802 565049
rect 191746 564975 191802 564984
rect 191288 564460 191340 564466
rect 191288 564402 191340 564408
rect 191748 563712 191800 563718
rect 191746 563680 191748 563689
rect 191800 563680 191802 563689
rect 191746 563615 191802 563624
rect 190918 562184 190974 562193
rect 190918 562119 190974 562128
rect 190932 561746 190960 562119
rect 190920 561740 190972 561746
rect 190920 561682 190972 561688
rect 190826 560960 190882 560969
rect 190826 560895 190882 560904
rect 190840 560318 190868 560895
rect 190828 560312 190880 560318
rect 190828 560254 190880 560260
rect 191746 559192 191802 559201
rect 191746 559127 191802 559136
rect 191760 558958 191788 559127
rect 191748 558952 191800 558958
rect 191748 558894 191800 558900
rect 191746 557832 191802 557841
rect 191746 557767 191802 557776
rect 191760 557598 191788 557767
rect 191748 557592 191800 557598
rect 191748 557534 191800 557540
rect 191746 556472 191802 556481
rect 191746 556407 191802 556416
rect 191760 556238 191788 556407
rect 191748 556232 191800 556238
rect 191748 556174 191800 556180
rect 191470 554976 191526 554985
rect 191470 554911 191526 554920
rect 191484 554878 191512 554911
rect 191472 554872 191524 554878
rect 191472 554814 191524 554820
rect 191102 552664 191158 552673
rect 191102 552599 191158 552608
rect 191116 552158 191144 552599
rect 191104 552152 191156 552158
rect 191104 552094 191156 552100
rect 191746 550760 191802 550769
rect 191746 550695 191802 550704
rect 191760 550662 191788 550695
rect 191748 550656 191800 550662
rect 191748 550598 191800 550604
rect 191654 549808 191710 549817
rect 191654 549743 191710 549752
rect 190642 548312 190698 548321
rect 190642 548247 190698 548256
rect 190656 547942 190684 548247
rect 190644 547936 190696 547942
rect 190644 547878 190696 547884
rect 191668 547874 191696 549743
rect 191746 549400 191802 549409
rect 191746 549335 191748 549344
rect 191800 549335 191802 549344
rect 191748 549306 191800 549312
rect 191668 547846 191788 547874
rect 191562 547088 191618 547097
rect 191562 547023 191618 547032
rect 191576 546514 191604 547023
rect 191656 546576 191708 546582
rect 191654 546544 191656 546553
rect 191708 546544 191710 546553
rect 191564 546508 191616 546514
rect 191654 546479 191710 546488
rect 191564 546450 191616 546456
rect 191654 545320 191710 545329
rect 191654 545255 191710 545264
rect 191668 545154 191696 545255
rect 191656 545148 191708 545154
rect 191656 545090 191708 545096
rect 191564 545080 191616 545086
rect 191564 545022 191616 545028
rect 191010 544232 191066 544241
rect 191010 544167 191066 544176
rect 191024 543794 191052 544167
rect 191576 544105 191604 545022
rect 191562 544096 191618 544105
rect 191562 544031 191618 544040
rect 191012 543788 191064 543794
rect 191012 543730 191064 543736
rect 191656 540592 191708 540598
rect 191654 540560 191656 540569
rect 191708 540560 191710 540569
rect 191654 540495 191710 540504
rect 191654 456240 191710 456249
rect 191654 456175 191710 456184
rect 191562 456104 191618 456113
rect 191562 456039 191618 456048
rect 190458 449168 190514 449177
rect 190458 449103 190514 449112
rect 190472 448526 190500 449103
rect 190460 448520 190512 448526
rect 190460 448462 190512 448468
rect 191576 447817 191604 456039
rect 191562 447808 191618 447817
rect 191562 447743 191618 447752
rect 191564 447092 191616 447098
rect 191564 447034 191616 447040
rect 191576 446457 191604 447034
rect 191562 446448 191618 446457
rect 191562 446383 191618 446392
rect 191562 445088 191618 445097
rect 190368 445052 190420 445058
rect 191562 445023 191564 445032
rect 190368 444994 190420 445000
rect 191616 445023 191618 445032
rect 191564 444994 191616 445000
rect 191378 442096 191434 442105
rect 191378 442031 191434 442040
rect 191392 441658 191420 442031
rect 191380 441652 191432 441658
rect 191668 441614 191696 456175
rect 191380 441594 191432 441600
rect 191484 441586 191696 441614
rect 190644 440904 190696 440910
rect 190644 440846 190696 440852
rect 190656 440745 190684 440846
rect 190642 440736 190698 440745
rect 190642 440671 190698 440680
rect 190644 438184 190696 438190
rect 190644 438126 190696 438132
rect 190656 438025 190684 438126
rect 190642 438016 190698 438025
rect 190642 437951 190698 437960
rect 191484 433945 191512 441586
rect 191656 440224 191708 440230
rect 191656 440166 191708 440172
rect 191668 439385 191696 440166
rect 191654 439376 191710 439385
rect 191654 439311 191710 439320
rect 191656 436824 191708 436830
rect 191562 436792 191618 436801
rect 191656 436766 191708 436772
rect 191562 436727 191618 436736
rect 191576 435305 191604 436727
rect 191668 436665 191696 436766
rect 191654 436656 191710 436665
rect 191654 436591 191710 436600
rect 191562 435296 191618 435305
rect 191562 435231 191618 435240
rect 191470 433936 191526 433945
rect 191470 433871 191526 433880
rect 191654 432304 191710 432313
rect 191654 432239 191710 432248
rect 191668 432002 191696 432239
rect 191656 431996 191708 432002
rect 191656 431938 191708 431944
rect 191760 431254 191788 547846
rect 193048 530602 193076 593399
rect 193036 530596 193088 530602
rect 193036 530538 193088 530544
rect 193140 527950 193168 599043
rect 193416 584458 193444 599082
rect 197636 599072 197688 599078
rect 194598 599040 194654 599049
rect 193508 598998 194166 599026
rect 193508 598505 193536 598998
rect 197174 599040 197230 599049
rect 194654 598998 194718 599026
rect 195624 599010 196006 599026
rect 195612 599004 196006 599010
rect 194598 598975 194654 598984
rect 195664 598998 196006 599004
rect 197230 598998 197294 599026
rect 201590 599040 201646 599049
rect 197688 599020 198030 599026
rect 197636 599014 198030 599020
rect 197648 598998 198030 599014
rect 197174 598975 197230 598984
rect 203062 599040 203118 599049
rect 201646 598998 201710 599026
rect 202998 598998 203062 599026
rect 201590 598975 201646 598984
rect 207110 599040 207166 599049
rect 203062 598975 203118 598984
rect 203352 598998 203734 599026
rect 195612 598946 195664 598952
rect 203352 598942 203380 598998
rect 210790 599040 210846 599049
rect 207166 598998 207414 599026
rect 210726 598998 210790 599026
rect 207110 598975 207166 598984
rect 219714 599040 219770 599049
rect 214760 599010 215142 599026
rect 210790 598975 210846 598984
rect 214748 599004 215142 599010
rect 214800 598998 215142 599004
rect 220910 599040 220966 599049
rect 219770 598998 220110 599026
rect 220846 598998 220910 599026
rect 219714 598975 219770 598984
rect 222856 599010 222884 599134
rect 231270 599134 231518 599162
rect 232240 599148 232268 600306
rect 232332 599162 232360 615466
rect 233896 600710 233924 615946
rect 237472 612876 237524 612882
rect 237472 612818 237524 612824
rect 234066 604616 234122 604625
rect 234066 604551 234122 604560
rect 233884 600704 233936 600710
rect 233884 600646 233936 600652
rect 232332 599134 232806 599162
rect 234080 599148 234108 604551
rect 235356 600704 235408 600710
rect 235356 600646 235408 600652
rect 235368 599148 235396 600646
rect 236366 599448 236422 599457
rect 236366 599383 236422 599392
rect 236380 599162 236408 599383
rect 236826 599176 236882 599185
rect 236118 599134 236408 599162
rect 236670 599134 236826 599162
rect 231214 599111 231270 599120
rect 237484 599162 237512 612818
rect 242820 604518 242848 703122
rect 249708 702908 249760 702914
rect 249708 702850 249760 702856
rect 242900 616888 242952 616894
rect 242900 616830 242952 616836
rect 238484 604512 238536 604518
rect 238484 604454 238536 604460
rect 241796 604512 241848 604518
rect 241796 604454 241848 604460
rect 242808 604512 242860 604518
rect 242808 604454 242860 604460
rect 237484 599134 237958 599162
rect 238496 599148 238524 604454
rect 241060 601792 241112 601798
rect 239218 601760 239274 601769
rect 241060 601734 241112 601740
rect 239218 601695 239274 601704
rect 239232 599148 239260 601695
rect 240046 599176 240102 599185
rect 239798 599134 240046 599162
rect 236826 599111 236882 599120
rect 241072 599148 241100 601734
rect 241808 599148 241836 604454
rect 242912 599162 242940 616830
rect 245476 605872 245528 605878
rect 245476 605814 245528 605820
rect 244924 603220 244976 603226
rect 244924 603162 244976 603168
rect 244186 600672 244242 600681
rect 244186 600607 244242 600616
rect 243910 599176 243966 599185
rect 242912 599134 243110 599162
rect 243662 599134 243910 599162
rect 240046 599111 240102 599120
rect 244200 599148 244228 600607
rect 244936 599148 244964 603162
rect 245488 599148 245516 605814
rect 249720 603158 249748 702850
rect 255964 702568 256016 702574
rect 255964 702510 256016 702516
rect 251824 700324 251876 700330
rect 251824 700266 251876 700272
rect 251836 615494 251864 700266
rect 251836 615466 251956 615494
rect 251928 614174 251956 615466
rect 251916 614168 251968 614174
rect 251916 614110 251968 614116
rect 249708 603152 249760 603158
rect 249708 603094 249760 603100
rect 246210 600536 246266 600545
rect 246210 600471 246266 600480
rect 246762 600536 246818 600545
rect 246762 600471 246818 600480
rect 246224 599148 246252 600471
rect 246776 599148 246804 600471
rect 248328 600364 248380 600370
rect 248328 600306 248380 600312
rect 248340 599593 248368 600306
rect 248326 599584 248382 599593
rect 248326 599519 248382 599528
rect 249338 599312 249394 599321
rect 249338 599247 249394 599256
rect 249352 599162 249380 599247
rect 249720 599162 249748 603094
rect 250074 600400 250130 600409
rect 250074 600335 250130 600344
rect 249352 599148 249748 599162
rect 250088 599148 250116 600335
rect 251928 599148 251956 614110
rect 254124 611380 254176 611386
rect 254124 611322 254176 611328
rect 253124 599270 253428 599298
rect 253124 599162 253152 599270
rect 249366 599134 249748 599148
rect 252494 599134 253152 599162
rect 243910 599111 243966 599120
rect 228640 599072 228692 599078
rect 223854 599040 223910 599049
rect 220910 598975 220966 598984
rect 222844 599004 222896 599010
rect 214748 598946 214800 598952
rect 224222 599040 224278 599049
rect 223910 598998 223974 599026
rect 223854 598975 223910 598984
rect 224278 598998 224526 599026
rect 228390 599020 228640 599026
rect 251456 599072 251508 599078
rect 228390 599014 228692 599020
rect 230018 599040 230074 599049
rect 228390 598998 228680 599014
rect 224222 598975 224278 598984
rect 230662 599040 230718 599049
rect 230074 598998 230414 599026
rect 230018 598975 230074 598984
rect 233238 599040 233294 599049
rect 230718 598998 230966 599026
rect 230662 598975 230718 598984
rect 234710 599040 234766 599049
rect 233294 598998 233542 599026
rect 233238 598975 233294 598984
rect 236826 599040 236882 599049
rect 234766 598998 234830 599026
rect 234710 598975 234766 598984
rect 240690 599040 240746 599049
rect 236882 598998 237222 599026
rect 240534 598998 240690 599026
rect 236826 598975 236882 598984
rect 242622 599040 242678 599049
rect 242374 598998 242622 599026
rect 240690 598975 240746 598984
rect 247774 599040 247830 599049
rect 247526 598998 247724 599026
rect 242622 598975 242678 598984
rect 222844 598946 222896 598952
rect 247696 598942 247724 598998
rect 250258 599040 250314 599049
rect 247830 598998 248078 599026
rect 248814 598998 249104 599026
rect 247774 598975 247830 598984
rect 249076 598942 249104 598998
rect 250314 598998 250654 599026
rect 251206 599020 251456 599026
rect 253296 599072 253348 599078
rect 251206 599014 251508 599020
rect 252834 599040 252890 599049
rect 251206 598998 251496 599014
rect 250258 598975 250314 598984
rect 252890 598998 253230 599026
rect 253296 599014 253348 599020
rect 252834 598975 252890 598984
rect 203340 598936 203392 598942
rect 203340 598878 203392 598884
rect 247684 598936 247736 598942
rect 247684 598878 247736 598884
rect 249064 598936 249116 598942
rect 249064 598878 249116 598884
rect 193494 598496 193550 598505
rect 193494 598431 193550 598440
rect 253308 592034 253336 599014
rect 253400 596834 253428 599270
rect 253480 598936 253532 598942
rect 253480 598878 253532 598884
rect 253492 597582 253520 598878
rect 253480 597576 253532 597582
rect 253480 597518 253532 597524
rect 253388 596828 253440 596834
rect 253388 596770 253440 596776
rect 253938 592308 253994 592317
rect 253938 592243 253994 592252
rect 253308 592006 253428 592034
rect 253400 591326 253428 592006
rect 253388 591320 253440 591326
rect 253388 591262 253440 591268
rect 193404 584452 193456 584458
rect 193404 584394 193456 584400
rect 253386 556200 253442 556209
rect 253386 556135 253442 556144
rect 253400 547874 253428 556135
rect 253308 547846 253428 547874
rect 251456 539368 251508 539374
rect 251456 539310 251508 539316
rect 250444 539300 250496 539306
rect 250444 539242 250496 539248
rect 193600 536217 193628 539172
rect 193586 536208 193642 536217
rect 193586 536143 193642 536152
rect 194152 536081 194180 539172
rect 194612 539158 194718 539186
rect 194138 536072 194194 536081
rect 194138 536007 194194 536016
rect 193128 527944 193180 527950
rect 193128 527886 193180 527892
rect 193312 526448 193364 526454
rect 193312 526390 193364 526396
rect 193128 514140 193180 514146
rect 193128 514082 193180 514088
rect 192576 497480 192628 497486
rect 192576 497422 192628 497428
rect 192484 480956 192536 480962
rect 192484 480898 192536 480904
rect 191932 449744 191984 449750
rect 191932 449686 191984 449692
rect 191944 448497 191972 449686
rect 191930 448488 191986 448497
rect 191840 448452 191892 448458
rect 191930 448423 191986 448432
rect 191840 448394 191892 448400
rect 191852 443601 191880 448394
rect 191838 443592 191894 443601
rect 191838 443527 191894 443536
rect 191748 431248 191800 431254
rect 191748 431190 191800 431196
rect 191760 430953 191788 431190
rect 191746 430944 191802 430953
rect 191746 430879 191802 430888
rect 191012 430568 191064 430574
rect 191012 430510 191064 430516
rect 191024 429593 191052 430510
rect 191010 429584 191066 429593
rect 191010 429519 191066 429528
rect 190828 429140 190880 429146
rect 190828 429082 190880 429088
rect 190840 428233 190868 429082
rect 190826 428224 190882 428233
rect 190826 428159 190882 428168
rect 190828 427780 190880 427786
rect 190828 427722 190880 427728
rect 190840 426873 190868 427722
rect 190826 426864 190882 426873
rect 190826 426799 190882 426808
rect 191748 425740 191800 425746
rect 191748 425682 191800 425688
rect 191760 425513 191788 425682
rect 191746 425504 191802 425513
rect 191746 425439 191802 425448
rect 191748 424380 191800 424386
rect 191748 424322 191800 424328
rect 191760 423881 191788 424322
rect 191746 423872 191802 423881
rect 191746 423807 191802 423816
rect 191012 423632 191064 423638
rect 191012 423574 191064 423580
rect 191024 422521 191052 423574
rect 191010 422512 191066 422521
rect 191010 422447 191066 422456
rect 191746 421152 191802 421161
rect 191746 421087 191802 421096
rect 191760 420918 191788 421087
rect 192496 420986 192524 480898
rect 192588 475561 192616 497422
rect 192574 475552 192630 475561
rect 192574 475487 192630 475496
rect 193036 464364 193088 464370
rect 193036 464306 193088 464312
rect 193048 443737 193076 464306
rect 193034 443728 193090 443737
rect 193034 443663 193090 443672
rect 193048 443018 193076 443663
rect 193036 443012 193088 443018
rect 193036 442954 193088 442960
rect 192484 420980 192536 420986
rect 192484 420922 192536 420928
rect 191748 420912 191800 420918
rect 191748 420854 191800 420860
rect 192496 419801 192524 420922
rect 192482 419792 192538 419801
rect 192482 419727 192538 419736
rect 191748 419484 191800 419490
rect 191748 419426 191800 419432
rect 191760 418441 191788 419426
rect 191746 418432 191802 418441
rect 191746 418367 191802 418376
rect 191746 417072 191802 417081
rect 191746 417007 191802 417016
rect 191760 416838 191788 417007
rect 191748 416832 191800 416838
rect 191748 416774 191800 416780
rect 190644 416084 190696 416090
rect 190644 416026 190696 416032
rect 190656 415449 190684 416026
rect 190642 415440 190698 415449
rect 190642 415375 190698 415384
rect 191472 415404 191524 415410
rect 191472 415346 191524 415352
rect 191484 414089 191512 415346
rect 191470 414080 191526 414089
rect 191470 414015 191526 414024
rect 191746 412720 191802 412729
rect 191746 412655 191748 412664
rect 191800 412655 191802 412664
rect 191748 412626 191800 412632
rect 193140 411369 193168 514082
rect 193324 460934 193352 526390
rect 194612 515409 194640 539158
rect 195440 532030 195468 539172
rect 195992 533458 196020 539172
rect 196176 539158 196742 539186
rect 195980 533452 196032 533458
rect 195980 533394 196032 533400
rect 195428 532024 195480 532030
rect 195428 531966 195480 531972
rect 196176 528554 196204 539158
rect 197280 535537 197308 539172
rect 197266 535528 197322 535537
rect 197266 535463 197322 535472
rect 198016 535362 198044 539172
rect 198200 539158 198582 539186
rect 198752 539158 199318 539186
rect 198200 538214 198228 539158
rect 198108 538186 198228 538214
rect 198004 535356 198056 535362
rect 198004 535298 198056 535304
rect 198108 533338 198136 538186
rect 195992 528526 196204 528554
rect 197372 533310 198136 533338
rect 195992 525162 196020 528526
rect 195980 525156 196032 525162
rect 195980 525098 196032 525104
rect 195244 522300 195296 522306
rect 195244 522242 195296 522248
rect 194598 515400 194654 515409
rect 194598 515335 194654 515344
rect 193324 460906 193536 460934
rect 193508 456794 193536 460906
rect 195058 458960 195114 458969
rect 195058 458895 195114 458904
rect 195072 456822 195100 458895
rect 193416 456766 193536 456794
rect 194600 456816 194652 456822
rect 193416 448458 193444 456766
rect 194600 456758 194652 456764
rect 195060 456816 195112 456822
rect 195060 456758 195112 456764
rect 193588 454096 193640 454102
rect 193588 454038 193640 454044
rect 193600 450228 193628 454038
rect 194612 450242 194640 456758
rect 194612 450214 194718 450242
rect 195256 449993 195284 522242
rect 197372 512689 197400 533310
rect 198002 530632 198058 530641
rect 198002 530567 198058 530576
rect 197358 512680 197414 512689
rect 197358 512615 197414 512624
rect 195334 511456 195390 511465
rect 195334 511391 195390 511400
rect 195348 461553 195376 511391
rect 198016 503033 198044 530567
rect 198096 511284 198148 511290
rect 198096 511226 198148 511232
rect 198002 503024 198058 503033
rect 198002 502959 198058 502968
rect 196624 492040 196676 492046
rect 196624 491982 196676 491988
rect 195334 461544 195390 461553
rect 195334 461479 195390 461488
rect 196636 459105 196664 491982
rect 198108 490686 198136 511226
rect 198096 490680 198148 490686
rect 198096 490622 198148 490628
rect 198752 487830 198780 539158
rect 199856 534041 199884 539172
rect 200408 538218 200436 539172
rect 200592 539158 201158 539186
rect 201604 539158 201710 539186
rect 202064 539158 202446 539186
rect 200396 538212 200448 538218
rect 200396 538154 200448 538160
rect 199842 534032 199898 534041
rect 199842 533967 199898 533976
rect 198832 533452 198884 533458
rect 198832 533394 198884 533400
rect 198844 488510 198872 533394
rect 200212 530596 200264 530602
rect 200212 530538 200264 530544
rect 199384 523728 199436 523734
rect 199384 523670 199436 523676
rect 198832 488504 198884 488510
rect 198832 488446 198884 488452
rect 198844 487898 198872 488446
rect 198832 487892 198884 487898
rect 198832 487834 198884 487840
rect 198740 487824 198792 487830
rect 198740 487766 198792 487772
rect 196714 482216 196770 482225
rect 196714 482151 196770 482160
rect 196622 459096 196678 459105
rect 196622 459031 196678 459040
rect 196728 456385 196756 482151
rect 197358 465760 197414 465769
rect 197358 465695 197414 465704
rect 197372 463758 197400 465695
rect 197360 463752 197412 463758
rect 197360 463694 197412 463700
rect 196714 456376 196770 456385
rect 196714 456311 196770 456320
rect 196072 455524 196124 455530
rect 196072 455466 196124 455472
rect 195610 452704 195666 452713
rect 195610 452639 195666 452648
rect 195624 450228 195652 452639
rect 196084 450242 196112 455466
rect 197372 450242 197400 463694
rect 197910 454064 197966 454073
rect 197910 453999 197966 454008
rect 197924 450242 197952 453999
rect 199292 452600 199344 452606
rect 199292 452542 199344 452548
rect 199304 451382 199332 452542
rect 199292 451376 199344 451382
rect 199292 451318 199344 451324
rect 196084 450214 196558 450242
rect 197372 450214 197478 450242
rect 197924 450214 198398 450242
rect 199304 450228 199332 451318
rect 199396 450401 199424 523670
rect 199476 487824 199528 487830
rect 199476 487766 199528 487772
rect 199488 452606 199516 487766
rect 200224 452674 200252 530538
rect 200592 528554 200620 539158
rect 201500 532772 201552 532778
rect 201500 532714 201552 532720
rect 200316 528526 200620 528554
rect 200316 490618 200344 528526
rect 200304 490612 200356 490618
rect 200304 490554 200356 490560
rect 201512 461514 201540 532714
rect 201604 527882 201632 539158
rect 202064 532778 202092 539158
rect 202984 538121 203012 539172
rect 203352 539158 203734 539186
rect 204286 539158 204484 539186
rect 202970 538112 203026 538121
rect 202970 538047 203026 538056
rect 202052 532772 202104 532778
rect 202052 532714 202104 532720
rect 202984 532030 203012 538047
rect 202972 532024 203024 532030
rect 202972 531966 203024 531972
rect 203352 530641 203380 539158
rect 203338 530632 203394 530641
rect 203338 530567 203394 530576
rect 201592 527876 201644 527882
rect 201592 527818 201644 527824
rect 202144 526448 202196 526454
rect 202144 526390 202196 526396
rect 202156 479602 202184 526390
rect 203522 522336 203578 522345
rect 204456 522306 204484 539158
rect 204640 539158 205022 539186
rect 204640 529242 204668 539158
rect 205560 536110 205588 539172
rect 205744 539158 206310 539186
rect 205548 536104 205600 536110
rect 205548 536046 205600 536052
rect 204902 532128 204958 532137
rect 204902 532063 204958 532072
rect 204628 529236 204680 529242
rect 204628 529178 204680 529184
rect 203522 522271 203578 522280
rect 204444 522300 204496 522306
rect 203536 497486 203564 522271
rect 204444 522242 204496 522248
rect 203524 497480 203576 497486
rect 203524 497422 203576 497428
rect 202234 480856 202290 480865
rect 202234 480791 202290 480800
rect 202144 479596 202196 479602
rect 202144 479538 202196 479544
rect 202248 462233 202276 480791
rect 204166 464536 204222 464545
rect 204166 464471 204222 464480
rect 201590 462224 201646 462233
rect 201590 462159 201646 462168
rect 202234 462224 202290 462233
rect 202234 462159 202290 462168
rect 201500 461508 201552 461514
rect 201500 461450 201552 461456
rect 201512 461038 201540 461450
rect 201500 461032 201552 461038
rect 201604 461009 201632 462159
rect 202326 461544 202382 461553
rect 202144 461508 202196 461514
rect 202326 461479 202382 461488
rect 202144 461450 202196 461456
rect 201500 460974 201552 460980
rect 201590 461000 201646 461009
rect 201590 460935 201646 460944
rect 201406 459096 201462 459105
rect 201406 459031 201462 459040
rect 201420 452985 201448 459031
rect 200854 452976 200910 452985
rect 200854 452911 200910 452920
rect 201406 452976 201462 452985
rect 201406 452911 201462 452920
rect 200212 452668 200264 452674
rect 200212 452610 200264 452616
rect 199476 452600 199528 452606
rect 199476 452542 199528 452548
rect 199382 450392 199438 450401
rect 199382 450327 199438 450336
rect 200224 450242 200252 452610
rect 200868 450242 200896 452911
rect 201604 451274 201632 460935
rect 202156 454034 202184 461450
rect 202144 454028 202196 454034
rect 202144 453970 202196 453976
rect 201604 451246 201816 451274
rect 201788 450242 201816 451246
rect 200224 450214 200422 450242
rect 200868 450214 201342 450242
rect 201788 450214 202262 450242
rect 195242 449984 195298 449993
rect 195242 449919 195298 449928
rect 202340 449750 202368 461479
rect 204180 460934 204208 464471
rect 204088 460906 204208 460934
rect 203154 452704 203210 452713
rect 203154 452639 203210 452648
rect 203168 450228 203196 452639
rect 204088 451353 204116 460906
rect 204536 458652 204588 458658
rect 204536 458594 204588 458600
rect 204548 458318 204576 458594
rect 204536 458312 204588 458318
rect 204536 458254 204588 458260
rect 204074 451344 204130 451353
rect 204074 451279 204130 451288
rect 204088 450228 204116 451279
rect 204548 450242 204576 458254
rect 204916 454753 204944 532063
rect 205640 527944 205692 527950
rect 205640 527886 205692 527892
rect 204994 522472 205050 522481
rect 204994 522407 205050 522416
rect 205008 458833 205036 522407
rect 205088 502988 205140 502994
rect 205088 502930 205140 502936
rect 205100 464409 205128 502930
rect 205086 464400 205142 464409
rect 205086 464335 205142 464344
rect 205548 463004 205600 463010
rect 205548 462946 205600 462952
rect 204994 458824 205050 458833
rect 204994 458759 205050 458768
rect 205560 458658 205588 462946
rect 205548 458652 205600 458658
rect 205548 458594 205600 458600
rect 204902 454744 204958 454753
rect 204902 454679 204958 454688
rect 204548 450214 205022 450242
rect 205652 449970 205680 527886
rect 205744 514146 205772 539158
rect 206282 535528 206338 535537
rect 206282 535463 206338 535472
rect 206376 535492 206428 535498
rect 205732 514140 205784 514146
rect 205732 514082 205784 514088
rect 206296 468489 206324 535463
rect 206376 535434 206428 535440
rect 206388 493338 206416 535434
rect 206848 532710 206876 539172
rect 207400 538257 207428 539172
rect 207386 538248 207442 538257
rect 207386 538183 207442 538192
rect 208136 535537 208164 539172
rect 208412 539158 208702 539186
rect 209056 539158 209438 539186
rect 208122 535528 208178 535537
rect 208122 535463 208178 535472
rect 206836 532704 206888 532710
rect 206836 532646 206888 532652
rect 207664 530596 207716 530602
rect 207664 530538 207716 530544
rect 206376 493332 206428 493338
rect 206376 493274 206428 493280
rect 207676 485081 207704 530538
rect 208412 523734 208440 539158
rect 209056 528554 209084 539158
rect 209976 535498 210004 539172
rect 210344 539158 210726 539186
rect 211172 539158 211278 539186
rect 209964 535492 210016 535498
rect 209964 535434 210016 535440
rect 210344 528554 210372 539158
rect 208504 528526 209084 528554
rect 209884 528526 210372 528554
rect 208504 527134 208532 528526
rect 208492 527128 208544 527134
rect 208492 527070 208544 527076
rect 208400 523728 208452 523734
rect 208400 523670 208452 523676
rect 207662 485072 207718 485081
rect 207662 485007 207718 485016
rect 208504 478174 208532 527070
rect 209884 483682 209912 528526
rect 210424 516860 210476 516866
rect 210424 516802 210476 516808
rect 209872 483676 209924 483682
rect 209872 483618 209924 483624
rect 208492 478168 208544 478174
rect 208492 478110 208544 478116
rect 206282 468480 206338 468489
rect 206282 468415 206338 468424
rect 208398 461680 208454 461689
rect 208398 461615 208454 461624
rect 207020 454028 207072 454034
rect 207020 453970 207072 453976
rect 207032 450228 207060 453970
rect 207940 452736 207992 452742
rect 207940 452678 207992 452684
rect 207952 450228 207980 452678
rect 208412 450242 208440 461615
rect 210436 454102 210464 516802
rect 210608 483676 210660 483682
rect 210608 483618 210660 483624
rect 210514 481672 210570 481681
rect 210514 481607 210570 481616
rect 209780 454096 209832 454102
rect 209780 454038 209832 454044
rect 210424 454096 210476 454102
rect 210424 454038 210476 454044
rect 208412 450214 208886 450242
rect 209792 450228 209820 454038
rect 210528 451926 210556 481607
rect 210620 479602 210648 483618
rect 210608 479596 210660 479602
rect 210608 479538 210660 479544
rect 211172 478242 211200 539158
rect 212000 536722 212028 539172
rect 212566 539158 212672 539186
rect 211988 536716 212040 536722
rect 211988 536658 212040 536664
rect 212000 534478 212028 536658
rect 211988 534472 212040 534478
rect 211988 534414 212040 534420
rect 212540 533384 212592 533390
rect 212540 533326 212592 533332
rect 211802 531992 211858 532001
rect 211802 531927 211858 531936
rect 211160 478236 211212 478242
rect 211160 478178 211212 478184
rect 211816 471345 211844 531927
rect 211802 471336 211858 471345
rect 211802 471271 211858 471280
rect 212552 464370 212580 533326
rect 212644 532137 212672 539158
rect 212724 534472 212776 534478
rect 212724 534414 212776 534420
rect 212630 532128 212686 532137
rect 212630 532063 212686 532072
rect 212736 528554 212764 534414
rect 213104 533497 213132 539172
rect 213472 539158 213854 539186
rect 213932 539158 214406 539186
rect 214576 539158 215142 539186
rect 213090 533488 213146 533497
rect 213090 533423 213146 533432
rect 213472 533390 213500 539158
rect 213460 533384 213512 533390
rect 213460 533326 213512 533332
rect 213184 533248 213236 533254
rect 213184 533190 213236 533196
rect 212644 528526 212764 528554
rect 212644 501770 212672 528526
rect 212632 501764 212684 501770
rect 212632 501706 212684 501712
rect 212644 501634 212672 501706
rect 212632 501628 212684 501634
rect 212632 501570 212684 501576
rect 213196 491978 213224 533190
rect 213276 501764 213328 501770
rect 213276 501706 213328 501712
rect 213184 491972 213236 491978
rect 213184 491914 213236 491920
rect 213288 467945 213316 501706
rect 213932 468586 213960 539158
rect 214576 528554 214604 539158
rect 215680 538214 215708 539172
rect 216416 538286 216444 539172
rect 216784 539158 216982 539186
rect 217336 539158 217718 539186
rect 218164 539158 218270 539186
rect 216404 538280 216456 538286
rect 216404 538222 216456 538228
rect 215312 538186 215708 538214
rect 215312 536790 215340 538186
rect 215300 536784 215352 536790
rect 215300 536726 215352 536732
rect 214024 528526 214604 528554
rect 214024 509930 214052 528526
rect 214012 509924 214064 509930
rect 214012 509866 214064 509872
rect 214654 509824 214710 509833
rect 214654 509759 214710 509768
rect 214564 505844 214616 505850
rect 214564 505786 214616 505792
rect 213920 468580 213972 468586
rect 213920 468522 213972 468528
rect 212630 467936 212686 467945
rect 212630 467871 212686 467880
rect 213274 467936 213330 467945
rect 213274 467871 213330 467880
rect 212540 464364 212592 464370
rect 212540 464306 212592 464312
rect 211160 455456 211212 455462
rect 211160 455398 211212 455404
rect 210516 451920 210568 451926
rect 210516 451862 210568 451868
rect 210528 450242 210556 451862
rect 211172 450242 211200 455398
rect 212644 450242 212672 467871
rect 213828 461644 213880 461650
rect 213828 461586 213880 461592
rect 213840 459678 213868 461586
rect 213276 459672 213328 459678
rect 213276 459614 213328 459620
rect 213828 459672 213880 459678
rect 213828 459614 213880 459620
rect 213288 450242 213316 459614
rect 214576 457570 214604 505786
rect 214668 486577 214696 509759
rect 214654 486568 214710 486577
rect 214654 486503 214710 486512
rect 215312 480962 215340 536726
rect 215944 535492 215996 535498
rect 215944 535434 215996 535440
rect 215956 503062 215984 535434
rect 216036 534744 216088 534750
rect 216036 534686 216088 534692
rect 216048 515438 216076 534686
rect 216680 533384 216732 533390
rect 216680 533326 216732 533332
rect 216036 515432 216088 515438
rect 216036 515374 216088 515380
rect 215944 503056 215996 503062
rect 215944 502998 215996 503004
rect 215944 490680 215996 490686
rect 215944 490622 215996 490628
rect 215300 480956 215352 480962
rect 215300 480898 215352 480904
rect 215300 465724 215352 465730
rect 215300 465666 215352 465672
rect 215312 459678 215340 465666
rect 215482 464400 215538 464409
rect 215482 464335 215538 464344
rect 215300 459672 215352 459678
rect 215300 459614 215352 459620
rect 214564 457564 214616 457570
rect 214564 457506 214616 457512
rect 214564 454028 214616 454034
rect 214564 453970 214616 453976
rect 210528 450214 210726 450242
rect 211172 450214 211646 450242
rect 212644 450214 212750 450242
rect 213288 450214 213670 450242
rect 214576 450228 214604 453970
rect 215496 450228 215524 464335
rect 215956 459785 215984 490622
rect 216692 469849 216720 533326
rect 216784 518226 216812 539158
rect 217336 533390 217364 539158
rect 217414 535528 217470 535537
rect 217414 535463 217470 535472
rect 217324 533384 217376 533390
rect 217324 533326 217376 533332
rect 217428 528554 217456 535463
rect 217336 528526 217456 528554
rect 216772 518220 216824 518226
rect 216772 518162 216824 518168
rect 217336 476785 217364 528526
rect 218164 476882 218192 539158
rect 218992 535498 219020 539172
rect 219544 535537 219572 539172
rect 219728 539158 220110 539186
rect 219530 535528 219586 535537
rect 218980 535492 219032 535498
rect 219530 535463 219586 535472
rect 218980 535434 219032 535440
rect 218794 530768 218850 530777
rect 218794 530703 218850 530712
rect 218704 518220 218756 518226
rect 218704 518162 218756 518168
rect 218716 492046 218744 518162
rect 218704 492040 218756 492046
rect 218704 491982 218756 491988
rect 218152 476876 218204 476882
rect 218152 476818 218204 476824
rect 217322 476776 217378 476785
rect 217322 476711 217378 476720
rect 218808 475425 218836 530703
rect 219728 528554 219756 539158
rect 220084 535560 220136 535566
rect 220084 535502 220136 535508
rect 219452 528526 219756 528554
rect 219452 505782 219480 528526
rect 220096 527785 220124 535502
rect 220082 527776 220138 527785
rect 220082 527711 220138 527720
rect 220084 525156 220136 525162
rect 220084 525098 220136 525104
rect 219440 505776 219492 505782
rect 219440 505718 219492 505724
rect 218794 475416 218850 475425
rect 218794 475351 218850 475360
rect 216772 471368 216824 471374
rect 216772 471310 216824 471316
rect 216678 469840 216734 469849
rect 216678 469775 216734 469784
rect 216784 463729 216812 471310
rect 218702 465896 218758 465905
rect 218702 465831 218758 465840
rect 217416 465112 217468 465118
rect 217416 465054 217468 465060
rect 216770 463720 216826 463729
rect 216770 463655 216826 463664
rect 216784 460934 216812 463655
rect 216784 460906 216904 460934
rect 215942 459776 215998 459785
rect 215942 459711 215998 459720
rect 215956 454034 215984 459711
rect 216036 459672 216088 459678
rect 216036 459614 216088 459620
rect 215944 454028 215996 454034
rect 215944 453970 215996 453976
rect 216048 450242 216076 459614
rect 216876 450242 216904 460906
rect 217428 460222 217456 465054
rect 217416 460216 217468 460222
rect 217416 460158 217468 460164
rect 218716 459921 218744 465831
rect 218058 459912 218114 459921
rect 218058 459847 218114 459856
rect 218702 459912 218758 459921
rect 218702 459847 218758 459856
rect 218072 450242 218100 459847
rect 218888 457496 218940 457502
rect 218888 457438 218940 457444
rect 218900 450242 218928 457438
rect 220096 455462 220124 525098
rect 220832 497486 220860 539172
rect 221384 538354 221412 539172
rect 221372 538348 221424 538354
rect 221372 538290 221424 538296
rect 222120 537441 222148 539172
rect 222304 539158 222686 539186
rect 222106 537432 222162 537441
rect 222106 537367 222162 537376
rect 222304 530602 222332 539158
rect 223408 535566 223436 539172
rect 223396 535560 223448 535566
rect 222934 535528 222990 535537
rect 222844 535492 222896 535498
rect 223396 535502 223448 535508
rect 223960 535498 223988 539172
rect 224696 538286 224724 539172
rect 224684 538280 224736 538286
rect 224684 538222 224736 538228
rect 222934 535463 222990 535472
rect 223948 535492 224000 535498
rect 222844 535434 222896 535440
rect 222292 530596 222344 530602
rect 222292 530538 222344 530544
rect 220820 497480 220872 497486
rect 220820 497422 220872 497428
rect 222108 491972 222160 491978
rect 222108 491914 222160 491920
rect 220084 455456 220136 455462
rect 220084 455398 220136 455404
rect 220096 451274 220124 455398
rect 222120 454209 222148 491914
rect 222856 461553 222884 535434
rect 222948 497457 222976 535463
rect 223948 535434 224000 535440
rect 224696 535401 224724 538222
rect 225248 536042 225276 539172
rect 225524 539158 225998 539186
rect 225236 536036 225288 536042
rect 225236 535978 225288 535984
rect 224682 535392 224738 535401
rect 224682 535327 224738 535336
rect 224696 534177 224724 535327
rect 223670 534168 223726 534177
rect 223670 534103 223726 534112
rect 224682 534168 224738 534177
rect 224682 534103 224738 534112
rect 222934 497448 222990 497457
rect 222934 497383 222990 497392
rect 223488 493332 223540 493338
rect 223488 493274 223540 493280
rect 222842 461544 222898 461553
rect 222842 461479 222898 461488
rect 223500 455122 223528 493274
rect 223580 465724 223632 465730
rect 223580 465666 223632 465672
rect 222568 455116 222620 455122
rect 222568 455058 222620 455064
rect 223488 455116 223540 455122
rect 223488 455058 223540 455064
rect 222106 454200 222162 454209
rect 222106 454135 222162 454144
rect 221188 453212 221240 453218
rect 221188 453154 221240 453160
rect 219820 451246 220124 451274
rect 219820 450242 219848 451246
rect 216048 450214 216430 450242
rect 216876 450214 217350 450242
rect 218072 450214 218454 450242
rect 218900 450214 219374 450242
rect 219820 450214 220294 450242
rect 221200 450228 221228 453154
rect 222120 451274 222148 454135
rect 222580 454102 222608 455058
rect 222568 454096 222620 454102
rect 222568 454038 222620 454044
rect 221660 451246 222148 451274
rect 221660 450242 221688 451246
rect 222580 450242 222608 454038
rect 223592 451274 223620 465666
rect 223684 456929 223712 534103
rect 225524 528554 225552 539158
rect 226536 535537 226564 539172
rect 226720 539158 227102 539186
rect 227732 539158 227838 539186
rect 228008 539158 228390 539186
rect 226522 535528 226578 535537
rect 226522 535463 226578 535472
rect 226248 528624 226300 528630
rect 226248 528566 226300 528572
rect 224972 528526 225552 528554
rect 224972 523705 225000 528526
rect 224958 523696 225014 523705
rect 224958 523631 225014 523640
rect 226156 482996 226208 483002
rect 226156 482938 226208 482944
rect 224958 463720 225014 463729
rect 224958 463655 225014 463664
rect 224972 460934 225000 463655
rect 224972 460906 225644 460934
rect 223670 456920 223726 456929
rect 223670 456855 223726 456864
rect 223684 454073 223712 456855
rect 225052 456816 225104 456822
rect 225052 456758 225104 456764
rect 223670 454064 223726 454073
rect 223670 453999 223726 454008
rect 223684 453218 223712 453999
rect 223672 453212 223724 453218
rect 223672 453154 223724 453160
rect 223592 451246 223712 451274
rect 223684 450242 223712 451246
rect 221660 450214 222134 450242
rect 222580 450214 223054 450242
rect 223684 450214 224158 450242
rect 225064 450228 225092 456758
rect 225616 450242 225644 460906
rect 226168 456822 226196 482938
rect 226260 463729 226288 528566
rect 226720 528554 226748 539158
rect 226984 536036 227036 536042
rect 226984 535978 227036 535984
rect 226352 528526 226748 528554
rect 226352 483002 226380 528526
rect 226996 488238 227024 535978
rect 227732 509833 227760 539158
rect 228008 528554 228036 539158
rect 229112 528630 229140 539172
rect 229664 535498 229692 539172
rect 229652 535492 229704 535498
rect 229652 535434 229704 535440
rect 230400 534750 230428 539172
rect 230492 539158 230966 539186
rect 231228 539158 231702 539186
rect 231964 539158 232254 539186
rect 232424 539158 232806 539186
rect 233344 539158 233542 539186
rect 233712 539158 234094 539186
rect 234724 539158 234830 539186
rect 235000 539158 235382 539186
rect 230388 534744 230440 534750
rect 230388 534686 230440 534692
rect 229742 530632 229798 530641
rect 229742 530567 229798 530576
rect 229100 528624 229152 528630
rect 229100 528566 229152 528572
rect 227824 528526 228036 528554
rect 227824 526454 227852 528526
rect 227812 526448 227864 526454
rect 227812 526390 227864 526396
rect 227718 509824 227774 509833
rect 227718 509759 227774 509768
rect 229756 498846 229784 530567
rect 229836 526448 229888 526454
rect 229836 526390 229888 526396
rect 229848 508570 229876 526390
rect 229836 508564 229888 508570
rect 229836 508506 229888 508512
rect 229744 498840 229796 498846
rect 229744 498782 229796 498788
rect 226984 488232 227036 488238
rect 226984 488174 227036 488180
rect 229100 488232 229152 488238
rect 229100 488174 229152 488180
rect 227076 487892 227128 487898
rect 227076 487834 227128 487840
rect 226340 482996 226392 483002
rect 226340 482938 226392 482944
rect 226432 481704 226484 481710
rect 226432 481646 226484 481652
rect 226246 463720 226302 463729
rect 226246 463655 226302 463664
rect 226156 456816 226208 456822
rect 226156 456758 226208 456764
rect 226444 450242 226472 481646
rect 227088 464370 227116 487834
rect 227812 479596 227864 479602
rect 227812 479538 227864 479544
rect 227718 468072 227774 468081
rect 227718 468007 227774 468016
rect 227732 466546 227760 468007
rect 227720 466540 227772 466546
rect 227720 466482 227772 466488
rect 227076 464364 227128 464370
rect 227076 464306 227128 464312
rect 227732 450242 227760 466482
rect 227824 454034 227852 479538
rect 229112 472122 229140 488174
rect 230492 475425 230520 539158
rect 231228 530602 231256 539158
rect 231860 532772 231912 532778
rect 231860 532714 231912 532720
rect 231216 530596 231268 530602
rect 231216 530538 231268 530544
rect 231122 526416 231178 526425
rect 231122 526351 231178 526360
rect 230478 475416 230534 475425
rect 230478 475351 230534 475360
rect 229100 472116 229152 472122
rect 229100 472058 229152 472064
rect 229112 460934 229140 472058
rect 231136 460934 231164 526351
rect 231872 478145 231900 532714
rect 231964 504422 231992 539158
rect 232424 532778 232452 539158
rect 233240 533384 233292 533390
rect 233240 533326 233292 533332
rect 232412 532772 232464 532778
rect 232412 532714 232464 532720
rect 232502 511320 232558 511329
rect 232502 511255 232558 511264
rect 231952 504416 232004 504422
rect 231952 504358 232004 504364
rect 231858 478136 231914 478145
rect 231858 478071 231914 478080
rect 232516 465633 232544 511255
rect 232596 488572 232648 488578
rect 232596 488514 232648 488520
rect 232502 465624 232558 465633
rect 232502 465559 232558 465568
rect 229112 460906 229232 460934
rect 231136 460906 231256 460934
rect 227812 454028 227864 454034
rect 227812 453970 227864 453976
rect 228732 454028 228784 454034
rect 228732 453970 228784 453976
rect 228744 451625 228772 453970
rect 228730 451616 228786 451625
rect 228730 451551 228786 451560
rect 225616 450214 225998 450242
rect 226444 450214 226918 450242
rect 227732 450214 227838 450242
rect 228744 450228 228772 451551
rect 229204 450242 229232 460906
rect 231228 456929 231256 460906
rect 232134 458824 232190 458833
rect 232134 458759 232190 458768
rect 231214 456920 231270 456929
rect 231214 456855 231270 456864
rect 230756 454028 230808 454034
rect 230756 453970 230808 453976
rect 229204 450214 229678 450242
rect 230768 450228 230796 453970
rect 231228 450242 231256 456855
rect 232148 450242 232176 458759
rect 232608 455569 232636 488514
rect 233252 479602 233280 533326
rect 233344 523734 233372 539158
rect 233424 535832 233476 535838
rect 233424 535774 233476 535780
rect 233436 533458 233464 535774
rect 233424 533452 233476 533458
rect 233424 533394 233476 533400
rect 233712 533390 233740 539158
rect 233884 535492 233936 535498
rect 233884 535434 233936 535440
rect 233700 533384 233752 533390
rect 233700 533326 233752 533332
rect 233332 523728 233384 523734
rect 233332 523670 233384 523676
rect 233240 479596 233292 479602
rect 233240 479538 233292 479544
rect 233238 465624 233294 465633
rect 233238 465559 233294 465568
rect 233252 465225 233280 465559
rect 233238 465216 233294 465225
rect 233238 465151 233294 465160
rect 233148 460216 233200 460222
rect 233148 460158 233200 460164
rect 233160 458833 233188 460158
rect 233146 458824 233202 458833
rect 233146 458759 233202 458768
rect 232594 455560 232650 455569
rect 232594 455495 232650 455504
rect 232608 454034 232636 455495
rect 232596 454028 232648 454034
rect 232596 453970 232648 453976
rect 233252 452849 233280 465151
rect 233238 452840 233294 452849
rect 233238 452775 233294 452784
rect 233252 450242 233280 452775
rect 233896 450673 233924 535434
rect 234620 533384 234672 533390
rect 234620 533326 234672 533332
rect 234632 514078 234660 533326
rect 234724 525162 234752 539158
rect 235000 533390 235028 539158
rect 234988 533384 235040 533390
rect 234988 533326 235040 533332
rect 234712 525156 234764 525162
rect 234712 525098 234764 525104
rect 234620 514072 234672 514078
rect 234620 514014 234672 514020
rect 236104 513330 236132 539172
rect 236656 535838 236684 539172
rect 236644 535832 236696 535838
rect 236644 535774 236696 535780
rect 237392 533390 237420 539172
rect 237484 539158 237958 539186
rect 237380 533384 237432 533390
rect 237380 533326 237432 533332
rect 237484 518226 237512 539158
rect 238680 535430 238708 539172
rect 239232 538218 239260 539172
rect 239324 539158 239798 539186
rect 240244 539158 240534 539186
rect 240704 539158 241086 539186
rect 241532 539158 241822 539186
rect 241900 539158 242374 539186
rect 242912 539158 243110 539186
rect 243188 539158 243662 539186
rect 239220 538212 239272 538218
rect 239220 538154 239272 538160
rect 238208 535424 238260 535430
rect 238208 535366 238260 535372
rect 238668 535424 238720 535430
rect 238668 535366 238720 535372
rect 237564 533384 237616 533390
rect 238220 533361 238248 535366
rect 237564 533326 237616 533332
rect 238206 533352 238262 533361
rect 237472 518220 237524 518226
rect 237472 518162 237524 518168
rect 237576 515438 237604 533326
rect 238206 533287 238262 533296
rect 238024 529236 238076 529242
rect 238024 529178 238076 529184
rect 237564 515432 237616 515438
rect 237564 515374 237616 515380
rect 236092 513324 236144 513330
rect 236092 513266 236144 513272
rect 235906 483848 235962 483857
rect 235906 483783 235962 483792
rect 235920 462233 235948 483783
rect 238036 471889 238064 529178
rect 239324 528554 239352 539158
rect 239404 538212 239456 538218
rect 239404 538154 239456 538160
rect 238772 528526 239352 528554
rect 238772 516798 238800 528526
rect 239416 525094 239444 538154
rect 240140 533384 240192 533390
rect 240140 533326 240192 533332
rect 239404 525088 239456 525094
rect 239404 525030 239456 525036
rect 239402 518936 239458 518945
rect 239402 518871 239458 518880
rect 238760 516792 238812 516798
rect 238760 516734 238812 516740
rect 238116 513324 238168 513330
rect 238116 513266 238168 513272
rect 237378 471880 237434 471889
rect 237378 471815 237434 471824
rect 238022 471880 238078 471889
rect 238022 471815 238078 471824
rect 237392 470665 237420 471815
rect 237378 470656 237434 470665
rect 237378 470591 237434 470600
rect 236000 465112 236052 465118
rect 236000 465054 236052 465060
rect 236012 463593 236040 465054
rect 235998 463584 236054 463593
rect 235998 463519 236054 463528
rect 234618 462224 234674 462233
rect 234618 462159 234674 462168
rect 235906 462224 235962 462233
rect 235906 462159 235962 462168
rect 234632 460934 234660 462159
rect 235920 461009 235948 462159
rect 235906 461000 235962 461009
rect 235906 460935 235962 460944
rect 237392 460934 237420 470591
rect 234632 460906 234936 460934
rect 237392 460906 237972 460934
rect 234436 457564 234488 457570
rect 234436 457506 234488 457512
rect 234448 452674 234476 457506
rect 234436 452668 234488 452674
rect 234436 452610 234488 452616
rect 233882 450664 233938 450673
rect 233882 450599 233938 450608
rect 231228 450214 231702 450242
rect 232148 450214 232622 450242
rect 233252 450214 233542 450242
rect 234448 450228 234476 452610
rect 234908 450242 234936 460906
rect 237470 458280 237526 458289
rect 237470 458215 237526 458224
rect 236460 452736 236512 452742
rect 236460 452678 236512 452684
rect 234908 450214 235382 450242
rect 236472 450228 236500 452678
rect 237484 450242 237512 458215
rect 237406 450214 237512 450242
rect 237944 450242 237972 460906
rect 238128 458289 238156 513266
rect 239416 491366 239444 518871
rect 239404 491360 239456 491366
rect 239404 491302 239456 491308
rect 239494 476232 239550 476241
rect 239494 476167 239550 476176
rect 239402 471200 239458 471209
rect 239402 471135 239458 471144
rect 238114 458280 238170 458289
rect 238114 458215 238170 458224
rect 239416 455938 239444 471135
rect 239508 462913 239536 476167
rect 240152 474026 240180 533326
rect 240244 502994 240272 539158
rect 240704 533390 240732 539158
rect 240692 533384 240744 533390
rect 240692 533326 240744 533332
rect 240232 502988 240284 502994
rect 240232 502930 240284 502936
rect 241428 491360 241480 491366
rect 241428 491302 241480 491308
rect 241440 484430 241468 491302
rect 241428 484424 241480 484430
rect 241428 484366 241480 484372
rect 240782 481536 240838 481545
rect 240782 481471 240838 481480
rect 240796 480282 240824 481471
rect 240784 480276 240836 480282
rect 240784 480218 240836 480224
rect 240140 474020 240192 474026
rect 240140 473962 240192 473968
rect 239494 462904 239550 462913
rect 239494 462839 239550 462848
rect 240796 457473 240824 480218
rect 241428 464432 241480 464438
rect 241428 464374 241480 464380
rect 240782 457464 240838 457473
rect 240782 457399 240838 457408
rect 238760 455932 238812 455938
rect 238760 455874 238812 455880
rect 239404 455932 239456 455938
rect 239404 455874 239456 455880
rect 238772 450242 238800 455874
rect 239416 455530 239444 455874
rect 239404 455524 239456 455530
rect 239404 455466 239456 455472
rect 238850 452840 238906 452849
rect 238850 452775 238906 452784
rect 238864 451217 238892 452775
rect 241440 451382 241468 464374
rect 241532 458862 241560 539158
rect 241900 528554 241928 539158
rect 241624 528526 241928 528554
rect 241624 487830 241652 528526
rect 242912 498846 242940 539158
rect 242992 535492 243044 535498
rect 242992 535434 243044 535440
rect 243004 534070 243032 535434
rect 242992 534064 243044 534070
rect 242992 534006 243044 534012
rect 243188 528601 243216 539158
rect 244384 538150 244412 539172
rect 244372 538144 244424 538150
rect 244372 538086 244424 538092
rect 244384 532098 244412 538086
rect 244936 535537 244964 539172
rect 245028 539158 245502 539186
rect 245672 539158 246238 539186
rect 244922 535528 244978 535537
rect 244922 535463 244978 535472
rect 245028 533338 245056 539158
rect 245106 537432 245162 537441
rect 245106 537367 245162 537376
rect 244476 533310 245056 533338
rect 244372 532092 244424 532098
rect 244372 532034 244424 532040
rect 243174 528592 243230 528601
rect 243174 528527 243230 528536
rect 243544 526516 243596 526522
rect 243544 526458 243596 526464
rect 242900 498840 242952 498846
rect 241702 498808 241758 498817
rect 242900 498782 242952 498788
rect 241702 498743 241758 498752
rect 241612 487824 241664 487830
rect 241612 487766 241664 487772
rect 241716 474842 241744 498743
rect 243556 494018 243584 526458
rect 244278 505744 244334 505753
rect 244278 505679 244334 505688
rect 242900 494012 242952 494018
rect 242900 493954 242952 493960
rect 243544 494012 243596 494018
rect 243544 493954 243596 493960
rect 242912 492726 242940 493954
rect 242900 492720 242952 492726
rect 242900 492662 242952 492668
rect 241704 474836 241756 474842
rect 241704 474778 241756 474784
rect 242164 474836 242216 474842
rect 242164 474778 242216 474784
rect 242176 463593 242204 474778
rect 241610 463584 241666 463593
rect 241610 463519 241666 463528
rect 242162 463584 242218 463593
rect 242162 463519 242218 463528
rect 241624 462369 241652 463519
rect 241610 462360 241666 462369
rect 241610 462295 241666 462304
rect 241624 460934 241652 462295
rect 241624 460906 241744 460934
rect 241520 458856 241572 458862
rect 241520 458798 241572 458804
rect 240140 451376 240192 451382
rect 240140 451318 240192 451324
rect 241428 451376 241480 451382
rect 241428 451318 241480 451324
rect 238850 451208 238906 451217
rect 238850 451143 238906 451152
rect 237944 450214 238326 450242
rect 238772 450214 239246 450242
rect 240152 450228 240180 451318
rect 241060 451308 241112 451314
rect 241060 451250 241112 451256
rect 241072 450228 241100 451250
rect 241716 450242 241744 460906
rect 242912 450242 242940 492662
rect 243544 454708 243596 454714
rect 243544 454650 243596 454656
rect 243556 450242 243584 454650
rect 244292 452742 244320 505679
rect 244476 504490 244504 533310
rect 245120 528554 245148 537367
rect 244936 528526 245148 528554
rect 244936 519586 244964 528526
rect 245672 527950 245700 539158
rect 246776 536761 246804 539172
rect 247144 539158 247526 539186
rect 247696 539158 248078 539186
rect 248524 539158 248814 539186
rect 248984 539158 249366 539186
rect 249904 539158 250102 539186
rect 246762 536752 246818 536761
rect 246762 536687 246818 536696
rect 246302 535528 246358 535537
rect 246302 535463 246358 535472
rect 245660 527944 245712 527950
rect 245660 527886 245712 527892
rect 244924 519580 244976 519586
rect 244924 519522 244976 519528
rect 244464 504484 244516 504490
rect 244464 504426 244516 504432
rect 244370 496632 244426 496641
rect 244370 496567 244426 496576
rect 244384 495514 244412 496567
rect 244372 495508 244424 495514
rect 244372 495450 244424 495456
rect 244384 494766 244412 495450
rect 244372 494760 244424 494766
rect 244372 494702 244424 494708
rect 246316 493406 246344 535463
rect 246396 534744 246448 534750
rect 246396 534686 246448 534692
rect 246408 512650 246436 534686
rect 246948 533452 247000 533458
rect 246948 533394 247000 533400
rect 246396 512644 246448 512650
rect 246396 512586 246448 512592
rect 246304 493400 246356 493406
rect 246304 493342 246356 493348
rect 245568 481704 245620 481710
rect 245568 481646 245620 481652
rect 245580 468586 245608 481646
rect 245568 468580 245620 468586
rect 245568 468522 245620 468528
rect 246960 465730 246988 533394
rect 247040 533384 247092 533390
rect 247040 533326 247092 533332
rect 246948 465724 247000 465730
rect 246948 465666 247000 465672
rect 245660 464364 245712 464370
rect 245660 464306 245712 464312
rect 245672 460934 245700 464306
rect 245672 460906 246344 460934
rect 244922 452840 244978 452849
rect 244922 452775 244978 452784
rect 244280 452736 244332 452742
rect 244280 452678 244332 452684
rect 244292 450537 244320 452678
rect 244278 450528 244334 450537
rect 244278 450463 244334 450472
rect 241716 450214 242190 450242
rect 242912 450214 243110 450242
rect 243556 450214 244030 450242
rect 244936 450228 244964 452775
rect 246316 450242 246344 460906
rect 246316 450214 246790 450242
rect 245750 449984 245806 449993
rect 205652 449954 205942 449970
rect 205640 449948 205942 449954
rect 205692 449942 205942 449948
rect 245806 449942 245870 449970
rect 245750 449919 245806 449928
rect 205640 449890 205692 449896
rect 202328 449744 202380 449750
rect 247052 449721 247080 533326
rect 247144 491978 247172 539158
rect 247696 533390 247724 539158
rect 247684 533384 247736 533390
rect 247684 533326 247736 533332
rect 248524 529242 248552 539158
rect 248512 529236 248564 529242
rect 248512 529178 248564 529184
rect 248984 528554 249012 539158
rect 249064 534812 249116 534818
rect 249064 534754 249116 534760
rect 248432 528526 249012 528554
rect 247132 491972 247184 491978
rect 247132 491914 247184 491920
rect 248432 481710 248460 528526
rect 248512 527876 248564 527882
rect 248512 527818 248564 527824
rect 248420 481704 248472 481710
rect 248420 481646 248472 481652
rect 248524 470594 248552 527818
rect 249076 474065 249104 534754
rect 249904 526425 249932 539158
rect 249890 526416 249946 526425
rect 249890 526351 249946 526360
rect 250456 500274 250484 539242
rect 250640 535498 250668 539172
rect 251192 539158 251390 539186
rect 250628 535492 250680 535498
rect 250628 535434 250680 535440
rect 250444 500268 250496 500274
rect 250444 500210 250496 500216
rect 250444 476876 250496 476882
rect 250444 476818 250496 476824
rect 248602 474056 248658 474065
rect 248602 473991 248658 474000
rect 249062 474056 249118 474065
rect 249062 473991 249118 474000
rect 248432 470566 248552 470594
rect 248432 466478 248460 470566
rect 248420 466472 248472 466478
rect 248420 466414 248472 466420
rect 247408 458244 247460 458250
rect 247408 458186 247460 458192
rect 247420 450242 247448 458186
rect 248432 450242 248460 466414
rect 248616 454034 248644 473991
rect 249064 462392 249116 462398
rect 249064 462334 249116 462340
rect 248604 454028 248656 454034
rect 248604 453970 248656 453976
rect 249076 453966 249104 462334
rect 249708 454028 249760 454034
rect 249708 453970 249760 453976
rect 249064 453960 249116 453966
rect 249064 453902 249116 453908
rect 247420 450214 247894 450242
rect 248432 450214 248814 450242
rect 249614 449984 249670 449993
rect 249720 449970 249748 453970
rect 250456 450294 250484 476818
rect 251086 452568 251142 452577
rect 251086 452503 251142 452512
rect 251100 451926 251128 452503
rect 251088 451920 251140 451926
rect 251088 451862 251140 451868
rect 250626 451480 250682 451489
rect 250626 451415 250682 451424
rect 250640 451314 250668 451415
rect 250628 451308 250680 451314
rect 250628 451250 250680 451256
rect 250444 450288 250496 450294
rect 250444 450230 250496 450236
rect 250640 450228 250668 451250
rect 251192 450498 251220 539158
rect 251468 539073 251496 539310
rect 251454 539064 251510 539073
rect 251454 538999 251510 539008
rect 251928 533390 251956 539172
rect 252020 539158 252494 539186
rect 251916 533384 251968 533390
rect 251916 533326 251968 533332
rect 252020 528554 252048 539158
rect 253216 536110 253244 539172
rect 253204 536104 253256 536110
rect 253204 536046 253256 536052
rect 252466 529136 252522 529145
rect 252466 529071 252522 529080
rect 251284 528526 252048 528554
rect 251284 526454 251312 528526
rect 251272 526448 251324 526454
rect 251272 526390 251324 526396
rect 251272 523728 251324 523734
rect 251272 523670 251324 523676
rect 251284 479534 251312 523670
rect 251824 493400 251876 493406
rect 251824 493342 251876 493348
rect 251272 479528 251324 479534
rect 251272 479470 251324 479476
rect 251284 478922 251312 479470
rect 251272 478916 251324 478922
rect 251272 478858 251324 478864
rect 251548 454028 251600 454034
rect 251548 453970 251600 453976
rect 251560 452985 251588 453970
rect 251546 452976 251602 452985
rect 251546 452911 251602 452920
rect 251180 450492 251232 450498
rect 251180 450434 251232 450440
rect 251560 450228 251588 452911
rect 249670 449956 249748 449970
rect 249670 449942 249734 449956
rect 249614 449919 249670 449928
rect 251836 449750 251864 493342
rect 252480 481681 252508 529071
rect 252560 484424 252612 484430
rect 252558 484392 252560 484401
rect 252612 484392 252614 484401
rect 252558 484327 252614 484336
rect 252466 481672 252522 481681
rect 252466 481607 252522 481616
rect 252480 480865 252508 481607
rect 252466 480856 252522 480865
rect 252466 480791 252522 480800
rect 252560 479596 252612 479602
rect 252560 479538 252612 479544
rect 251916 478916 251968 478922
rect 251916 478858 251968 478864
rect 251928 454034 251956 478858
rect 252572 459610 252600 479538
rect 253308 476241 253336 547846
rect 253386 541104 253442 541113
rect 253386 541039 253442 541048
rect 253400 493338 253428 541039
rect 253952 516866 253980 592243
rect 254030 586936 254086 586945
rect 254030 586871 254086 586880
rect 254044 526522 254072 586871
rect 254136 582321 254164 611322
rect 255320 610020 255372 610026
rect 255320 609962 255372 609968
rect 254676 603220 254728 603226
rect 254676 603162 254728 603168
rect 254582 599584 254638 599593
rect 254582 599519 254638 599528
rect 254596 583030 254624 599519
rect 254688 588606 254716 603162
rect 254766 600672 254822 600681
rect 254766 600607 254822 600616
rect 254780 592657 254808 600607
rect 255332 593042 255360 609962
rect 255976 598913 256004 702510
rect 267660 697610 267688 703520
rect 268384 703112 268436 703118
rect 268384 703054 268436 703060
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 259460 612808 259512 612814
rect 259460 612750 259512 612756
rect 255962 598904 256018 598913
rect 255962 598839 256018 598848
rect 255410 593872 255466 593881
rect 255410 593807 255466 593816
rect 255424 593434 255452 593807
rect 255412 593428 255464 593434
rect 255412 593370 255464 593376
rect 255410 593056 255466 593065
rect 255332 593014 255410 593042
rect 255410 592991 255466 593000
rect 255424 592686 255452 592991
rect 255412 592680 255464 592686
rect 254766 592648 254822 592657
rect 255412 592622 255464 592628
rect 254766 592583 254822 592592
rect 255976 589937 256004 598839
rect 256606 597680 256662 597689
rect 256606 597615 256662 597624
rect 256620 595474 256648 597615
rect 256608 595468 256660 595474
rect 256608 595410 256660 595416
rect 256606 595232 256662 595241
rect 256662 595190 256740 595218
rect 256606 595167 256662 595176
rect 255410 589928 255466 589937
rect 255410 589863 255466 589872
rect 255962 589928 256018 589937
rect 255962 589863 256018 589872
rect 255424 589354 255452 589863
rect 255502 589384 255558 589393
rect 255412 589348 255464 589354
rect 255502 589319 255558 589328
rect 255412 589290 255464 589296
rect 254676 588600 254728 588606
rect 254676 588542 254728 588548
rect 255516 587217 255544 589319
rect 255962 588024 256018 588033
rect 255962 587959 256018 587968
rect 255502 587208 255558 587217
rect 255502 587143 255558 587152
rect 255318 585168 255374 585177
rect 255318 585103 255374 585112
rect 254584 583024 254636 583030
rect 254584 582966 254636 582972
rect 254122 582312 254178 582321
rect 254122 582247 254178 582256
rect 255332 579578 255360 585103
rect 255412 584452 255464 584458
rect 255412 584394 255464 584400
rect 255424 584225 255452 584394
rect 255502 584352 255558 584361
rect 255502 584287 255558 584296
rect 255410 584216 255466 584225
rect 255410 584151 255466 584160
rect 255516 583778 255544 584287
rect 255504 583772 255556 583778
rect 255504 583714 255556 583720
rect 255410 582584 255466 582593
rect 255410 582519 255466 582528
rect 255424 582418 255452 582519
rect 255412 582412 255464 582418
rect 255412 582354 255464 582360
rect 255502 580272 255558 580281
rect 255502 580207 255558 580216
rect 255410 579864 255466 579873
rect 255410 579799 255466 579808
rect 255424 579698 255452 579799
rect 255516 579766 255544 580207
rect 255504 579760 255556 579766
rect 255504 579702 255556 579708
rect 255412 579692 255464 579698
rect 255412 579634 255464 579640
rect 255332 579550 255452 579578
rect 255318 578640 255374 578649
rect 255318 578575 255374 578584
rect 255332 578270 255360 578575
rect 255320 578264 255372 578270
rect 255320 578206 255372 578212
rect 255424 578150 255452 579550
rect 255332 578122 255452 578150
rect 254122 554976 254178 554985
rect 254122 554911 254178 554920
rect 254032 526516 254084 526522
rect 254032 526458 254084 526464
rect 253940 516860 253992 516866
rect 253940 516802 253992 516808
rect 254136 496126 254164 554911
rect 254214 545184 254270 545193
rect 254214 545119 254270 545128
rect 254228 530670 254256 545119
rect 254216 530664 254268 530670
rect 254216 530606 254268 530612
rect 254676 525156 254728 525162
rect 254676 525098 254728 525104
rect 254584 515432 254636 515438
rect 254584 515374 254636 515380
rect 254124 496120 254176 496126
rect 254124 496062 254176 496068
rect 253388 493332 253440 493338
rect 253388 493274 253440 493280
rect 253294 476232 253350 476241
rect 253294 476167 253350 476176
rect 253480 469260 253532 469266
rect 253480 469202 253532 469208
rect 252560 459604 252612 459610
rect 252560 459546 252612 459552
rect 252098 455424 252154 455433
rect 252098 455359 252154 455368
rect 251916 454028 251968 454034
rect 251916 453970 251968 453976
rect 252112 450242 252140 455359
rect 253388 453960 253440 453966
rect 253388 453902 253440 453908
rect 252112 450214 252494 450242
rect 253400 450228 253428 453902
rect 251824 449744 251876 449750
rect 202328 449686 202380 449692
rect 247038 449712 247094 449721
rect 251824 449686 251876 449692
rect 247038 449647 247094 449656
rect 253492 449614 253520 469202
rect 254214 462904 254270 462913
rect 254214 462839 254270 462848
rect 253572 459604 253624 459610
rect 253572 459546 253624 459552
rect 253480 449608 253532 449614
rect 253480 449550 253532 449556
rect 193404 448452 193456 448458
rect 193404 448394 193456 448400
rect 253584 429865 253612 459546
rect 254124 450288 254176 450294
rect 254124 450230 254176 450236
rect 253940 449744 253992 449750
rect 253940 449686 253992 449692
rect 253952 448769 253980 449686
rect 253938 448760 253994 448769
rect 253938 448695 253994 448704
rect 254030 448624 254086 448633
rect 254030 448559 254086 448568
rect 253570 429856 253626 429865
rect 253570 429791 253626 429800
rect 192850 411360 192906 411369
rect 192850 411295 192852 411304
rect 192904 411295 192906 411304
rect 193126 411360 193182 411369
rect 193126 411295 193182 411304
rect 192852 411266 192904 411272
rect 190460 410576 190512 410582
rect 190460 410518 190512 410524
rect 190472 410009 190500 410518
rect 190458 410000 190514 410009
rect 190380 409958 190458 409986
rect 190276 398880 190328 398886
rect 190276 398822 190328 398828
rect 189724 398132 189776 398138
rect 189724 398074 189776 398080
rect 189722 396128 189778 396137
rect 189722 396063 189778 396072
rect 189736 385694 189764 396063
rect 189724 385688 189776 385694
rect 189724 385630 189776 385636
rect 189736 380905 189764 385630
rect 189722 380896 189778 380905
rect 189722 380831 189778 380840
rect 189170 380216 189226 380225
rect 190288 380186 190316 398822
rect 189170 380151 189226 380160
rect 190276 380180 190328 380186
rect 189184 379506 189212 380151
rect 190276 380122 190328 380128
rect 189172 379500 189224 379506
rect 189172 379442 189224 379448
rect 189170 346488 189226 346497
rect 189170 346423 189226 346432
rect 189184 342922 189212 346423
rect 189172 342916 189224 342922
rect 189172 342858 189224 342864
rect 189078 330440 189134 330449
rect 189078 330375 189134 330384
rect 190274 311128 190330 311137
rect 190274 311063 190330 311072
rect 189080 309188 189132 309194
rect 189080 309130 189132 309136
rect 189092 308514 189120 309130
rect 189080 308508 189132 308514
rect 189080 308450 189132 308456
rect 189724 307828 189776 307834
rect 189724 307770 189776 307776
rect 188988 298852 189040 298858
rect 188988 298794 189040 298800
rect 189736 298110 189764 307770
rect 189814 301064 189870 301073
rect 189814 300999 189870 301008
rect 189724 298104 189776 298110
rect 189724 298046 189776 298052
rect 189828 291854 189856 300999
rect 190182 295488 190238 295497
rect 190182 295423 190238 295432
rect 189816 291848 189868 291854
rect 189816 291790 189868 291796
rect 188988 290080 189040 290086
rect 188988 290022 189040 290028
rect 188896 273284 188948 273290
rect 188896 273226 188948 273232
rect 188434 272504 188490 272513
rect 188434 272439 188490 272448
rect 188342 251832 188398 251841
rect 188342 251767 188398 251776
rect 187698 244896 187754 244905
rect 187698 244831 187754 244840
rect 187608 242276 187660 242282
rect 187608 242218 187660 242224
rect 187712 241097 187740 244831
rect 188356 244497 188384 251767
rect 188342 244488 188398 244497
rect 188342 244423 188398 244432
rect 187698 241088 187754 241097
rect 187698 241023 187754 241032
rect 187608 221468 187660 221474
rect 187608 221410 187660 221416
rect 187056 196648 187108 196654
rect 187056 196590 187108 196596
rect 186964 154692 187016 154698
rect 186964 154634 187016 154640
rect 186976 144430 187004 154634
rect 187516 153264 187568 153270
rect 187516 153206 187568 153212
rect 186964 144424 187016 144430
rect 186964 144366 187016 144372
rect 187528 126274 187556 153206
rect 187516 126268 187568 126274
rect 187516 126210 187568 126216
rect 187620 108934 187648 221410
rect 187700 158024 187752 158030
rect 187700 157966 187752 157972
rect 187712 157350 187740 157966
rect 187700 157344 187752 157350
rect 187700 157286 187752 157292
rect 188356 155281 188384 244423
rect 188448 239873 188476 272439
rect 189000 260234 189028 290022
rect 190196 287570 190224 295423
rect 190184 287564 190236 287570
rect 190184 287506 190236 287512
rect 189722 285696 189778 285705
rect 189722 285631 189778 285640
rect 189736 281489 189764 285631
rect 189722 281480 189778 281489
rect 189722 281415 189778 281424
rect 188988 260228 189040 260234
rect 188988 260170 189040 260176
rect 188528 255332 188580 255338
rect 188528 255274 188580 255280
rect 188540 240961 188568 255274
rect 189080 243568 189132 243574
rect 189080 243510 189132 243516
rect 189092 242962 189120 243510
rect 189080 242956 189132 242962
rect 189080 242898 189132 242904
rect 188526 240952 188582 240961
rect 188526 240887 188582 240896
rect 188434 239864 188490 239873
rect 188434 239799 188490 239808
rect 189092 207670 189120 242898
rect 189736 227118 189764 281415
rect 189816 276140 189868 276146
rect 189816 276082 189868 276088
rect 189828 238105 189856 276082
rect 190288 274689 190316 311063
rect 190380 309194 190408 409958
rect 190458 409935 190514 409944
rect 191746 408640 191802 408649
rect 191746 408575 191802 408584
rect 191760 408542 191788 408575
rect 191748 408536 191800 408542
rect 191748 408478 191800 408484
rect 191656 407176 191708 407182
rect 191656 407118 191708 407124
rect 191668 405657 191696 407118
rect 191746 407008 191802 407017
rect 191746 406943 191802 406952
rect 191760 406434 191788 406943
rect 191748 406428 191800 406434
rect 191748 406370 191800 406376
rect 191654 405648 191710 405657
rect 191654 405583 191710 405592
rect 191746 404288 191802 404297
rect 191746 404223 191802 404232
rect 191760 403034 191788 404223
rect 191748 403028 191800 403034
rect 191748 402970 191800 402976
rect 193126 402928 193182 402937
rect 193126 402863 193182 402872
rect 193140 401878 193168 402863
rect 193128 401872 193180 401878
rect 193128 401814 193180 401820
rect 191562 401568 191618 401577
rect 191562 401503 191618 401512
rect 191576 400926 191604 401503
rect 191564 400920 191616 400926
rect 191564 400862 191616 400868
rect 191746 400208 191802 400217
rect 191746 400143 191802 400152
rect 191760 398886 191788 400143
rect 191748 398880 191800 398886
rect 191748 398822 191800 398828
rect 191746 398576 191802 398585
rect 191746 398511 191802 398520
rect 191760 398138 191788 398511
rect 191748 398132 191800 398138
rect 191748 398074 191800 398080
rect 192484 396092 192536 396098
rect 192484 396034 192536 396040
rect 191840 394732 191892 394738
rect 191840 394674 191892 394680
rect 191010 394496 191066 394505
rect 191010 394431 191066 394440
rect 191024 393378 191052 394431
rect 191012 393372 191064 393378
rect 191012 393314 191064 393320
rect 191746 391776 191802 391785
rect 191746 391711 191802 391720
rect 191760 390590 191788 391711
rect 191852 390930 191880 394674
rect 191932 393304 191984 393310
rect 191932 393246 191984 393252
rect 191944 393145 191972 393246
rect 191930 393136 191986 393145
rect 191930 393071 191986 393080
rect 191840 390924 191892 390930
rect 191840 390866 191892 390872
rect 191748 390584 191800 390590
rect 191748 390526 191800 390532
rect 191838 387696 191894 387705
rect 191838 387631 191894 387640
rect 191852 387433 191880 387631
rect 191838 387424 191894 387433
rect 191838 387359 191894 387368
rect 190458 375456 190514 375465
rect 190458 375391 190514 375400
rect 190472 326369 190500 375391
rect 191944 373994 191972 393071
rect 192496 391105 192524 396034
rect 192482 391096 192538 391105
rect 192482 391031 192538 391040
rect 192022 390688 192078 390697
rect 192022 390623 192078 390632
rect 192036 387705 192064 390623
rect 192022 387696 192078 387705
rect 192022 387631 192078 387640
rect 191852 373966 191972 373994
rect 191104 373312 191156 373318
rect 191104 373254 191156 373260
rect 190550 372736 190606 372745
rect 190550 372671 190606 372680
rect 190564 336025 190592 372671
rect 191116 356046 191144 373254
rect 191104 356040 191156 356046
rect 191104 355982 191156 355988
rect 191102 342952 191158 342961
rect 191102 342887 191158 342896
rect 190550 336016 190606 336025
rect 190550 335951 190606 335960
rect 190458 326360 190514 326369
rect 190458 326295 190514 326304
rect 191116 323649 191144 342887
rect 191852 331294 191880 373966
rect 191840 331288 191892 331294
rect 191840 331230 191892 331236
rect 193036 331288 193088 331294
rect 193036 331230 193088 331236
rect 193048 329089 193076 331230
rect 193034 329080 193090 329089
rect 193034 329015 193090 329024
rect 193036 328228 193088 328234
rect 193036 328170 193088 328176
rect 191102 323640 191158 323649
rect 191102 323575 191158 323584
rect 190368 309188 190420 309194
rect 190368 309130 190420 309136
rect 191104 300824 191156 300830
rect 191104 300766 191156 300772
rect 190920 300212 190972 300218
rect 190920 300154 190972 300160
rect 190932 299849 190960 300154
rect 191116 299849 191144 300766
rect 190918 299840 190974 299849
rect 190918 299775 190974 299784
rect 191102 299840 191158 299849
rect 191102 299775 191158 299784
rect 191748 298852 191800 298858
rect 191748 298794 191800 298800
rect 191760 298761 191788 298794
rect 191746 298752 191802 298761
rect 191746 298687 191802 298696
rect 191746 297664 191802 297673
rect 191746 297599 191802 297608
rect 191760 297430 191788 297599
rect 191748 297424 191800 297430
rect 191748 297366 191800 297372
rect 192022 296032 192078 296041
rect 192022 295967 192078 295976
rect 192036 295361 192064 295967
rect 192022 295352 192078 295361
rect 192022 295287 192078 295296
rect 191746 294400 191802 294409
rect 191746 294335 191802 294344
rect 191760 294030 191788 294335
rect 191748 294024 191800 294030
rect 191748 293966 191800 293972
rect 191562 293312 191618 293321
rect 191562 293247 191618 293256
rect 191576 292670 191604 293247
rect 191564 292664 191616 292670
rect 191564 292606 191616 292612
rect 193048 292233 193076 328170
rect 193140 324970 193168 401814
rect 193310 398032 193366 398041
rect 193310 397967 193366 397976
rect 193128 324964 193180 324970
rect 193128 324906 193180 324912
rect 193324 315353 193352 397967
rect 254044 396953 254072 448559
rect 254136 441614 254164 450230
rect 254228 447545 254256 462839
rect 254308 458856 254360 458862
rect 254308 458798 254360 458804
rect 254214 447536 254270 447545
rect 254214 447471 254270 447480
rect 254136 441586 254256 441614
rect 254228 427961 254256 441586
rect 254214 427952 254270 427961
rect 254214 427887 254270 427896
rect 254122 405376 254178 405385
rect 254122 405311 254178 405320
rect 254030 396944 254086 396953
rect 254030 396879 254086 396888
rect 254030 395584 254086 395593
rect 254030 395519 254086 395528
rect 253664 392624 253716 392630
rect 253664 392566 253716 392572
rect 253572 391332 253624 391338
rect 253572 391274 253624 391280
rect 193402 391096 193458 391105
rect 193458 391054 193614 391082
rect 193402 391031 193458 391040
rect 194140 390992 194192 390998
rect 212446 390960 212502 390969
rect 194192 390940 194534 390946
rect 194140 390934 194534 390940
rect 194152 390918 194534 390934
rect 195992 390930 196374 390946
rect 195980 390924 196374 390930
rect 196032 390918 196374 390924
rect 249706 390960 249762 390969
rect 212502 390918 212566 390946
rect 212446 390895 212502 390904
rect 249706 390895 249762 390904
rect 195980 390866 196032 390872
rect 195242 387696 195298 387705
rect 195242 387631 195298 387640
rect 195256 351937 195284 387631
rect 195440 386306 195468 390388
rect 195428 386300 195480 386306
rect 195428 386242 195480 386248
rect 195242 351928 195298 351937
rect 195242 351863 195298 351872
rect 194600 351212 194652 351218
rect 194600 351154 194652 351160
rect 193310 315344 193366 315353
rect 193310 315279 193366 315288
rect 193402 314936 193458 314945
rect 193402 314871 193458 314880
rect 193034 292224 193090 292233
rect 193034 292159 193090 292168
rect 193048 291417 193076 292159
rect 190366 291408 190422 291417
rect 190366 291343 190422 291352
rect 193034 291408 193090 291417
rect 193034 291343 193090 291352
rect 189998 274680 190054 274689
rect 189998 274615 190054 274624
rect 190274 274680 190330 274689
rect 190274 274615 190330 274624
rect 189814 238096 189870 238105
rect 189814 238031 189870 238040
rect 190012 237969 190040 274615
rect 190380 246344 190408 291343
rect 191654 291136 191710 291145
rect 191654 291071 191710 291080
rect 191196 290080 191248 290086
rect 191194 290048 191196 290057
rect 191248 290048 191250 290057
rect 191194 289983 191250 289992
rect 191668 289882 191696 291071
rect 191656 289876 191708 289882
rect 191656 289818 191708 289824
rect 191748 289808 191800 289814
rect 191748 289750 191800 289756
rect 191760 288969 191788 289750
rect 191746 288960 191802 288969
rect 191746 288895 191802 288904
rect 191748 287020 191800 287026
rect 191748 286962 191800 286968
rect 191760 286793 191788 286962
rect 191746 286784 191802 286793
rect 191746 286719 191802 286728
rect 191746 284608 191802 284617
rect 191746 284543 191802 284552
rect 191760 284374 191788 284543
rect 191748 284368 191800 284374
rect 191748 284310 191800 284316
rect 191746 283520 191802 283529
rect 191746 283455 191802 283464
rect 191760 282946 191788 283455
rect 191748 282940 191800 282946
rect 191748 282882 191800 282888
rect 191746 282432 191802 282441
rect 191746 282367 191802 282376
rect 191760 281586 191788 282367
rect 192024 281648 192076 281654
rect 192024 281590 192076 281596
rect 191748 281580 191800 281586
rect 191748 281522 191800 281528
rect 191746 281344 191802 281353
rect 191746 281279 191802 281288
rect 191760 280838 191788 281279
rect 191748 280832 191800 280838
rect 191748 280774 191800 280780
rect 192036 280265 192064 281590
rect 192022 280256 192078 280265
rect 192022 280191 192078 280200
rect 191746 279168 191802 279177
rect 191746 279103 191802 279112
rect 191760 278798 191788 279103
rect 191748 278792 191800 278798
rect 191748 278734 191800 278740
rect 191562 278080 191618 278089
rect 191562 278015 191618 278024
rect 191576 277438 191604 278015
rect 191564 277432 191616 277438
rect 191564 277374 191616 277380
rect 191746 276992 191802 277001
rect 191746 276927 191802 276936
rect 191760 276078 191788 276927
rect 191748 276072 191800 276078
rect 191748 276014 191800 276020
rect 191746 275904 191802 275913
rect 191746 275839 191802 275848
rect 191760 274689 191788 275839
rect 191746 274680 191802 274689
rect 191746 274615 191802 274624
rect 191746 273728 191802 273737
rect 191746 273663 191802 273672
rect 191760 273290 191788 273663
rect 191748 273284 191800 273290
rect 191748 273226 191800 273232
rect 191286 272640 191342 272649
rect 191286 272575 191342 272584
rect 191300 271930 191328 272575
rect 191288 271924 191340 271930
rect 191288 271866 191340 271872
rect 191746 271552 191802 271561
rect 191746 271487 191802 271496
rect 191760 270706 191788 271487
rect 191748 270700 191800 270706
rect 191748 270642 191800 270648
rect 191196 270496 191248 270502
rect 191194 270464 191196 270473
rect 191248 270464 191250 270473
rect 191194 270399 191250 270408
rect 193416 269385 193444 314871
rect 194414 305688 194470 305697
rect 193864 305652 193916 305658
rect 194414 305623 194470 305632
rect 193864 305594 193916 305600
rect 193588 305108 193640 305114
rect 193588 305050 193640 305056
rect 193600 300150 193628 305050
rect 193876 301580 193904 305594
rect 194428 301580 194456 305623
rect 194612 303793 194640 351154
rect 195256 349761 195284 351863
rect 195242 349752 195298 349761
rect 195242 349687 195298 349696
rect 195992 328234 196020 390866
rect 196544 390374 197294 390402
rect 196544 373994 196572 390374
rect 198200 387705 198228 390388
rect 197358 387696 197414 387705
rect 197358 387631 197414 387640
rect 198186 387696 198242 387705
rect 198186 387631 198242 387640
rect 197372 387433 197400 387631
rect 197358 387424 197414 387433
rect 197358 387359 197414 387368
rect 197360 386300 197412 386306
rect 197360 386242 197412 386248
rect 196084 373966 196572 373994
rect 196084 365634 196112 373966
rect 196072 365628 196124 365634
rect 196072 365570 196124 365576
rect 196084 365226 196112 365570
rect 196072 365220 196124 365226
rect 196072 365162 196124 365168
rect 196624 365220 196676 365226
rect 196624 365162 196676 365168
rect 196636 356794 196664 365162
rect 197372 360194 197400 386242
rect 199120 384441 199148 390388
rect 200224 389230 200252 390388
rect 200212 389224 200264 389230
rect 200212 389166 200264 389172
rect 201144 386073 201172 390388
rect 201604 390374 202078 390402
rect 201604 389230 201632 390374
rect 201592 389224 201644 389230
rect 201592 389166 201644 389172
rect 201130 386064 201186 386073
rect 201130 385999 201186 386008
rect 199106 384432 199162 384441
rect 199106 384367 199162 384376
rect 201604 373994 201632 389166
rect 202984 389094 203012 390388
rect 203536 390374 203918 390402
rect 202972 389088 203024 389094
rect 202972 389030 203024 389036
rect 203536 386073 203564 390374
rect 204350 389872 204406 389881
rect 204350 389807 204406 389816
rect 203522 386064 203578 386073
rect 203522 385999 203578 386008
rect 201512 373966 201632 373994
rect 201512 367062 201540 373966
rect 203536 373318 203564 385999
rect 203524 373312 203576 373318
rect 203524 373254 203576 373260
rect 201500 367056 201552 367062
rect 201500 366998 201552 367004
rect 199382 366344 199438 366353
rect 199382 366279 199438 366288
rect 197360 360188 197412 360194
rect 197360 360130 197412 360136
rect 196624 356788 196676 356794
rect 196624 356730 196676 356736
rect 198740 353320 198792 353326
rect 198740 353262 198792 353268
rect 197360 344344 197412 344350
rect 197360 344286 197412 344292
rect 198004 344344 198056 344350
rect 198004 344286 198056 344292
rect 196622 340096 196678 340105
rect 196622 340031 196678 340040
rect 195980 328228 196032 328234
rect 195980 328170 196032 328176
rect 196636 310729 196664 340031
rect 196714 319424 196770 319433
rect 196714 319359 196770 319368
rect 196622 310720 196678 310729
rect 196622 310655 196678 310664
rect 195058 309088 195114 309097
rect 195058 309023 195114 309032
rect 195072 307873 195100 309023
rect 195058 307864 195114 307873
rect 195058 307799 195114 307808
rect 194598 303784 194654 303793
rect 194598 303719 194654 303728
rect 195072 301580 195100 307799
rect 196256 307760 196308 307766
rect 196256 307702 196308 307708
rect 196268 307086 196296 307702
rect 196256 307080 196308 307086
rect 196256 307022 196308 307028
rect 195610 303784 195666 303793
rect 195610 303719 195666 303728
rect 195624 301580 195652 303719
rect 196268 301580 196296 307022
rect 196636 301594 196664 310655
rect 196728 307766 196756 319359
rect 196716 307760 196768 307766
rect 196716 307702 196768 307708
rect 197372 306374 197400 344286
rect 197450 331256 197506 331265
rect 197450 331191 197506 331200
rect 197464 327049 197492 331191
rect 197450 327040 197506 327049
rect 197450 326975 197506 326984
rect 198016 312497 198044 344286
rect 198752 325694 198780 353262
rect 198752 325666 199332 325694
rect 198002 312488 198058 312497
rect 198002 312423 198058 312432
rect 197372 306346 198320 306374
rect 197452 305040 197504 305046
rect 197452 304982 197504 304988
rect 196636 301566 196834 301594
rect 197464 301580 197492 304982
rect 198292 301594 198320 306346
rect 199198 306368 199254 306377
rect 199198 306303 199254 306312
rect 198292 301566 198674 301594
rect 193680 300960 193732 300966
rect 193680 300902 193732 300908
rect 197636 300960 197688 300966
rect 199014 300928 199070 300937
rect 197688 300908 198030 300914
rect 197636 300902 198030 300908
rect 193588 300144 193640 300150
rect 193588 300086 193640 300092
rect 193692 299441 193720 300902
rect 197648 300886 198030 300902
rect 199212 300914 199240 306303
rect 199304 303362 199332 325666
rect 199396 306377 199424 366279
rect 202142 363624 202198 363633
rect 202142 363559 202198 363568
rect 200762 359408 200818 359417
rect 200762 359343 200818 359352
rect 200776 334121 200804 359343
rect 201682 349888 201738 349897
rect 201682 349823 201738 349832
rect 201498 338736 201554 338745
rect 201498 338671 201554 338680
rect 200118 334112 200174 334121
rect 200118 334047 200174 334056
rect 200762 334112 200818 334121
rect 200762 334047 200818 334056
rect 199382 306368 199438 306377
rect 199382 306303 199438 306312
rect 199304 303334 199516 303362
rect 199488 301594 199516 303334
rect 200132 301594 200160 334047
rect 200212 332716 200264 332722
rect 200212 332658 200264 332664
rect 200224 325694 200252 332658
rect 200224 325666 200712 325694
rect 200684 301594 200712 325666
rect 201512 303498 201540 338671
rect 201590 331800 201646 331809
rect 201590 331735 201646 331744
rect 201604 303618 201632 331735
rect 201696 303657 201724 349823
rect 202156 343097 202184 363559
rect 202142 343088 202198 343097
rect 202142 343023 202198 343032
rect 204364 335354 204392 389807
rect 204824 389201 204852 390388
rect 204810 389192 204866 389201
rect 205928 389162 205956 390388
rect 206204 390374 206862 390402
rect 207032 390374 207782 390402
rect 208412 390374 208702 390402
rect 204810 389127 204866 389136
rect 205916 389156 205968 389162
rect 204824 386345 204852 389127
rect 205916 389098 205968 389104
rect 204810 386336 204866 386345
rect 204810 386271 204866 386280
rect 206204 383654 206232 390374
rect 206204 383626 206508 383654
rect 206480 378865 206508 383626
rect 206466 378856 206522 378865
rect 206466 378791 206522 378800
rect 206284 359508 206336 359514
rect 206284 359450 206336 359456
rect 204902 347032 204958 347041
rect 204902 346967 204958 346976
rect 204180 335326 204392 335354
rect 202878 334792 202934 334801
rect 202878 334727 202934 334736
rect 201682 303648 201738 303657
rect 201592 303612 201644 303618
rect 201682 303583 201738 303592
rect 202786 303648 202842 303657
rect 202892 303618 202920 334727
rect 204180 334665 204208 335326
rect 204166 334656 204222 334665
rect 204166 334591 204222 334600
rect 204180 330546 204208 334591
rect 204168 330540 204220 330546
rect 204168 330482 204220 330488
rect 204260 323672 204312 323678
rect 204260 323614 204312 323620
rect 203062 322280 203118 322289
rect 203062 322215 203118 322224
rect 202786 303583 202842 303592
rect 202880 303612 202932 303618
rect 201592 303554 201644 303560
rect 201512 303470 201816 303498
rect 201592 303408 201644 303414
rect 201592 303350 201644 303356
rect 199488 301566 199870 301594
rect 200132 301566 200422 301594
rect 200684 301566 201066 301594
rect 201604 301580 201632 303350
rect 201788 301594 201816 303470
rect 201788 301566 202262 301594
rect 202800 301580 202828 303583
rect 202880 303554 202932 303560
rect 203076 301594 203104 322215
rect 204272 303618 204300 323614
rect 204350 317656 204406 317665
rect 204350 317591 204406 317600
rect 203708 303612 203760 303618
rect 203708 303554 203760 303560
rect 204260 303612 204312 303618
rect 204260 303554 204312 303560
rect 203720 301594 203748 303554
rect 204364 301594 204392 317591
rect 204916 314129 204944 346967
rect 205638 338056 205694 338065
rect 205638 337991 205694 338000
rect 205652 336841 205680 337991
rect 205638 336832 205694 336841
rect 205638 336767 205694 336776
rect 205652 325694 205680 336767
rect 205732 329928 205784 329934
rect 205732 329870 205784 329876
rect 205744 329118 205772 329870
rect 205732 329112 205784 329118
rect 205732 329054 205784 329060
rect 205652 325666 206048 325694
rect 204902 314120 204958 314129
rect 204902 314055 204958 314064
rect 205822 305144 205878 305153
rect 205822 305079 205878 305088
rect 204812 303612 204864 303618
rect 204812 303554 204864 303560
rect 204824 301594 204852 303554
rect 203076 301566 203458 301594
rect 203720 301566 204010 301594
rect 204364 301566 204654 301594
rect 204824 301566 205206 301594
rect 205836 301580 205864 305079
rect 206020 301594 206048 325666
rect 206296 305153 206324 359450
rect 206376 348492 206428 348498
rect 206376 348434 206428 348440
rect 206388 305658 206416 348434
rect 206480 342922 206508 378791
rect 207032 364342 207060 390374
rect 208412 375193 208440 390374
rect 209608 385665 209636 390388
rect 209792 390374 210542 390402
rect 209594 385656 209650 385665
rect 209594 385591 209650 385600
rect 208398 375184 208454 375193
rect 208398 375119 208454 375128
rect 207020 364336 207072 364342
rect 207020 364278 207072 364284
rect 209042 362264 209098 362273
rect 209042 362199 209098 362208
rect 206558 352608 206614 352617
rect 206558 352543 206614 352552
rect 206468 342916 206520 342922
rect 206468 342858 206520 342864
rect 206572 338065 206600 352543
rect 207664 349852 207716 349858
rect 207664 349794 207716 349800
rect 207676 340241 207704 349794
rect 207662 340232 207718 340241
rect 207662 340167 207718 340176
rect 207202 338872 207258 338881
rect 207202 338807 207258 338816
rect 206558 338056 206614 338065
rect 206558 337991 206614 338000
rect 207110 331936 207166 331945
rect 207110 331871 207166 331880
rect 206376 305652 206428 305658
rect 206376 305594 206428 305600
rect 206282 305144 206338 305153
rect 206282 305079 206338 305088
rect 207124 301594 207152 331871
rect 207216 325694 207244 338807
rect 207216 325666 207888 325694
rect 207572 308440 207624 308446
rect 207572 308382 207624 308388
rect 206020 301566 206402 301594
rect 207046 301566 207152 301594
rect 207584 301580 207612 308382
rect 207860 301594 207888 325666
rect 208398 313304 208454 313313
rect 208398 313239 208454 313248
rect 208412 301594 208440 313239
rect 209056 306649 209084 362199
rect 209792 349761 209820 390374
rect 211632 387734 211660 390388
rect 211620 387728 211672 387734
rect 211620 387670 211672 387676
rect 211632 383654 211660 387670
rect 213472 387569 213500 390388
rect 213932 390374 214406 390402
rect 213458 387560 213514 387569
rect 213458 387495 213514 387504
rect 211632 383626 211844 383654
rect 209778 349752 209834 349761
rect 209778 349687 209834 349696
rect 209136 348492 209188 348498
rect 209136 348434 209188 348440
rect 209148 311137 209176 348434
rect 210424 333260 210476 333266
rect 210424 333202 210476 333208
rect 209780 323604 209832 323610
rect 209780 323546 209832 323552
rect 209318 313984 209374 313993
rect 209318 313919 209374 313928
rect 209332 313313 209360 313919
rect 209318 313304 209374 313313
rect 209318 313239 209374 313248
rect 209134 311128 209190 311137
rect 209134 311063 209190 311072
rect 209042 306640 209098 306649
rect 209042 306575 209098 306584
rect 209056 301594 209084 306575
rect 209792 301594 209820 323546
rect 210436 309369 210464 333202
rect 211342 328672 211398 328681
rect 211342 328607 211398 328616
rect 210238 309360 210294 309369
rect 210238 309295 210294 309304
rect 210422 309360 210478 309369
rect 210422 309295 210478 309304
rect 210252 301594 210280 309295
rect 211066 303648 211122 303657
rect 211066 303583 211122 303592
rect 207860 301566 208242 301594
rect 208412 301566 208886 301594
rect 209056 301566 209438 301594
rect 209792 301566 210082 301594
rect 210252 301566 210634 301594
rect 211080 301034 211108 303583
rect 211356 301594 211384 328607
rect 211434 326360 211490 326369
rect 211434 326295 211490 326304
rect 211278 301566 211384 301594
rect 211448 301594 211476 326295
rect 211816 323678 211844 383626
rect 213932 369782 213960 390374
rect 215312 389298 215340 390388
rect 215404 390374 216246 390402
rect 216692 390374 217350 390402
rect 215300 389292 215352 389298
rect 215300 389234 215352 389240
rect 214564 381608 214616 381614
rect 214564 381550 214616 381556
rect 213920 369776 213972 369782
rect 213920 369718 213972 369724
rect 214576 355978 214604 381550
rect 214654 369064 214710 369073
rect 214654 368999 214710 369008
rect 214668 356726 214696 368999
rect 214656 356720 214708 356726
rect 214656 356662 214708 356668
rect 214564 355972 214616 355978
rect 214564 355914 214616 355920
rect 213184 355428 213236 355434
rect 213184 355370 213236 355376
rect 211894 348392 211950 348401
rect 211894 348327 211950 348336
rect 211908 328681 211936 348327
rect 212632 336796 212684 336802
rect 212632 336738 212684 336744
rect 211894 328672 211950 328681
rect 211894 328607 211950 328616
rect 211804 323672 211856 323678
rect 211804 323614 211856 323620
rect 212446 309768 212502 309777
rect 212446 309703 212502 309712
rect 212460 302569 212488 309703
rect 212446 302560 212502 302569
rect 212446 302495 212502 302504
rect 211448 301566 211830 301594
rect 212460 301580 212488 302495
rect 212644 301594 212672 336738
rect 213196 303686 213224 355370
rect 214564 355360 214616 355366
rect 214564 355302 214616 355308
rect 213828 354000 213880 354006
rect 213828 353942 213880 353948
rect 213840 325694 213868 353942
rect 214576 346526 214604 355302
rect 214564 346520 214616 346526
rect 214564 346462 214616 346468
rect 213840 325666 213960 325694
rect 213932 325009 213960 325666
rect 213918 325000 213974 325009
rect 213918 324935 213974 324944
rect 213184 303680 213236 303686
rect 213184 303622 213236 303628
rect 213196 301594 213224 303622
rect 213932 301594 213960 324935
rect 214576 303686 214604 346462
rect 215312 325038 215340 389234
rect 215404 381993 215432 390374
rect 216692 383489 216720 390374
rect 218256 386306 218284 390388
rect 218716 390374 219190 390402
rect 218716 387802 218744 390374
rect 218704 387796 218756 387802
rect 218704 387738 218756 387744
rect 217324 386300 217376 386306
rect 217324 386242 217376 386248
rect 218244 386300 218296 386306
rect 218244 386242 218296 386248
rect 216678 383480 216734 383489
rect 216678 383415 216734 383424
rect 215390 381984 215446 381993
rect 215390 381919 215446 381928
rect 215404 381041 215432 381919
rect 215390 381032 215446 381041
rect 215390 380967 215446 380976
rect 215942 381032 215998 381041
rect 215942 380967 215998 380976
rect 215956 340202 215984 380967
rect 216680 362228 216732 362234
rect 216680 362170 216732 362176
rect 216692 360097 216720 362170
rect 216678 360088 216734 360097
rect 216678 360023 216734 360032
rect 217336 353258 217364 386242
rect 217414 360088 217470 360097
rect 217414 360023 217470 360032
rect 217324 353252 217376 353258
rect 217324 353194 217376 353200
rect 216588 351212 216640 351218
rect 216588 351154 216640 351160
rect 215944 340196 215996 340202
rect 215944 340138 215996 340144
rect 215482 336016 215538 336025
rect 215482 335951 215538 335960
rect 215496 325694 215524 335951
rect 215496 325666 216168 325694
rect 215300 325032 215352 325038
rect 215300 324974 215352 324980
rect 215392 305652 215444 305658
rect 215392 305594 215444 305600
rect 214838 304192 214894 304201
rect 214838 304127 214894 304136
rect 214564 303680 214616 303686
rect 214564 303622 214616 303628
rect 212644 301566 213026 301594
rect 213196 301566 213670 301594
rect 213932 301566 214222 301594
rect 214852 301580 214880 304127
rect 215404 301580 215432 305594
rect 216140 301594 216168 325666
rect 216600 303414 216628 351154
rect 217336 337414 217364 353194
rect 217428 345166 217456 360023
rect 217416 345160 217468 345166
rect 217416 345102 217468 345108
rect 217428 345014 217456 345102
rect 217428 344986 217640 345014
rect 217324 337408 217376 337414
rect 217324 337350 217376 337356
rect 217414 336016 217470 336025
rect 217414 335951 217470 335960
rect 217428 311914 217456 335951
rect 217612 325694 217640 344986
rect 217612 325666 217916 325694
rect 217416 311908 217468 311914
rect 217416 311850 217468 311856
rect 217232 303680 217284 303686
rect 217232 303622 217284 303628
rect 216588 303408 216640 303414
rect 216588 303350 216640 303356
rect 216600 302938 216628 303350
rect 216588 302932 216640 302938
rect 216588 302874 216640 302880
rect 216862 301608 216918 301617
rect 216140 301566 216614 301594
rect 217244 301580 217272 303622
rect 217428 301594 217456 311850
rect 217428 301566 217810 301594
rect 216862 301543 216918 301552
rect 215668 301096 215720 301102
rect 215720 301044 216062 301050
rect 215668 301038 216062 301044
rect 211068 301028 211120 301034
rect 215680 301022 216062 301038
rect 211068 300970 211120 300976
rect 216876 300966 216904 301543
rect 199070 300900 199240 300914
rect 216864 300960 216916 300966
rect 217888 300937 217916 325666
rect 218716 311817 218744 387738
rect 219992 387320 220044 387326
rect 219992 387262 220044 387268
rect 220004 383654 220032 387262
rect 220096 384305 220124 390388
rect 220924 390374 221030 390402
rect 220176 387864 220228 387870
rect 220176 387806 220228 387812
rect 220082 384296 220138 384305
rect 220082 384231 220138 384240
rect 220004 383626 220124 383654
rect 220096 350538 220124 383626
rect 220188 382129 220216 387806
rect 220174 382120 220230 382129
rect 220174 382055 220230 382064
rect 220084 350532 220136 350538
rect 220084 350474 220136 350480
rect 220188 349897 220216 382055
rect 220924 380361 220952 390374
rect 221936 387870 221964 390388
rect 222212 390374 222870 390402
rect 223592 390374 223974 390402
rect 221924 387864 221976 387870
rect 221924 387806 221976 387812
rect 220910 380352 220966 380361
rect 220910 380287 220966 380296
rect 220266 373416 220322 373425
rect 220266 373351 220322 373360
rect 220174 349888 220230 349897
rect 220174 349823 220230 349832
rect 220280 345681 220308 373351
rect 222212 372502 222240 390374
rect 223592 378146 223620 390374
rect 224880 384849 224908 390388
rect 225800 387802 225828 390388
rect 226352 390374 226734 390402
rect 225788 387796 225840 387802
rect 225788 387738 225840 387744
rect 225800 387326 225828 387738
rect 225788 387320 225840 387326
rect 225788 387262 225840 387268
rect 224866 384840 224922 384849
rect 224866 384775 224922 384784
rect 223580 378140 223632 378146
rect 223580 378082 223632 378088
rect 224224 378140 224276 378146
rect 224224 378082 224276 378088
rect 222200 372496 222252 372502
rect 222200 372438 222252 372444
rect 222212 371278 222240 372438
rect 222200 371272 222252 371278
rect 222200 371214 222252 371220
rect 222844 371272 222896 371278
rect 222844 371214 222896 371220
rect 221462 370560 221518 370569
rect 221462 370495 221518 370504
rect 220266 345672 220322 345681
rect 220266 345607 220322 345616
rect 220084 339516 220136 339522
rect 220084 339458 220136 339464
rect 219438 338192 219494 338201
rect 219438 338127 219494 338136
rect 219348 331968 219400 331974
rect 219348 331910 219400 331916
rect 218702 311808 218758 311817
rect 218702 311743 218758 311752
rect 218060 311160 218112 311166
rect 218060 311102 218112 311108
rect 218072 307057 218100 311102
rect 218704 309188 218756 309194
rect 218704 309130 218756 309136
rect 218058 307048 218114 307057
rect 218058 306983 218114 306992
rect 218716 305697 218744 309130
rect 218702 305688 218758 305697
rect 218702 305623 218758 305632
rect 219360 304366 219388 331910
rect 218428 304360 218480 304366
rect 218428 304302 218480 304308
rect 219348 304360 219400 304366
rect 219348 304302 219400 304308
rect 218150 301200 218206 301209
rect 218440 301186 218468 304302
rect 218980 303408 219032 303414
rect 218980 303350 219032 303356
rect 218992 301580 219020 303350
rect 219452 301594 219480 338127
rect 220096 323610 220124 339458
rect 220818 336696 220874 336705
rect 220818 336631 220874 336640
rect 220832 335481 220860 336631
rect 220818 335472 220874 335481
rect 220818 335407 220874 335416
rect 220084 323604 220136 323610
rect 220084 323546 220136 323552
rect 220174 308000 220230 308009
rect 220174 307935 220230 307944
rect 219452 301566 219650 301594
rect 220188 301580 220216 307935
rect 220832 301580 220860 335407
rect 220910 327720 220966 327729
rect 220910 327655 220966 327664
rect 220924 303686 220952 327655
rect 221476 325694 221504 370495
rect 221554 348528 221610 348537
rect 221554 348463 221610 348472
rect 221568 336705 221596 348463
rect 221554 336696 221610 336705
rect 221554 336631 221610 336640
rect 222290 330440 222346 330449
rect 222290 330375 222346 330384
rect 221016 325666 221504 325694
rect 221016 324465 221044 325666
rect 221002 324456 221058 324465
rect 221002 324391 221058 324400
rect 220912 303680 220964 303686
rect 220912 303622 220964 303628
rect 221016 301594 221044 324391
rect 221740 303680 221792 303686
rect 221740 303622 221792 303628
rect 221752 301594 221780 303622
rect 222304 301594 222332 330375
rect 222856 311137 222884 371214
rect 224236 360913 224264 378082
rect 224222 360904 224278 360913
rect 224222 360839 224278 360848
rect 224314 351112 224370 351121
rect 224314 351047 224370 351056
rect 224222 338736 224278 338745
rect 224222 338671 224278 338680
rect 223578 338056 223634 338065
rect 223578 337991 223634 338000
rect 223592 337385 223620 337991
rect 223578 337376 223634 337385
rect 223578 337311 223634 337320
rect 223486 312488 223542 312497
rect 223486 312423 223542 312432
rect 222842 311128 222898 311137
rect 222842 311063 222898 311072
rect 223394 306776 223450 306785
rect 223394 306711 223450 306720
rect 223408 304978 223436 306711
rect 223396 304972 223448 304978
rect 223396 304914 223448 304920
rect 223500 302297 223528 312423
rect 223592 303686 223620 337311
rect 224236 320113 224264 338671
rect 224328 338065 224356 351047
rect 224314 338056 224370 338065
rect 224314 337991 224370 338000
rect 223670 320104 223726 320113
rect 223670 320039 223726 320048
rect 224222 320104 224278 320113
rect 224222 320039 224278 320048
rect 223684 318889 223712 320039
rect 223670 318880 223726 318889
rect 223670 318815 223726 318824
rect 223580 303680 223632 303686
rect 223580 303622 223632 303628
rect 223486 302288 223542 302297
rect 223486 302223 223542 302232
rect 223500 301594 223528 302223
rect 221016 301566 221398 301594
rect 221752 301566 222042 301594
rect 222304 301566 222594 301594
rect 223238 301566 223528 301594
rect 223684 301594 223712 318815
rect 224880 308446 224908 384775
rect 226352 364274 226380 390374
rect 227640 387870 227668 390388
rect 227732 390374 228574 390402
rect 229112 390374 229678 390402
rect 227628 387864 227680 387870
rect 227628 387806 227680 387812
rect 227732 372570 227760 390374
rect 228364 387864 228416 387870
rect 228364 387806 228416 387812
rect 228376 383722 228404 387806
rect 228364 383716 228416 383722
rect 228364 383658 228416 383664
rect 228376 377466 228404 383658
rect 229112 382226 229140 390374
rect 230584 389337 230612 390388
rect 230570 389328 230626 389337
rect 230492 389286 230570 389314
rect 229100 382220 229152 382226
rect 229100 382162 229152 382168
rect 228364 377460 228416 377466
rect 228364 377402 228416 377408
rect 229742 376000 229798 376009
rect 229742 375935 229798 375944
rect 227720 372564 227772 372570
rect 227720 372506 227772 372512
rect 227626 371920 227682 371929
rect 227626 371855 227682 371864
rect 226340 364268 226392 364274
rect 226340 364210 226392 364216
rect 226352 363662 226380 364210
rect 226340 363656 226392 363662
rect 226340 363598 226392 363604
rect 226246 346488 226302 346497
rect 226246 346423 226302 346432
rect 225142 327856 225198 327865
rect 225142 327791 225198 327800
rect 224868 308440 224920 308446
rect 224868 308382 224920 308388
rect 224132 303680 224184 303686
rect 224132 303622 224184 303628
rect 225052 303680 225104 303686
rect 225052 303622 225104 303628
rect 224144 301594 224172 303622
rect 223684 301566 223882 301594
rect 224144 301566 224434 301594
rect 225064 301580 225092 303622
rect 225156 301594 225184 327791
rect 225972 307828 226024 307834
rect 225972 307770 226024 307776
rect 225984 301594 226012 307770
rect 226260 303686 226288 346423
rect 226338 334656 226394 334665
rect 226338 334591 226394 334600
rect 226352 306374 226380 334591
rect 226982 320784 227038 320793
rect 226982 320719 227038 320728
rect 226352 306346 226472 306374
rect 226248 303680 226300 303686
rect 226248 303622 226300 303628
rect 226444 301594 226472 306346
rect 226996 301594 227024 320719
rect 227640 304978 227668 371855
rect 227732 371278 227760 372506
rect 227720 371272 227772 371278
rect 227720 371214 227772 371220
rect 228456 371272 228508 371278
rect 228456 371214 228508 371220
rect 228364 367804 228416 367810
rect 228364 367746 228416 367752
rect 228376 305114 228404 367746
rect 228468 363730 228496 371214
rect 228456 363724 228508 363730
rect 228456 363666 228508 363672
rect 229008 356720 229060 356726
rect 229008 356662 229060 356668
rect 228364 305108 228416 305114
rect 228364 305050 228416 305056
rect 227628 304972 227680 304978
rect 227628 304914 227680 304920
rect 228376 301594 228404 305050
rect 229020 304298 229048 356662
rect 229756 328545 229784 375935
rect 229282 328536 229338 328545
rect 229282 328471 229338 328480
rect 229742 328536 229798 328545
rect 229742 328471 229798 328480
rect 229296 325694 229324 328471
rect 229296 325666 229968 325694
rect 229836 304972 229888 304978
rect 229836 304914 229888 304920
rect 229008 304292 229060 304298
rect 229008 304234 229060 304240
rect 229020 303634 229048 304234
rect 229020 303606 229140 303634
rect 229112 301594 229140 303606
rect 225156 301566 225630 301594
rect 225984 301566 226274 301594
rect 226444 301566 226826 301594
rect 226996 301566 227470 301594
rect 228376 301566 228666 301594
rect 229112 301566 229218 301594
rect 229848 301580 229876 304914
rect 229940 301594 229968 325666
rect 230492 309806 230520 389286
rect 230570 389263 230626 389272
rect 231504 385014 231532 390388
rect 231872 390374 232438 390402
rect 230572 385008 230624 385014
rect 230572 384950 230624 384956
rect 231492 385008 231544 385014
rect 231492 384950 231544 384956
rect 230584 381546 230612 384950
rect 231872 382974 231900 390374
rect 233344 388482 233372 390388
rect 233332 388476 233384 388482
rect 233332 388418 233384 388424
rect 234264 387870 234292 390388
rect 234632 390374 235382 390402
rect 236012 390374 236302 390402
rect 232504 387864 232556 387870
rect 232504 387806 232556 387812
rect 234252 387864 234304 387870
rect 234252 387806 234304 387812
rect 232516 386374 232544 387806
rect 232504 386368 232556 386374
rect 232504 386310 232556 386316
rect 231860 382968 231912 382974
rect 231860 382910 231912 382916
rect 231122 381576 231178 381585
rect 230572 381540 230624 381546
rect 231122 381511 231178 381520
rect 230572 381482 230624 381488
rect 231136 341465 231164 381511
rect 232516 374649 232544 386310
rect 232594 382936 232650 382945
rect 232594 382871 232650 382880
rect 232502 374640 232558 374649
rect 232502 374575 232558 374584
rect 232502 351928 232558 351937
rect 232502 351863 232558 351872
rect 231122 341456 231178 341465
rect 231122 341391 231178 341400
rect 230572 334076 230624 334082
rect 230572 334018 230624 334024
rect 230480 309800 230532 309806
rect 230480 309742 230532 309748
rect 230584 303686 230612 334018
rect 230662 332616 230718 332625
rect 230662 332551 230718 332560
rect 230572 303680 230624 303686
rect 230572 303622 230624 303628
rect 230676 301594 230704 332551
rect 231858 331256 231914 331265
rect 231858 331191 231914 331200
rect 231872 325694 231900 331191
rect 231872 325666 232360 325694
rect 231122 309224 231178 309233
rect 231122 309159 231178 309168
rect 231136 302190 231164 309159
rect 232228 304632 232280 304638
rect 232228 304574 232280 304580
rect 231308 303680 231360 303686
rect 232240 303657 232268 304574
rect 231308 303622 231360 303628
rect 232226 303648 232282 303657
rect 231124 302184 231176 302190
rect 231124 302126 231176 302132
rect 231320 301594 231348 303622
rect 232226 303583 232282 303592
rect 229940 301566 230414 301594
rect 230676 301566 231058 301594
rect 231320 301566 231610 301594
rect 232240 301580 232268 303583
rect 232332 301594 232360 325666
rect 232516 303754 232544 351863
rect 232608 347041 232636 382871
rect 234342 377360 234398 377369
rect 234342 377295 234398 377304
rect 233882 358048 233938 358057
rect 233882 357983 233938 357992
rect 233896 348498 233924 357983
rect 233884 348492 233936 348498
rect 233884 348434 233936 348440
rect 232594 347032 232650 347041
rect 232594 346967 232650 346976
rect 234356 339454 234384 377295
rect 234632 371142 234660 390374
rect 236012 375358 236040 390374
rect 237208 388657 237236 390388
rect 236642 388648 236698 388657
rect 236642 388583 236698 388592
rect 237194 388648 237250 388657
rect 237194 388583 237250 388592
rect 236656 378146 236684 388583
rect 238128 388414 238156 390388
rect 239048 389298 239076 390388
rect 239508 390374 239982 390402
rect 240152 390374 241086 390402
rect 242006 390374 242204 390402
rect 238760 389292 238812 389298
rect 238760 389234 238812 389240
rect 239036 389292 239088 389298
rect 239036 389234 239088 389240
rect 238116 388408 238168 388414
rect 238116 388350 238168 388356
rect 238022 387016 238078 387025
rect 238022 386951 238078 386960
rect 236644 378140 236696 378146
rect 236644 378082 236696 378088
rect 236000 375352 236052 375358
rect 236000 375294 236052 375300
rect 236644 375352 236696 375358
rect 236644 375294 236696 375300
rect 236656 374746 236684 375294
rect 236644 374740 236696 374746
rect 236644 374682 236696 374688
rect 235262 373280 235318 373289
rect 235262 373215 235318 373224
rect 234620 371136 234672 371142
rect 234620 371078 234672 371084
rect 234632 370530 234660 371078
rect 234620 370524 234672 370530
rect 234620 370466 234672 370472
rect 234528 369164 234580 369170
rect 234528 369106 234580 369112
rect 234436 347064 234488 347070
rect 234436 347006 234488 347012
rect 234344 339448 234396 339454
rect 234344 339390 234396 339396
rect 233882 329896 233938 329905
rect 233882 329831 233938 329840
rect 233896 329118 233924 329831
rect 233884 329112 233936 329118
rect 233884 329054 233936 329060
rect 233884 318096 233936 318102
rect 233884 318038 233936 318044
rect 232504 303748 232556 303754
rect 232504 303690 232556 303696
rect 233896 303686 233924 318038
rect 233976 303748 234028 303754
rect 233976 303690 234028 303696
rect 233884 303680 233936 303686
rect 233884 303622 233936 303628
rect 233424 303204 233476 303210
rect 233424 303146 233476 303152
rect 233436 302258 233464 303146
rect 233424 302252 233476 302258
rect 233424 302194 233476 302200
rect 232332 301566 232806 301594
rect 233436 301580 233464 302194
rect 233988 301580 234016 303690
rect 234448 303210 234476 347006
rect 234436 303204 234488 303210
rect 234436 303146 234488 303152
rect 234540 301753 234568 369106
rect 235276 349858 235304 373215
rect 236642 356688 236698 356697
rect 236642 356623 236698 356632
rect 235264 349852 235316 349858
rect 235264 349794 235316 349800
rect 236656 344350 236684 356623
rect 236644 344344 236696 344350
rect 236644 344286 236696 344292
rect 238036 342961 238064 386951
rect 238772 381614 238800 389234
rect 239404 388408 239456 388414
rect 239404 388350 239456 388356
rect 238760 381608 238812 381614
rect 238760 381550 238812 381556
rect 239416 375329 239444 388350
rect 239508 386306 239536 390374
rect 239496 386300 239548 386306
rect 239496 386242 239548 386248
rect 239402 375320 239458 375329
rect 239402 375255 239458 375264
rect 238114 370696 238170 370705
rect 238114 370631 238170 370640
rect 238128 351218 238156 370631
rect 239416 357474 239444 375255
rect 239404 357468 239456 357474
rect 239404 357410 239456 357416
rect 238116 351212 238168 351218
rect 238116 351154 238168 351160
rect 238022 342952 238078 342961
rect 238022 342887 238078 342896
rect 234804 339448 234856 339454
rect 234804 339390 234856 339396
rect 234816 338774 234844 339390
rect 234804 338768 234856 338774
rect 234804 338710 234856 338716
rect 234710 314800 234766 314809
rect 234710 314735 234766 314744
rect 234620 303680 234672 303686
rect 234620 303622 234672 303628
rect 234526 301744 234582 301753
rect 234526 301679 234582 301688
rect 234632 301580 234660 303622
rect 234724 301594 234752 314735
rect 234816 306374 234844 338710
rect 237380 337476 237432 337482
rect 237380 337418 237432 337424
rect 236000 331900 236052 331906
rect 236000 331842 236052 331848
rect 235262 327720 235318 327729
rect 235262 327655 235318 327664
rect 235276 314809 235304 327655
rect 235262 314800 235318 314809
rect 235262 314735 235318 314744
rect 234816 306346 235488 306374
rect 235460 301594 235488 306346
rect 236012 301594 236040 331842
rect 236644 317484 236696 317490
rect 236644 317426 236696 317432
rect 236656 307086 236684 317426
rect 236644 307080 236696 307086
rect 236644 307022 236696 307028
rect 237392 303686 237420 337418
rect 237470 318064 237526 318073
rect 237470 317999 237526 318008
rect 237484 310593 237512 317999
rect 239416 311166 239444 357410
rect 239508 354686 239536 386242
rect 240152 371210 240180 390374
rect 240968 387252 241020 387258
rect 240968 387194 241020 387200
rect 240782 381712 240838 381721
rect 240782 381647 240838 381656
rect 240140 371204 240192 371210
rect 240140 371146 240192 371152
rect 240140 356788 240192 356794
rect 240140 356730 240192 356736
rect 239496 354680 239548 354686
rect 239496 354622 239548 354628
rect 239404 311160 239456 311166
rect 239404 311102 239456 311108
rect 237470 310584 237526 310593
rect 237470 310519 237526 310528
rect 237380 303680 237432 303686
rect 237380 303622 237432 303628
rect 237484 301594 237512 310519
rect 239508 307834 239536 354622
rect 240046 339824 240102 339833
rect 240046 339759 240102 339768
rect 239496 307828 239548 307834
rect 239496 307770 239548 307776
rect 240060 303929 240088 339759
rect 240152 307737 240180 356730
rect 240138 307728 240194 307737
rect 240138 307663 240194 307672
rect 240796 304638 240824 381647
rect 240876 371204 240928 371210
rect 240876 371146 240928 371152
rect 240888 318102 240916 371146
rect 240980 365702 241008 387194
rect 242176 385014 242204 390374
rect 242912 387734 242940 390388
rect 243096 390374 243846 390402
rect 242900 387728 242952 387734
rect 242900 387670 242952 387676
rect 242912 387258 242940 387670
rect 242900 387252 242952 387258
rect 242900 387194 242952 387200
rect 242164 385008 242216 385014
rect 242164 384950 242216 384956
rect 241520 374672 241572 374678
rect 241520 374614 241572 374620
rect 240968 365696 241020 365702
rect 240968 365638 241020 365644
rect 241532 326466 241560 374614
rect 242176 369850 242204 384950
rect 243096 382265 243124 390374
rect 244752 389065 244780 390388
rect 244738 389056 244794 389065
rect 244738 388991 244794 389000
rect 245566 388376 245622 388385
rect 245566 388311 245622 388320
rect 244924 387864 244976 387870
rect 244924 387806 244976 387812
rect 244936 386209 244964 387806
rect 244922 386200 244978 386209
rect 244922 386135 244978 386144
rect 243082 382256 243138 382265
rect 243082 382191 243138 382200
rect 243096 381041 243124 382191
rect 243082 381032 243138 381041
rect 243082 380967 243138 380976
rect 244186 381032 244242 381041
rect 244186 380967 244242 380976
rect 242164 369844 242216 369850
rect 242164 369786 242216 369792
rect 241520 326460 241572 326466
rect 241520 326402 241572 326408
rect 241532 325718 241560 326402
rect 241520 325712 241572 325718
rect 241520 325654 241572 325660
rect 240876 318096 240928 318102
rect 240876 318038 240928 318044
rect 242176 312662 242204 369786
rect 242256 365016 242308 365022
rect 242256 364958 242308 364964
rect 242268 334014 242296 364958
rect 244200 354074 244228 380967
rect 244936 373386 244964 386135
rect 244924 373380 244976 373386
rect 244924 373322 244976 373328
rect 244924 370524 244976 370530
rect 244924 370466 244976 370472
rect 244188 354068 244240 354074
rect 244188 354010 244240 354016
rect 243084 340196 243136 340202
rect 243084 340138 243136 340144
rect 242256 334008 242308 334014
rect 242256 333950 242308 333956
rect 242164 312656 242216 312662
rect 242164 312598 242216 312604
rect 241428 307828 241480 307834
rect 241428 307770 241480 307776
rect 241242 307728 241298 307737
rect 241242 307663 241298 307672
rect 241256 306513 241284 307663
rect 241242 306504 241298 306513
rect 241242 306439 241298 306448
rect 240784 304632 240836 304638
rect 240784 304574 240836 304580
rect 240046 303920 240102 303929
rect 240046 303855 240102 303864
rect 237932 303680 237984 303686
rect 237932 303622 237984 303628
rect 237944 301594 237972 303622
rect 238850 302288 238906 302297
rect 238850 302223 238906 302232
rect 234724 301566 235198 301594
rect 235460 301566 235842 301594
rect 236012 301566 236394 301594
rect 237484 301566 237590 301594
rect 237944 301566 238234 301594
rect 238864 301580 238892 302223
rect 239402 302152 239458 302161
rect 239402 302087 239458 302096
rect 239416 301580 239444 302087
rect 240060 301580 240088 303855
rect 240600 302320 240652 302326
rect 240600 302262 240652 302268
rect 240612 301580 240640 302262
rect 241256 301580 241284 306439
rect 241440 302433 241468 307770
rect 241794 305008 241850 305017
rect 241794 304943 241850 304952
rect 241426 302424 241482 302433
rect 241426 302359 241482 302368
rect 241808 301580 241836 304943
rect 242268 303686 242296 333950
rect 242348 326460 242400 326466
rect 242348 326402 242400 326408
rect 242256 303680 242308 303686
rect 242256 303622 242308 303628
rect 242360 301578 242388 326402
rect 242440 304360 242492 304366
rect 242440 304302 242492 304308
rect 242452 301580 242480 304302
rect 243096 301617 243124 340138
rect 244464 336048 244516 336054
rect 244464 335990 244516 335996
rect 243176 328500 243228 328506
rect 243176 328442 243228 328448
rect 243082 301608 243138 301617
rect 242348 301572 242400 301578
rect 243018 301566 243082 301594
rect 243188 301594 243216 328442
rect 244370 310448 244426 310457
rect 244370 310383 244426 310392
rect 244384 309233 244412 310383
rect 244370 309224 244426 309233
rect 244370 309159 244426 309168
rect 244188 303680 244240 303686
rect 244188 303622 244240 303628
rect 243188 301566 243662 301594
rect 244200 301580 244228 303622
rect 243082 301543 243138 301552
rect 242348 301514 242400 301520
rect 243096 301483 243124 301543
rect 236734 301472 236790 301481
rect 236790 301430 237038 301458
rect 244384 301442 244412 309159
rect 244476 305833 244504 335990
rect 244936 334665 244964 370466
rect 245016 344412 245068 344418
rect 245016 344354 245068 344360
rect 245028 335374 245056 344354
rect 245016 335368 245068 335374
rect 245016 335310 245068 335316
rect 244922 334656 244978 334665
rect 244922 334591 244978 334600
rect 245028 310457 245056 335310
rect 245014 310448 245070 310457
rect 245014 310383 245070 310392
rect 245580 306513 245608 388311
rect 245672 387870 245700 390388
rect 245764 390374 246606 390402
rect 247052 390374 247710 390402
rect 245660 387864 245712 387870
rect 245660 387806 245712 387812
rect 245764 373998 245792 390374
rect 245844 388476 245896 388482
rect 245844 388418 245896 388424
rect 245856 386374 245884 388418
rect 245844 386368 245896 386374
rect 245844 386310 245896 386316
rect 246948 386368 247000 386374
rect 246948 386310 247000 386316
rect 245752 373992 245804 373998
rect 245752 373934 245804 373940
rect 245764 372638 245792 373934
rect 245752 372632 245804 372638
rect 245752 372574 245804 372580
rect 246304 372632 246356 372638
rect 246304 372574 246356 372580
rect 246316 330546 246344 372574
rect 246304 330540 246356 330546
rect 246304 330482 246356 330488
rect 245660 329928 245712 329934
rect 245660 329870 245712 329876
rect 245566 306504 245622 306513
rect 245566 306439 245622 306448
rect 245580 306374 245608 306439
rect 245304 306346 245608 306374
rect 244462 305824 244518 305833
rect 244462 305759 244518 305768
rect 244476 305017 244504 305759
rect 244462 305008 244518 305017
rect 244462 304943 244518 304952
rect 245304 301594 245332 306346
rect 244858 301566 245332 301594
rect 245672 301594 245700 329870
rect 246396 323672 246448 323678
rect 246396 323614 246448 323620
rect 246304 317484 246356 317490
rect 246304 317426 246356 317432
rect 246210 307048 246266 307057
rect 246210 306983 246266 306992
rect 246224 301594 246252 306983
rect 246316 302161 246344 317426
rect 246408 307057 246436 323614
rect 246394 307048 246450 307057
rect 246394 306983 246450 306992
rect 246960 304337 246988 386310
rect 247052 372609 247080 390374
rect 248616 389065 248644 390388
rect 249536 389065 249564 390388
rect 248602 389056 248658 389065
rect 248602 388991 248658 389000
rect 249522 389056 249578 389065
rect 249522 388991 249578 389000
rect 247222 388512 247278 388521
rect 247222 388447 247278 388456
rect 247684 388476 247736 388482
rect 247130 378720 247186 378729
rect 247130 378655 247186 378664
rect 247144 376718 247172 378655
rect 247132 376712 247184 376718
rect 247132 376654 247184 376660
rect 247038 372600 247094 372609
rect 247038 372535 247094 372544
rect 247052 371210 247080 372535
rect 247040 371204 247092 371210
rect 247040 371146 247092 371152
rect 247144 332654 247172 376654
rect 247236 366353 247264 388447
rect 247684 388418 247736 388424
rect 247696 379438 247724 388418
rect 249536 383654 249564 388991
rect 249536 383626 249656 383654
rect 247684 379432 247736 379438
rect 247684 379374 247736 379380
rect 249062 374640 249118 374649
rect 249062 374575 249118 374584
rect 248328 371204 248380 371210
rect 248328 371146 248380 371152
rect 247222 366344 247278 366353
rect 247222 366279 247278 366288
rect 247132 332648 247184 332654
rect 247132 332590 247184 332596
rect 247684 332648 247736 332654
rect 247684 332590 247736 332596
rect 247696 307873 247724 332590
rect 248340 330449 248368 371146
rect 248972 365696 249024 365702
rect 248972 365638 249024 365644
rect 248326 330440 248382 330449
rect 248326 330375 248382 330384
rect 247776 314016 247828 314022
rect 247776 313958 247828 313964
rect 247682 307864 247738 307873
rect 247682 307799 247738 307808
rect 246946 304328 247002 304337
rect 246946 304263 247002 304272
rect 247222 304192 247278 304201
rect 247222 304127 247278 304136
rect 246302 302152 246358 302161
rect 246302 302087 246358 302096
rect 245672 301566 246054 301594
rect 246224 301566 246606 301594
rect 247236 301580 247264 304127
rect 247696 301594 247724 307799
rect 247788 304298 247816 313958
rect 248694 311808 248750 311817
rect 248694 311743 248750 311752
rect 248602 310992 248658 311001
rect 248602 310927 248658 310936
rect 247776 304292 247828 304298
rect 247776 304234 247828 304240
rect 248616 301594 248644 310927
rect 248708 303686 248736 311743
rect 248696 303680 248748 303686
rect 248696 303622 248748 303628
rect 247696 301566 247802 301594
rect 248446 301566 248644 301594
rect 245120 301442 245410 301458
rect 244372 301436 244424 301442
rect 236734 301407 236790 301416
rect 244372 301378 244424 301384
rect 245108 301436 245410 301442
rect 245160 301430 245410 301436
rect 245108 301378 245160 301384
rect 218206 301172 218468 301186
rect 218206 301158 218454 301172
rect 218150 301135 218206 301144
rect 227720 300960 227772 300966
rect 216864 300902 216916 300908
rect 217874 300928 217930 300937
rect 199070 300886 199226 300900
rect 199014 300863 199070 300872
rect 248984 300914 249012 365638
rect 249076 329225 249104 374575
rect 249628 361622 249656 383626
rect 249720 373994 249748 390895
rect 251824 390584 251876 390590
rect 251824 390526 251876 390532
rect 250470 390374 250760 390402
rect 250442 389464 250498 389473
rect 250442 389399 250498 389408
rect 249720 373969 249840 373994
rect 249706 373966 249840 373969
rect 249706 373960 249762 373966
rect 249706 373895 249762 373904
rect 249708 371884 249760 371890
rect 249708 371826 249760 371832
rect 249616 361616 249668 361622
rect 249614 361584 249616 361593
rect 249668 361584 249670 361593
rect 249614 361519 249670 361528
rect 249062 329216 249118 329225
rect 249062 329151 249118 329160
rect 249616 313336 249668 313342
rect 249616 313278 249668 313284
rect 249628 311817 249656 313278
rect 249614 311808 249670 311817
rect 249614 311743 249670 311752
rect 249720 311001 249748 371826
rect 249812 365702 249840 373966
rect 250456 368393 250484 389399
rect 250732 389094 250760 390374
rect 250720 389088 250772 389094
rect 250720 389030 250772 389036
rect 250732 380866 250760 389030
rect 251376 388482 251404 390388
rect 251364 388476 251416 388482
rect 251364 388418 251416 388424
rect 250720 380860 250772 380866
rect 250720 380802 250772 380808
rect 251836 374678 251864 390526
rect 252310 390374 252508 390402
rect 252008 387864 252060 387870
rect 252008 387806 252060 387812
rect 251824 374672 251876 374678
rect 251824 374614 251876 374620
rect 251916 373312 251968 373318
rect 251916 373254 251968 373260
rect 250442 368384 250498 368393
rect 250442 368319 250498 368328
rect 249800 365696 249852 365702
rect 249800 365638 249852 365644
rect 250456 344350 250484 368319
rect 251824 363724 251876 363730
rect 251824 363666 251876 363672
rect 250444 344344 250496 344350
rect 250444 344286 250496 344292
rect 249890 331256 249946 331265
rect 249890 331191 249946 331200
rect 249904 327758 249932 331191
rect 249892 327752 249944 327758
rect 249892 327694 249944 327700
rect 251836 326466 251864 363666
rect 251928 338842 251956 373254
rect 252020 362914 252048 387806
rect 252480 384985 252508 390374
rect 253400 389162 253428 390388
rect 253388 389156 253440 389162
rect 253388 389098 253440 389104
rect 253400 387870 253428 389098
rect 253388 387864 253440 387870
rect 253388 387806 253440 387812
rect 253584 386306 253612 391274
rect 253676 389094 253704 392566
rect 253938 392048 253994 392057
rect 253938 391983 253994 391992
rect 253664 389088 253716 389094
rect 253664 389030 253716 389036
rect 253572 386300 253624 386306
rect 253572 386242 253624 386248
rect 252466 384976 252522 384985
rect 252466 384911 252522 384920
rect 252480 378826 252508 384911
rect 252468 378820 252520 378826
rect 252468 378762 252520 378768
rect 253952 365673 253980 391983
rect 254044 389473 254072 395519
rect 254030 389464 254086 389473
rect 254030 389399 254086 389408
rect 254136 366382 254164 405311
rect 254228 389337 254256 427887
rect 254320 392873 254348 458798
rect 254596 449274 254624 515374
rect 254688 458862 254716 525098
rect 254676 458856 254728 458862
rect 254676 458798 254728 458804
rect 255228 451308 255280 451314
rect 255228 451250 255280 451256
rect 255240 450566 255268 451250
rect 255228 450560 255280 450566
rect 255228 450502 255280 450508
rect 254584 449268 254636 449274
rect 254584 449210 254636 449216
rect 254490 447536 254546 447545
rect 254490 447471 254492 447480
rect 254544 447471 254546 447480
rect 254492 447442 254544 447448
rect 255332 415177 255360 578122
rect 255410 577688 255466 577697
rect 255410 577623 255466 577632
rect 255424 577114 255452 577623
rect 255412 577108 255464 577114
rect 255412 577050 255464 577056
rect 255410 577008 255466 577017
rect 255410 576943 255466 576952
rect 255424 576910 255452 576943
rect 255412 576904 255464 576910
rect 255412 576846 255464 576852
rect 255410 575920 255466 575929
rect 255410 575855 255466 575864
rect 255424 575550 255452 575855
rect 255412 575544 255464 575550
rect 255412 575486 255464 575492
rect 255410 574696 255466 574705
rect 255410 574631 255466 574640
rect 255424 574122 255452 574631
rect 255594 574152 255650 574161
rect 255412 574116 255464 574122
rect 255594 574087 255650 574096
rect 255412 574058 255464 574064
rect 255502 571976 255558 571985
rect 255502 571911 255558 571920
rect 255410 571568 255466 571577
rect 255410 571503 255466 571512
rect 255424 571470 255452 571503
rect 255412 571464 255464 571470
rect 255412 571406 255464 571412
rect 255516 571402 255544 571911
rect 255504 571396 255556 571402
rect 255504 571338 255556 571344
rect 255412 571328 255464 571334
rect 255412 571270 255464 571276
rect 255424 570625 255452 571270
rect 255410 570616 255466 570625
rect 255410 570551 255466 570560
rect 255502 569256 255558 569265
rect 255502 569191 255558 569200
rect 255410 568712 255466 568721
rect 255516 568682 255544 569191
rect 255410 568647 255466 568656
rect 255504 568676 255556 568682
rect 255424 568614 255452 568647
rect 255504 568618 255556 568624
rect 255412 568608 255464 568614
rect 255412 568550 255464 568556
rect 255608 567194 255636 574087
rect 255976 573374 256004 587959
rect 256712 586514 256740 595190
rect 256712 586486 256832 586514
rect 255964 573368 256016 573374
rect 255964 573310 256016 573316
rect 255686 572928 255742 572937
rect 255686 572863 255742 572872
rect 255700 567866 255728 572863
rect 255688 567860 255740 567866
rect 255688 567802 255740 567808
rect 255424 567166 255636 567194
rect 255424 431254 255452 567166
rect 255594 566264 255650 566273
rect 255594 566199 255650 566208
rect 255502 565992 255558 566001
rect 255502 565927 255504 565936
rect 255556 565927 255558 565936
rect 255504 565898 255556 565904
rect 255608 565894 255636 566199
rect 255596 565888 255648 565894
rect 255596 565830 255648 565836
rect 255502 564768 255558 564777
rect 255502 564703 255558 564712
rect 255516 564466 255544 564703
rect 255504 564460 255556 564466
rect 255504 564402 255556 564408
rect 255686 561776 255742 561785
rect 255686 561711 255742 561720
rect 255502 560824 255558 560833
rect 255502 560759 255558 560768
rect 255516 560318 255544 560759
rect 255504 560312 255556 560318
rect 255504 560254 255556 560260
rect 255594 559600 255650 559609
rect 255594 559535 255650 559544
rect 255502 559192 255558 559201
rect 255502 559127 255558 559136
rect 255516 559026 255544 559127
rect 255504 559020 255556 559026
rect 255504 558962 255556 558968
rect 255608 558958 255636 559535
rect 255596 558952 255648 558958
rect 255596 558894 255648 558900
rect 255700 558770 255728 561711
rect 255516 558742 255728 558770
rect 255516 546938 255544 558742
rect 255594 557968 255650 557977
rect 255594 557903 255650 557912
rect 255608 557598 255636 557903
rect 255596 557592 255648 557598
rect 255596 557534 255648 557540
rect 255594 556880 255650 556889
rect 255594 556815 255650 556824
rect 255608 556238 255636 556815
rect 255596 556232 255648 556238
rect 255596 556174 255648 556180
rect 255686 554160 255742 554169
rect 255686 554095 255742 554104
rect 255594 553616 255650 553625
rect 255594 553551 255650 553560
rect 255608 553518 255636 553551
rect 255596 553512 255648 553518
rect 255596 553454 255648 553460
rect 255700 553450 255728 554095
rect 255688 553444 255740 553450
rect 255688 553386 255740 553392
rect 255594 552800 255650 552809
rect 255594 552735 255650 552744
rect 255608 552702 255636 552735
rect 255596 552696 255648 552702
rect 255596 552638 255648 552644
rect 255594 550896 255650 550905
rect 255594 550831 255650 550840
rect 255608 550730 255636 550831
rect 255596 550724 255648 550730
rect 255596 550666 255648 550672
rect 255594 549944 255650 549953
rect 255594 549879 255596 549888
rect 255648 549879 255650 549888
rect 255596 549850 255648 549856
rect 255594 548448 255650 548457
rect 255594 548383 255650 548392
rect 255608 547942 255636 548383
rect 255596 547936 255648 547942
rect 255596 547878 255648 547884
rect 255870 547904 255926 547913
rect 255870 547839 255926 547848
rect 255516 546910 255820 546938
rect 255502 546816 255558 546825
rect 255502 546751 255558 546760
rect 255516 546514 255544 546751
rect 255504 546508 255556 546514
rect 255504 546450 255556 546456
rect 255502 545864 255558 545873
rect 255502 545799 255558 545808
rect 255516 545290 255544 545799
rect 255504 545284 255556 545290
rect 255504 545226 255556 545232
rect 255594 542872 255650 542881
rect 255594 542807 255650 542816
rect 255608 542502 255636 542807
rect 255596 542496 255648 542502
rect 255502 542464 255558 542473
rect 255596 542438 255648 542444
rect 255502 542399 255504 542408
rect 255556 542399 255558 542408
rect 255504 542370 255556 542376
rect 255502 540152 255558 540161
rect 255502 540087 255558 540096
rect 255516 539646 255544 540087
rect 255504 539640 255556 539646
rect 255504 539582 255556 539588
rect 255502 539472 255558 539481
rect 255502 539407 255558 539416
rect 255516 538354 255544 539407
rect 255792 539306 255820 546910
rect 255780 539300 255832 539306
rect 255780 539242 255832 539248
rect 255504 538348 255556 538354
rect 255504 538290 255556 538296
rect 255884 533458 255912 547839
rect 256606 543824 256662 543833
rect 256662 543782 256740 543810
rect 256606 543759 256662 543768
rect 255872 533452 255924 533458
rect 255872 533394 255924 533400
rect 255504 471300 255556 471306
rect 255504 471242 255556 471248
rect 255516 447250 255544 471242
rect 255594 457464 255650 457473
rect 255594 457399 255650 457408
rect 255608 449206 255636 457399
rect 255688 449608 255740 449614
rect 255688 449550 255740 449556
rect 255596 449200 255648 449206
rect 255596 449142 255648 449148
rect 255608 448905 255636 449142
rect 255594 448896 255650 448905
rect 255594 448831 255650 448840
rect 255516 447222 255636 447250
rect 255504 447092 255556 447098
rect 255504 447034 255556 447040
rect 255516 446185 255544 447034
rect 255502 446176 255558 446185
rect 255502 446111 255558 446120
rect 255608 444825 255636 447222
rect 255594 444816 255650 444825
rect 255594 444751 255650 444760
rect 255504 443692 255556 443698
rect 255504 443634 255556 443640
rect 255516 443465 255544 443634
rect 255502 443456 255558 443465
rect 255502 443391 255558 443400
rect 255700 442105 255728 449550
rect 255686 442096 255742 442105
rect 255686 442031 255742 442040
rect 255504 439544 255556 439550
rect 255504 439486 255556 439492
rect 255516 439113 255544 439486
rect 255502 439104 255558 439113
rect 255502 439039 255558 439048
rect 255504 438184 255556 438190
rect 255504 438126 255556 438132
rect 255516 437753 255544 438126
rect 255502 437744 255558 437753
rect 255502 437679 255558 437688
rect 255502 437608 255558 437617
rect 255502 437543 255558 437552
rect 255516 437510 255544 437543
rect 255504 437504 255556 437510
rect 255504 437446 255556 437452
rect 255516 436393 255544 437446
rect 255700 436762 255728 442031
rect 255688 436756 255740 436762
rect 255688 436698 255740 436704
rect 255502 436384 255558 436393
rect 255502 436319 255558 436328
rect 255504 435396 255556 435402
rect 255504 435338 255556 435344
rect 255516 435033 255544 435338
rect 255502 435024 255558 435033
rect 255502 434959 255558 434968
rect 255504 434716 255556 434722
rect 255504 434658 255556 434664
rect 255516 433673 255544 434658
rect 255502 433664 255558 433673
rect 255502 433599 255558 433608
rect 255964 432676 256016 432682
rect 255964 432618 256016 432624
rect 255976 432041 256004 432618
rect 255962 432032 256018 432041
rect 255962 431967 256018 431976
rect 255412 431248 255464 431254
rect 255412 431190 255464 431196
rect 255424 430681 255452 431190
rect 255410 430672 255466 430681
rect 255410 430607 255466 430616
rect 255410 426592 255466 426601
rect 255410 426527 255466 426536
rect 255424 426494 255452 426527
rect 255412 426488 255464 426494
rect 255412 426430 255464 426436
rect 255504 426420 255556 426426
rect 255504 426362 255556 426368
rect 255516 425241 255544 426362
rect 255502 425232 255558 425241
rect 255502 425167 255558 425176
rect 255502 423600 255558 423609
rect 255502 423535 255558 423544
rect 255516 422346 255544 423535
rect 255504 422340 255556 422346
rect 255504 422282 255556 422288
rect 255502 422240 255558 422249
rect 255502 422175 255558 422184
rect 255516 420986 255544 422175
rect 255504 420980 255556 420986
rect 255504 420922 255556 420928
rect 255502 420880 255558 420889
rect 255502 420815 255558 420824
rect 255516 419558 255544 420815
rect 255504 419552 255556 419558
rect 255410 419520 255466 419529
rect 255504 419494 255556 419500
rect 255410 419455 255412 419464
rect 255464 419455 255466 419464
rect 255412 419426 255464 419432
rect 255410 418160 255466 418169
rect 255410 418095 255466 418104
rect 255424 417450 255452 418095
rect 255412 417444 255464 417450
rect 255412 417386 255464 417392
rect 255412 416832 255464 416838
rect 255410 416800 255412 416809
rect 255464 416800 255466 416809
rect 255410 416735 255466 416744
rect 255318 415168 255374 415177
rect 255318 415103 255374 415112
rect 255412 413840 255464 413846
rect 255410 413808 255412 413817
rect 255464 413808 255466 413817
rect 255410 413743 255466 413752
rect 255412 412480 255464 412486
rect 255410 412448 255412 412457
rect 255464 412448 255466 412457
rect 255410 412383 255466 412392
rect 255502 411088 255558 411097
rect 255502 411023 255558 411032
rect 255410 409728 255466 409737
rect 255410 409663 255466 409672
rect 255424 408542 255452 409663
rect 255412 408536 255464 408542
rect 255412 408478 255464 408484
rect 255410 408368 255466 408377
rect 255410 408303 255466 408312
rect 255424 407862 255452 408303
rect 255412 407856 255464 407862
rect 255412 407798 255464 407804
rect 255516 407794 255544 411023
rect 255504 407788 255556 407794
rect 255504 407730 255556 407736
rect 255502 407008 255558 407017
rect 255502 406943 255558 406952
rect 255516 405754 255544 406943
rect 255504 405748 255556 405754
rect 255504 405690 255556 405696
rect 255320 402960 255372 402966
rect 255320 402902 255372 402908
rect 255332 402665 255360 402902
rect 255318 402656 255374 402665
rect 255318 402591 255374 402600
rect 255410 401296 255466 401305
rect 255410 401231 255466 401240
rect 255424 400246 255452 401231
rect 255412 400240 255464 400246
rect 255412 400182 255464 400188
rect 255410 399936 255466 399945
rect 255410 399871 255466 399880
rect 255424 398886 255452 399871
rect 255412 398880 255464 398886
rect 255412 398822 255464 398828
rect 255410 398576 255466 398585
rect 255410 398511 255466 398520
rect 255424 398274 255452 398511
rect 255412 398268 255464 398274
rect 255412 398210 255464 398216
rect 255502 394224 255558 394233
rect 255502 394159 255558 394168
rect 255516 393378 255544 394159
rect 255504 393372 255556 393378
rect 255504 393314 255556 393320
rect 254306 392864 254362 392873
rect 254306 392799 254362 392808
rect 254320 392018 254348 392799
rect 254308 392012 254360 392018
rect 254308 391954 254360 391960
rect 255320 392012 255372 392018
rect 255320 391954 255372 391960
rect 254214 389328 254270 389337
rect 254214 389263 254270 389272
rect 254124 366376 254176 366382
rect 254124 366318 254176 366324
rect 253938 365664 253994 365673
rect 253938 365599 253994 365608
rect 252008 362908 252060 362914
rect 252008 362850 252060 362856
rect 253952 344418 253980 365599
rect 255332 358766 255360 391954
rect 256712 363633 256740 543782
rect 256804 530641 256832 586486
rect 259472 584458 259500 612750
rect 263600 603152 263652 603158
rect 263600 603094 263652 603100
rect 261024 593428 261076 593434
rect 261024 593370 261076 593376
rect 260748 585200 260800 585206
rect 260748 585142 260800 585148
rect 259460 584452 259512 584458
rect 259460 584394 259512 584400
rect 259368 583092 259420 583098
rect 259368 583034 259420 583040
rect 259380 582418 259408 583034
rect 258172 582412 258224 582418
rect 258172 582354 258224 582360
rect 259368 582412 259420 582418
rect 259368 582354 259420 582360
rect 256882 567488 256938 567497
rect 256882 567423 256938 567432
rect 256896 534750 256924 567423
rect 258080 549908 258132 549914
rect 258080 549850 258132 549856
rect 256884 534744 256936 534750
rect 256884 534686 256936 534692
rect 256790 530632 256846 530641
rect 256790 530567 256846 530576
rect 256792 497480 256844 497486
rect 256792 497422 256844 497428
rect 256698 363624 256754 363633
rect 256698 363559 256754 363568
rect 255320 358760 255372 358766
rect 255320 358702 255372 358708
rect 253940 344412 253992 344418
rect 253940 344354 253992 344360
rect 253940 342916 253992 342922
rect 253940 342858 253992 342864
rect 251916 338836 251968 338842
rect 251916 338778 251968 338784
rect 252008 337476 252060 337482
rect 252008 337418 252060 337424
rect 251824 326460 251876 326466
rect 251824 326402 251876 326408
rect 251916 326392 251968 326398
rect 251916 326334 251968 326340
rect 250994 320240 251050 320249
rect 250994 320175 251050 320184
rect 251008 317490 251036 320175
rect 251824 320136 251876 320142
rect 251824 320078 251876 320084
rect 251836 318850 251864 320078
rect 251824 318844 251876 318850
rect 251824 318786 251876 318792
rect 250996 317484 251048 317490
rect 250996 317426 251048 317432
rect 249706 310992 249762 311001
rect 249706 310927 249762 310936
rect 249720 310593 249748 310927
rect 249706 310584 249762 310593
rect 249706 310519 249762 310528
rect 249340 303680 249392 303686
rect 249340 303622 249392 303628
rect 249352 301594 249380 303622
rect 250166 302424 250222 302433
rect 250166 302359 250222 302368
rect 249352 301566 249642 301594
rect 250180 301580 250208 302359
rect 251836 301753 251864 318786
rect 251928 304842 251956 326334
rect 252020 320142 252048 337418
rect 253204 329112 253256 329118
rect 253204 329054 253256 329060
rect 252466 321600 252522 321609
rect 252466 321535 252522 321544
rect 252008 320136 252060 320142
rect 252008 320078 252060 320084
rect 252480 306374 252508 321535
rect 252744 312656 252796 312662
rect 252744 312598 252796 312604
rect 252652 309800 252704 309806
rect 252652 309742 252704 309748
rect 252388 306346 252508 306374
rect 251916 304836 251968 304842
rect 251916 304778 251968 304784
rect 252006 302424 252062 302433
rect 252006 302359 252062 302368
rect 251822 301744 251878 301753
rect 251822 301679 251878 301688
rect 251730 301200 251786 301209
rect 252020 301186 252048 302359
rect 252388 302234 252416 306346
rect 252468 305108 252520 305114
rect 252468 305050 252520 305056
rect 252480 304366 252508 305050
rect 252468 304360 252520 304366
rect 252468 304302 252520 304308
rect 252558 304328 252614 304337
rect 252558 304263 252614 304272
rect 252572 303793 252600 304263
rect 252558 303784 252614 303793
rect 252558 303719 252614 303728
rect 252388 302206 252508 302234
rect 251786 301172 252048 301186
rect 251786 301158 252034 301172
rect 251730 301135 251786 301144
rect 250994 301064 251050 301073
rect 250838 301022 250994 301050
rect 250994 300999 251050 301008
rect 249248 300960 249300 300966
rect 227772 300908 228022 300914
rect 227720 300902 228022 300908
rect 227732 300886 228022 300902
rect 248984 300908 249248 300914
rect 251638 300928 251694 300937
rect 248984 300902 249300 300908
rect 248984 300900 249288 300902
rect 248998 300886 249288 300900
rect 251390 300886 251638 300914
rect 217874 300863 217930 300872
rect 251638 300863 251694 300872
rect 252480 300150 252508 302206
rect 252572 301580 252600 303719
rect 252468 300144 252520 300150
rect 252468 300086 252520 300092
rect 252664 299474 252692 309742
rect 252756 306374 252784 312598
rect 253216 311273 253244 329054
rect 253386 325816 253442 325825
rect 253386 325751 253442 325760
rect 253400 321473 253428 325751
rect 253386 321464 253442 321473
rect 253386 321399 253442 321408
rect 253202 311264 253258 311273
rect 253202 311199 253258 311208
rect 253386 311128 253442 311137
rect 253386 311063 253442 311072
rect 252756 306346 252876 306374
rect 252848 302234 252876 306346
rect 253400 305046 253428 311063
rect 253388 305040 253440 305046
rect 253388 304982 253440 304988
rect 252848 302206 252968 302234
rect 252664 299446 252876 299474
rect 193678 299432 193734 299441
rect 193678 299367 193734 299376
rect 252848 298081 252876 299446
rect 252834 298072 252890 298081
rect 252834 298007 252890 298016
rect 252834 297664 252890 297673
rect 252572 297622 252834 297650
rect 193402 269376 193458 269385
rect 193402 269311 193458 269320
rect 193416 269142 193444 269311
rect 193404 269136 193456 269142
rect 193404 269078 193456 269084
rect 192576 268388 192628 268394
rect 192576 268330 192628 268336
rect 191194 268288 191250 268297
rect 191194 268223 191250 268232
rect 190644 256692 190696 256698
rect 190644 256634 190696 256640
rect 190656 256329 190684 256634
rect 190642 256320 190698 256329
rect 190642 256255 190698 256264
rect 190642 254144 190698 254153
rect 190642 254079 190698 254088
rect 190656 253978 190684 254079
rect 190644 253972 190696 253978
rect 190644 253914 190696 253920
rect 190380 246316 190500 246344
rect 189998 237960 190054 237969
rect 189998 237895 190054 237904
rect 189724 227112 189776 227118
rect 189724 227054 189776 227060
rect 189080 207664 189132 207670
rect 189080 207606 189132 207612
rect 189724 193860 189776 193866
rect 189724 193802 189776 193808
rect 188896 157344 188948 157350
rect 188896 157286 188948 157292
rect 188436 156052 188488 156058
rect 188436 155994 188488 156000
rect 188342 155272 188398 155281
rect 188342 155207 188398 155216
rect 187700 154692 187752 154698
rect 187700 154634 187752 154640
rect 187712 153785 187740 154634
rect 187698 153776 187754 153785
rect 187698 153711 187754 153720
rect 187700 146940 187752 146946
rect 187700 146882 187752 146888
rect 187712 145897 187740 146882
rect 187698 145888 187754 145897
rect 187698 145823 187754 145832
rect 187700 135312 187752 135318
rect 187700 135254 187752 135260
rect 187712 133278 187740 135254
rect 188448 134910 188476 155994
rect 188436 134904 188488 134910
rect 188436 134846 188488 134852
rect 187700 133272 187752 133278
rect 187700 133214 187752 133220
rect 188908 131481 188936 157286
rect 189632 151156 189684 151162
rect 189632 151098 189684 151104
rect 189644 149705 189672 151098
rect 189078 149696 189134 149705
rect 189078 149631 189134 149640
rect 189630 149696 189686 149705
rect 189630 149631 189686 149640
rect 188986 147792 189042 147801
rect 188986 147727 189042 147736
rect 188894 131472 188950 131481
rect 188894 131407 188950 131416
rect 189000 121446 189028 147727
rect 189092 121650 189120 149631
rect 189170 134600 189226 134609
rect 189170 134535 189172 134544
rect 189224 134535 189226 134544
rect 189172 134506 189224 134512
rect 189080 121644 189132 121650
rect 189080 121586 189132 121592
rect 188988 121440 189040 121446
rect 188988 121382 189040 121388
rect 189092 121258 189120 121586
rect 189000 121230 189120 121258
rect 187700 119400 187752 119406
rect 187700 119342 187752 119348
rect 187712 114510 187740 119342
rect 189000 118658 189028 121230
rect 188988 118652 189040 118658
rect 188988 118594 189040 118600
rect 188436 116136 188488 116142
rect 188436 116078 188488 116084
rect 188344 114572 188396 114578
rect 188344 114514 188396 114520
rect 187700 114504 187752 114510
rect 187700 114446 187752 114452
rect 187608 108928 187660 108934
rect 187608 108870 187660 108876
rect 187608 105596 187660 105602
rect 187608 105538 187660 105544
rect 186964 101448 187016 101454
rect 186964 101390 187016 101396
rect 186318 89720 186374 89729
rect 186318 89655 186374 89664
rect 186976 82754 187004 101390
rect 186964 82748 187016 82754
rect 186964 82690 187016 82696
rect 186964 78668 187016 78674
rect 186964 78610 187016 78616
rect 186976 70281 187004 78610
rect 187620 71058 187648 105538
rect 187698 93120 187754 93129
rect 187698 93055 187754 93064
rect 187712 87961 187740 93055
rect 187698 87952 187754 87961
rect 187698 87887 187754 87896
rect 188356 73137 188384 114514
rect 188448 111110 188476 116078
rect 189736 115977 189764 193802
rect 190472 162217 190500 246316
rect 191104 242888 191156 242894
rect 191104 242830 191156 242836
rect 191116 179790 191144 242830
rect 191208 238649 191236 268223
rect 191562 266112 191618 266121
rect 191562 266047 191618 266056
rect 191576 265674 191604 266047
rect 191564 265668 191616 265674
rect 191564 265610 191616 265616
rect 191746 265024 191802 265033
rect 191746 264959 191748 264968
rect 191800 264959 191802 264968
rect 191748 264930 191800 264936
rect 191748 264172 191800 264178
rect 191748 264114 191800 264120
rect 191760 263945 191788 264114
rect 191746 263936 191802 263945
rect 191746 263871 191802 263880
rect 191746 262848 191802 262857
rect 191746 262783 191802 262792
rect 191760 262274 191788 262783
rect 191748 262268 191800 262274
rect 191748 262210 191800 262216
rect 191564 262200 191616 262206
rect 191564 262142 191616 262148
rect 191576 261769 191604 262142
rect 191562 261760 191618 261769
rect 191562 261695 191618 261704
rect 191748 260160 191800 260166
rect 191748 260102 191800 260108
rect 191760 259593 191788 260102
rect 191746 259584 191802 259593
rect 191746 259519 191802 259528
rect 191654 252648 191710 252657
rect 191654 252583 191710 252592
rect 191564 251184 191616 251190
rect 191564 251126 191616 251132
rect 191576 250889 191604 251126
rect 191562 250880 191618 250889
rect 191562 250815 191618 250824
rect 191668 249801 191696 252583
rect 191746 251968 191802 251977
rect 191746 251903 191802 251912
rect 191760 251870 191788 251903
rect 191748 251864 191800 251870
rect 191748 251806 191800 251812
rect 191654 249792 191710 249801
rect 191654 249727 191710 249736
rect 191668 249082 191696 249727
rect 191656 249076 191708 249082
rect 191656 249018 191708 249024
rect 191288 248872 191340 248878
rect 191288 248814 191340 248820
rect 191194 238640 191250 238649
rect 191194 238575 191250 238584
rect 191300 224262 191328 248814
rect 191746 247616 191802 247625
rect 191746 247551 191802 247560
rect 191760 247110 191788 247551
rect 191748 247104 191800 247110
rect 191748 247046 191800 247052
rect 192484 246356 192536 246362
rect 192484 246298 192536 246304
rect 191746 243264 191802 243273
rect 191746 243199 191802 243208
rect 191760 242962 191788 243199
rect 191748 242956 191800 242962
rect 191748 242898 191800 242904
rect 192022 240136 192078 240145
rect 192022 240071 192078 240080
rect 192036 237969 192064 240071
rect 192022 237960 192078 237969
rect 192022 237895 192078 237904
rect 191288 224256 191340 224262
rect 191288 224198 191340 224204
rect 192496 180033 192524 246298
rect 192588 234530 192616 268330
rect 193220 260228 193272 260234
rect 193220 260170 193272 260176
rect 192668 253224 192720 253230
rect 192668 253166 192720 253172
rect 192680 242078 192708 253166
rect 193128 244928 193180 244934
rect 193128 244870 193180 244876
rect 192668 242072 192720 242078
rect 192668 242014 192720 242020
rect 193140 240786 193168 244870
rect 193128 240780 193180 240786
rect 193128 240722 193180 240728
rect 192576 234524 192628 234530
rect 192576 234466 192628 234472
rect 192576 202156 192628 202162
rect 192576 202098 192628 202104
rect 192482 180024 192538 180033
rect 192482 179959 192538 179968
rect 191104 179784 191156 179790
rect 191104 179726 191156 179732
rect 192482 165744 192538 165753
rect 192482 165679 192538 165688
rect 190458 162208 190514 162217
rect 190458 162143 190514 162152
rect 191838 159352 191894 159361
rect 191838 159287 191894 159296
rect 191852 153270 191880 159287
rect 192496 158710 192524 165679
rect 192588 159361 192616 202098
rect 193126 162072 193182 162081
rect 193126 162007 193182 162016
rect 192574 159352 192630 159361
rect 192574 159287 192630 159296
rect 192484 158704 192536 158710
rect 192484 158646 192536 158652
rect 192496 157298 192524 158646
rect 192496 157270 192616 157298
rect 192484 153876 192536 153882
rect 192484 153818 192536 153824
rect 191840 153264 191892 153270
rect 191840 153206 191892 153212
rect 191746 149152 191802 149161
rect 191746 149087 191802 149096
rect 190368 148436 190420 148442
rect 190368 148378 190420 148384
rect 189814 136776 189870 136785
rect 189814 136711 189870 136720
rect 189828 131102 189856 136711
rect 190380 132494 190408 148378
rect 191654 145888 191710 145897
rect 191654 145823 191710 145832
rect 191668 145625 191696 145823
rect 191654 145616 191710 145625
rect 191654 145551 191710 145560
rect 191102 144256 191158 144265
rect 191102 144191 191158 144200
rect 191116 137873 191144 144191
rect 191102 137864 191158 137873
rect 191102 137799 191158 137808
rect 190458 134736 190514 134745
rect 190458 134671 190514 134680
rect 190288 132466 190408 132494
rect 189816 131096 189868 131102
rect 189816 131038 189868 131044
rect 190288 125769 190316 132466
rect 190472 131850 190500 134671
rect 190460 131844 190512 131850
rect 190460 131786 190512 131792
rect 190366 129840 190422 129849
rect 190366 129775 190422 129784
rect 190274 125760 190330 125769
rect 190274 125695 190330 125704
rect 190380 125594 190408 129775
rect 190368 125588 190420 125594
rect 190368 125530 190420 125536
rect 191012 121440 191064 121446
rect 191012 121382 191064 121388
rect 191024 120329 191052 121382
rect 191010 120320 191066 120329
rect 191010 120255 191066 120264
rect 191116 117609 191144 137799
rect 191564 136604 191616 136610
rect 191564 136546 191616 136552
rect 191576 136377 191604 136546
rect 191562 136368 191618 136377
rect 191562 136303 191618 136312
rect 191562 135552 191618 135561
rect 191562 135487 191618 135496
rect 191576 135318 191604 135487
rect 191564 135312 191616 135318
rect 191564 135254 191616 135260
rect 191196 134904 191248 134910
rect 191196 134846 191248 134852
rect 191208 133929 191236 134846
rect 191194 133920 191250 133929
rect 191194 133855 191250 133864
rect 191668 128489 191696 145551
rect 191760 129742 191788 149087
rect 192496 148374 192524 153818
rect 192588 151814 192616 157270
rect 192588 151786 192892 151814
rect 192484 148368 192536 148374
rect 192484 148310 192536 148316
rect 191748 129736 191800 129742
rect 191748 129678 191800 129684
rect 191760 129305 191788 129678
rect 191746 129296 191802 129305
rect 191746 129231 191802 129240
rect 191654 128480 191710 128489
rect 191654 128415 191710 128424
rect 191746 127664 191802 127673
rect 191746 127599 191802 127608
rect 191760 127022 191788 127599
rect 191748 127016 191800 127022
rect 191748 126958 191800 126964
rect 191562 126576 191618 126585
rect 191562 126511 191618 126520
rect 191576 126274 191604 126511
rect 191564 126268 191616 126274
rect 191564 126210 191616 126216
rect 192496 124953 192524 148310
rect 192864 139913 192892 151786
rect 193036 149048 193088 149054
rect 193036 148990 193088 148996
rect 193048 147937 193076 148990
rect 193034 147928 193090 147937
rect 193034 147863 193090 147872
rect 192942 146976 192998 146985
rect 192942 146911 192998 146920
rect 192850 139904 192906 139913
rect 192850 139839 192906 139848
rect 192482 124944 192538 124953
rect 192482 124879 192538 124888
rect 191748 124092 191800 124098
rect 191748 124034 191800 124040
rect 191760 123049 191788 124034
rect 192956 123865 192984 146911
rect 193036 140548 193088 140554
rect 193036 140490 193088 140496
rect 193048 138281 193076 140490
rect 193034 138272 193090 138281
rect 193034 138207 193090 138216
rect 192942 123856 192998 123865
rect 192942 123791 192998 123800
rect 191746 123040 191802 123049
rect 191746 122975 191802 122984
rect 191746 122224 191802 122233
rect 191746 122159 191802 122168
rect 191760 121650 191788 122159
rect 191748 121644 191800 121650
rect 191748 121586 191800 121592
rect 191194 121408 191250 121417
rect 191194 121343 191196 121352
rect 191248 121343 191250 121352
rect 191196 121314 191248 121320
rect 191748 120080 191800 120086
rect 191748 120022 191800 120028
rect 191760 119513 191788 120022
rect 191746 119504 191802 119513
rect 191746 119439 191802 119448
rect 191746 118688 191802 118697
rect 191746 118623 191802 118632
rect 191760 117978 191788 118623
rect 191748 117972 191800 117978
rect 191748 117914 191800 117920
rect 191102 117600 191158 117609
rect 191102 117535 191158 117544
rect 191562 116784 191618 116793
rect 191562 116719 191618 116728
rect 189814 116512 189870 116521
rect 189814 116447 189870 116456
rect 189722 115968 189778 115977
rect 189722 115903 189778 115912
rect 189724 111852 189776 111858
rect 189724 111794 189776 111800
rect 188436 111104 188488 111110
rect 188436 111046 188488 111052
rect 189078 110800 189134 110809
rect 189078 110735 189134 110744
rect 189092 109002 189120 110735
rect 189080 108996 189132 109002
rect 189080 108938 189132 108944
rect 188434 107808 188490 107817
rect 188434 107743 188490 107752
rect 188448 78577 188476 107743
rect 188528 102196 188580 102202
rect 188528 102138 188580 102144
rect 188540 80034 188568 102138
rect 188804 98048 188856 98054
rect 188804 97990 188856 97996
rect 188816 93129 188844 97990
rect 189078 93256 189134 93265
rect 189078 93191 189134 93200
rect 188802 93120 188858 93129
rect 188802 93055 188858 93064
rect 189092 92585 189120 93191
rect 189078 92576 189134 92585
rect 189078 92511 189134 92520
rect 189736 89457 189764 111794
rect 189828 99657 189856 116447
rect 191576 116142 191604 116719
rect 191564 116136 191616 116142
rect 191564 116078 191616 116084
rect 191760 115954 191788 117914
rect 191576 115926 191788 115954
rect 190368 110492 190420 110498
rect 190368 110434 190420 110440
rect 189814 99648 189870 99657
rect 189814 99583 189870 99592
rect 190182 99512 190238 99521
rect 190182 99447 190238 99456
rect 189722 89448 189778 89457
rect 189722 89383 189778 89392
rect 188528 80028 188580 80034
rect 188528 79970 188580 79976
rect 188434 78568 188490 78577
rect 188434 78503 188490 78512
rect 188342 73128 188398 73137
rect 188342 73063 188398 73072
rect 187608 71052 187660 71058
rect 187608 70994 187660 71000
rect 186962 70272 187018 70281
rect 186962 70207 187018 70216
rect 188448 46918 188476 78503
rect 190196 75206 190224 99447
rect 190274 92576 190330 92585
rect 190274 92511 190330 92520
rect 190184 75200 190236 75206
rect 190184 75142 190236 75148
rect 190196 73166 190224 75142
rect 190184 73160 190236 73166
rect 190184 73102 190236 73108
rect 190288 66910 190316 92511
rect 190380 78674 190408 110434
rect 190644 110424 190696 110430
rect 190644 110366 190696 110372
rect 190656 109721 190684 110366
rect 190642 109712 190698 109721
rect 190642 109647 190698 109656
rect 190828 107636 190880 107642
rect 190828 107578 190880 107584
rect 190840 107001 190868 107578
rect 190826 106992 190882 107001
rect 190826 106927 190882 106936
rect 191196 106276 191248 106282
rect 191196 106218 191248 106224
rect 191208 106185 191236 106218
rect 191194 106176 191250 106185
rect 191194 106111 191250 106120
rect 191010 103456 191066 103465
rect 191010 103391 191066 103400
rect 191024 102202 191052 103391
rect 191012 102196 191064 102202
rect 191012 102138 191064 102144
rect 191102 93664 191158 93673
rect 191102 93599 191158 93608
rect 191116 92585 191144 93599
rect 191102 92576 191158 92585
rect 191102 92511 191158 92520
rect 191576 79354 191604 115926
rect 191748 115660 191800 115666
rect 191748 115602 191800 115608
rect 191760 115161 191788 115602
rect 191746 115152 191802 115161
rect 191746 115087 191802 115096
rect 191748 114504 191800 114510
rect 191748 114446 191800 114452
rect 191760 113257 191788 114446
rect 191838 114064 191894 114073
rect 191838 113999 191894 114008
rect 191746 113248 191802 113257
rect 191746 113183 191802 113192
rect 191748 112464 191800 112470
rect 191746 112432 191748 112441
rect 191800 112432 191802 112441
rect 191746 112367 191802 112376
rect 191748 111784 191800 111790
rect 191748 111726 191800 111732
rect 191760 110537 191788 111726
rect 191746 110528 191802 110537
rect 191852 110498 191880 113999
rect 191746 110463 191802 110472
rect 191840 110492 191892 110498
rect 191840 110434 191892 110440
rect 191748 108928 191800 108934
rect 191746 108896 191748 108905
rect 191800 108896 191802 108905
rect 191746 108831 191802 108840
rect 191748 105596 191800 105602
rect 191748 105538 191800 105544
rect 191760 105097 191788 105538
rect 191746 105088 191802 105097
rect 191746 105023 191802 105032
rect 191746 101552 191802 101561
rect 191746 101487 191802 101496
rect 191760 100774 191788 101487
rect 191748 100768 191800 100774
rect 191654 100736 191710 100745
rect 191748 100710 191800 100716
rect 191654 100671 191710 100680
rect 191668 99521 191696 100671
rect 191654 99512 191710 99521
rect 191654 99447 191710 99456
rect 191748 98116 191800 98122
rect 191748 98058 191800 98064
rect 191760 98025 191788 98058
rect 191746 98016 191802 98025
rect 191656 97980 191708 97986
rect 191746 97951 191802 97960
rect 191656 97922 191708 97928
rect 191668 97209 191696 97922
rect 191654 97200 191710 97209
rect 191654 97135 191710 97144
rect 191932 95940 191984 95946
rect 191932 95882 191984 95888
rect 191654 95840 191710 95849
rect 191654 95775 191710 95784
rect 191564 79348 191616 79354
rect 191564 79290 191616 79296
rect 190368 78668 190420 78674
rect 190368 78610 190420 78616
rect 190276 66904 190328 66910
rect 190276 66846 190328 66852
rect 188436 46912 188488 46918
rect 188436 46854 188488 46860
rect 186136 43444 186188 43450
rect 186136 43386 186188 43392
rect 184756 42084 184808 42090
rect 184756 42026 184808 42032
rect 191668 26926 191696 95775
rect 191840 94512 191892 94518
rect 191746 94480 191802 94489
rect 191840 94454 191892 94460
rect 191746 94415 191802 94424
rect 191656 26920 191708 26926
rect 191656 26862 191708 26868
rect 184204 8968 184256 8974
rect 184204 8910 184256 8916
rect 191760 6186 191788 94415
rect 191852 92478 191880 94454
rect 191944 92546 191972 95882
rect 192024 93900 192076 93906
rect 192024 93842 192076 93848
rect 191932 92540 191984 92546
rect 191932 92482 191984 92488
rect 191840 92472 191892 92478
rect 191840 92414 191892 92420
rect 192036 89622 192064 93842
rect 192024 89616 192076 89622
rect 192024 89558 192076 89564
rect 193048 83502 193076 138207
rect 193140 102649 193168 162007
rect 193232 148442 193260 260170
rect 193680 244996 193732 245002
rect 193680 244938 193732 244944
rect 193692 244882 193720 244938
rect 193692 244854 193812 244882
rect 193678 242856 193734 242865
rect 193678 242791 193734 242800
rect 193588 242276 193640 242282
rect 193588 242218 193640 242224
rect 193310 240136 193366 240145
rect 193310 240071 193366 240080
rect 193324 189786 193352 240071
rect 193600 238754 193628 242218
rect 193692 241534 193720 242791
rect 193680 241528 193732 241534
rect 193680 241470 193732 241476
rect 193600 238726 193720 238754
rect 193692 237386 193720 238726
rect 193784 238542 193812 244854
rect 252376 242344 252428 242350
rect 252376 242286 252428 242292
rect 198004 242072 198056 242078
rect 198096 242072 198148 242078
rect 198004 242014 198056 242020
rect 198094 242040 198096 242049
rect 242992 242072 243044 242078
rect 198148 242040 198150 242049
rect 194810 241590 195376 241618
rect 195348 240038 195376 241590
rect 195336 240032 195388 240038
rect 195336 239974 195388 239980
rect 193772 238536 193824 238542
rect 193772 238478 193824 238484
rect 193680 237380 193732 237386
rect 193680 237322 193732 237328
rect 194600 224256 194652 224262
rect 194600 224198 194652 224204
rect 193312 189780 193364 189786
rect 193312 189722 193364 189728
rect 193862 174584 193918 174593
rect 193862 174519 193918 174528
rect 193876 153785 193904 174519
rect 193862 153776 193918 153785
rect 193862 153711 193918 153720
rect 193220 148436 193272 148442
rect 193220 148378 193272 148384
rect 193588 144424 193640 144430
rect 193588 144366 193640 144372
rect 193600 140964 193628 144366
rect 194140 144288 194192 144294
rect 194140 144230 194192 144236
rect 194152 140964 194180 144230
rect 194612 142497 194640 224198
rect 195244 198008 195296 198014
rect 195244 197950 195296 197956
rect 194876 170672 194928 170678
rect 194876 170614 194928 170620
rect 194888 170406 194916 170614
rect 194876 170400 194928 170406
rect 194876 170342 194928 170348
rect 194598 142488 194654 142497
rect 194598 142423 194654 142432
rect 194612 142154 194640 142423
rect 194612 142126 194732 142154
rect 193218 140856 193274 140865
rect 193218 140791 193274 140800
rect 193232 137970 193260 140791
rect 194704 140434 194732 142126
rect 194888 140554 194916 170342
rect 195256 141137 195284 197950
rect 195348 186998 195376 239974
rect 196070 238096 196126 238105
rect 196070 238031 196126 238040
rect 195978 225584 196034 225593
rect 195978 225519 196034 225528
rect 195992 221474 196020 225519
rect 195980 221468 196032 221474
rect 195980 221410 196032 221416
rect 195336 186992 195388 186998
rect 195336 186934 195388 186940
rect 195336 184204 195388 184210
rect 195336 184146 195388 184152
rect 195348 170678 195376 184146
rect 196084 175234 196112 238031
rect 196624 237312 196676 237318
rect 196624 237254 196676 237260
rect 196636 236774 196664 237254
rect 197188 236774 197216 241604
rect 196624 236768 196676 236774
rect 196624 236710 196676 236716
rect 197176 236768 197228 236774
rect 197176 236710 197228 236716
rect 196636 215937 196664 236710
rect 197360 236700 197412 236706
rect 197360 236642 197412 236648
rect 197372 234433 197400 236642
rect 197358 234424 197414 234433
rect 197358 234359 197414 234368
rect 196622 215928 196678 215937
rect 196622 215863 196678 215872
rect 196624 195288 196676 195294
rect 196624 195230 196676 195236
rect 196072 175228 196124 175234
rect 196072 175170 196124 175176
rect 195336 170672 195388 170678
rect 195336 170614 195388 170620
rect 196636 167074 196664 195230
rect 197358 193896 197414 193905
rect 197358 193831 197414 193840
rect 196808 175228 196860 175234
rect 196808 175170 196860 175176
rect 196820 173942 196848 175170
rect 196808 173936 196860 173942
rect 196808 173878 196860 173884
rect 196716 170400 196768 170406
rect 196716 170342 196768 170348
rect 195980 167068 196032 167074
rect 195980 167010 196032 167016
rect 196624 167068 196676 167074
rect 196624 167010 196676 167016
rect 195428 143540 195480 143546
rect 195428 143482 195480 143488
rect 195242 141128 195298 141137
rect 195242 141063 195298 141072
rect 195440 140964 195468 143482
rect 195992 140964 196020 167010
rect 196530 146432 196586 146441
rect 196530 146367 196586 146376
rect 196544 140964 196572 146367
rect 196728 142361 196756 170342
rect 196820 169017 196848 173878
rect 196806 169008 196862 169017
rect 196806 168943 196862 168952
rect 196714 142352 196770 142361
rect 196714 142287 196770 142296
rect 196728 140978 196756 142287
rect 197372 140978 197400 193831
rect 198016 178702 198044 242014
rect 198094 241975 198150 241984
rect 242990 242040 242992 242049
rect 243044 242040 243046 242049
rect 250166 242040 250222 242049
rect 242990 241975 243046 241984
rect 249812 241998 250166 242026
rect 199594 241590 200068 241618
rect 200040 196654 200068 241590
rect 201972 238406 202000 241604
rect 201500 238400 201552 238406
rect 201500 238342 201552 238348
rect 201960 238400 202012 238406
rect 201960 238342 202012 238348
rect 200028 196648 200080 196654
rect 200028 196590 200080 196596
rect 198924 179784 198976 179790
rect 198924 179726 198976 179732
rect 198004 178696 198056 178702
rect 198004 178638 198056 178644
rect 198740 159248 198792 159254
rect 198740 159190 198792 159196
rect 198752 158846 198780 159190
rect 198740 158840 198792 158846
rect 198740 158782 198792 158788
rect 198752 149818 198780 158782
rect 198936 151814 198964 179726
rect 200672 168496 200724 168502
rect 200672 168438 200724 168444
rect 200684 166977 200712 168438
rect 200118 166968 200174 166977
rect 200118 166903 200174 166912
rect 200670 166968 200726 166977
rect 200670 166903 200726 166912
rect 199384 164892 199436 164898
rect 199384 164834 199436 164840
rect 199396 159254 199424 164834
rect 199384 159248 199436 159254
rect 199384 159190 199436 159196
rect 198936 151786 199056 151814
rect 198752 149790 198964 149818
rect 198830 149696 198886 149705
rect 198830 149631 198886 149640
rect 198372 144968 198424 144974
rect 198372 144910 198424 144916
rect 197910 144800 197966 144809
rect 197910 144735 197966 144744
rect 197924 143546 197952 144735
rect 197912 143540 197964 143546
rect 197912 143482 197964 143488
rect 196728 140950 197110 140978
rect 197372 140950 197846 140978
rect 198384 140964 198412 144910
rect 198844 140978 198872 149631
rect 198936 141386 198964 149790
rect 199028 142934 199056 151786
rect 200132 144022 200160 166903
rect 200210 157992 200266 158001
rect 200210 157927 200266 157936
rect 200120 144016 200172 144022
rect 200120 143958 200172 143964
rect 199016 142928 199068 142934
rect 199016 142870 199068 142876
rect 198936 141358 199240 141386
rect 199212 140978 199240 141358
rect 198844 140950 198950 140978
rect 199212 140950 199686 140978
rect 200224 140964 200252 157927
rect 201512 151162 201540 238342
rect 204168 225004 204220 225010
rect 204168 224946 204220 224952
rect 204180 222154 204208 224946
rect 204364 224942 204392 241604
rect 205640 234524 205692 234530
rect 205640 234466 205692 234472
rect 205652 234122 205680 234466
rect 206756 234122 206784 241604
rect 207662 241088 207718 241097
rect 207662 241023 207718 241032
rect 207296 240780 207348 240786
rect 207296 240722 207348 240728
rect 205640 234116 205692 234122
rect 205640 234058 205692 234064
rect 206744 234116 206796 234122
rect 206744 234058 206796 234064
rect 204902 226944 204958 226953
rect 204902 226879 204958 226888
rect 204352 224936 204404 224942
rect 204352 224878 204404 224884
rect 204168 222148 204220 222154
rect 204168 222090 204220 222096
rect 203524 203584 203576 203590
rect 203524 203526 203576 203532
rect 203536 167686 203564 203526
rect 204720 169788 204772 169794
rect 204720 169730 204772 169736
rect 204732 168502 204760 169730
rect 204260 168496 204312 168502
rect 204260 168438 204312 168444
rect 204720 168496 204772 168502
rect 204720 168438 204772 168444
rect 202880 167680 202932 167686
rect 202880 167622 202932 167628
rect 203524 167680 203576 167686
rect 203524 167622 203576 167628
rect 202788 159384 202840 159390
rect 202788 159326 202840 159332
rect 202800 155990 202828 159326
rect 201684 155984 201736 155990
rect 201684 155926 201736 155932
rect 202788 155984 202840 155990
rect 202788 155926 202840 155932
rect 201696 151814 201724 155926
rect 201696 151786 202184 151814
rect 201500 151156 201552 151162
rect 201500 151098 201552 151104
rect 201592 151088 201644 151094
rect 201592 151030 201644 151036
rect 201314 144120 201370 144129
rect 201314 144055 201370 144064
rect 200396 144016 200448 144022
rect 200396 143958 200448 143964
rect 200408 140978 200436 143958
rect 200408 140950 200790 140978
rect 201328 140964 201356 144055
rect 201604 140978 201632 151030
rect 202156 140978 202184 151786
rect 202892 142225 202920 167622
rect 204168 150476 204220 150482
rect 204168 150418 204220 150424
rect 204180 149802 204208 150418
rect 204168 149796 204220 149802
rect 204168 149738 204220 149744
rect 204272 144022 204300 168438
rect 204350 152008 204406 152017
rect 204350 151943 204406 151952
rect 204364 147674 204392 151943
rect 204364 147646 204484 147674
rect 204260 144016 204312 144022
rect 204260 143958 204312 143964
rect 202878 142216 202934 142225
rect 202878 142151 202934 142160
rect 203890 142216 203946 142225
rect 203890 142151 203946 142160
rect 203156 141432 203208 141438
rect 203156 141374 203208 141380
rect 203168 140978 203196 141374
rect 201604 140950 202078 140978
rect 202156 140950 202630 140978
rect 203168 140964 203472 140978
rect 203904 140964 203932 142151
rect 204456 140964 204484 147646
rect 204916 145761 204944 226879
rect 205652 170406 205680 234058
rect 207308 233238 207336 240722
rect 207676 234530 207704 241023
rect 207664 234524 207716 234530
rect 207664 234466 207716 234472
rect 207296 233232 207348 233238
rect 207296 233174 207348 233180
rect 207018 232520 207074 232529
rect 207018 232455 207074 232464
rect 207032 229129 207060 232455
rect 207018 229120 207074 229129
rect 207018 229055 207074 229064
rect 206284 224256 206336 224262
rect 206284 224198 206336 224204
rect 206296 174758 206324 224198
rect 205732 174752 205784 174758
rect 205732 174694 205784 174700
rect 206284 174752 206336 174758
rect 206284 174694 206336 174700
rect 205744 174554 205772 174694
rect 205732 174548 205784 174554
rect 205732 174490 205784 174496
rect 205744 172582 205772 174490
rect 205732 172576 205784 172582
rect 205732 172518 205784 172524
rect 205640 170400 205692 170406
rect 205640 170342 205692 170348
rect 204996 165640 205048 165646
rect 204996 165582 205048 165588
rect 205008 153785 205036 165582
rect 204994 153776 205050 153785
rect 204994 153711 205050 153720
rect 205744 151814 205772 172518
rect 207676 156233 207704 234466
rect 209148 231810 209176 241604
rect 211540 240106 211568 241604
rect 212446 240952 212502 240961
rect 212446 240887 212502 240896
rect 211528 240100 211580 240106
rect 211528 240042 211580 240048
rect 210422 236600 210478 236609
rect 210422 236535 210478 236544
rect 209136 231804 209188 231810
rect 209136 231746 209188 231752
rect 210436 227633 210464 236535
rect 210514 229120 210570 229129
rect 210514 229055 210570 229064
rect 210422 227624 210478 227633
rect 210422 227559 210478 227568
rect 209044 227112 209096 227118
rect 209044 227054 209096 227060
rect 207756 180124 207808 180130
rect 207756 180066 207808 180072
rect 207662 156224 207718 156233
rect 207662 156159 207718 156168
rect 205744 151786 205864 151814
rect 204902 145752 204958 145761
rect 204902 145687 204958 145696
rect 204916 145586 204944 145687
rect 204904 145580 204956 145586
rect 204904 145522 204956 145528
rect 204628 144016 204680 144022
rect 204628 143958 204680 143964
rect 204640 140978 204668 143958
rect 205836 140978 205864 151786
rect 206376 149796 206428 149802
rect 206376 149738 206428 149744
rect 203182 140950 203472 140964
rect 204640 140950 205022 140978
rect 205836 140950 206310 140978
rect 203444 140826 203472 140950
rect 205640 140888 205692 140894
rect 205574 140836 205640 140842
rect 205574 140830 205692 140836
rect 206388 140842 206416 149738
rect 207018 148064 207074 148073
rect 207018 147999 207074 148008
rect 207032 140978 207060 147999
rect 207676 141545 207704 156159
rect 207768 149705 207796 180066
rect 208400 164280 208452 164286
rect 208400 164222 208452 164228
rect 208412 162761 208440 164222
rect 208398 162752 208454 162761
rect 208398 162687 208454 162696
rect 207848 151088 207900 151094
rect 207848 151030 207900 151036
rect 207754 149696 207810 149705
rect 207754 149631 207810 149640
rect 207662 141536 207718 141545
rect 207662 141471 207718 141480
rect 207860 141409 207888 151030
rect 208412 147014 208440 162687
rect 208490 152416 208546 152425
rect 208490 152351 208546 152360
rect 208504 151910 208532 152351
rect 208492 151904 208544 151910
rect 208492 151846 208544 151852
rect 208400 147008 208452 147014
rect 208400 146950 208452 146956
rect 207846 141400 207902 141409
rect 207846 141335 207902 141344
rect 208122 141400 208178 141409
rect 208122 141335 208178 141344
rect 207032 140950 207414 140978
rect 208136 140964 208164 141335
rect 208504 140978 208532 151846
rect 208504 140950 208702 140978
rect 206558 140856 206614 140865
rect 205574 140828 205680 140830
rect 203432 140820 203484 140826
rect 203432 140762 203484 140768
rect 205560 140814 205680 140828
rect 206388 140814 206558 140842
rect 194876 140548 194928 140554
rect 194876 140490 194928 140496
rect 205180 140480 205232 140486
rect 194966 140448 195022 140457
rect 194704 140420 194966 140434
rect 194718 140406 194966 140420
rect 205560 140434 205588 140814
rect 206614 140814 206862 140842
rect 206558 140791 206614 140800
rect 209056 140593 209084 227054
rect 210436 226409 210464 227559
rect 210422 226400 210478 226409
rect 210422 226335 210478 226344
rect 210528 226234 210556 229055
rect 211066 226400 211122 226409
rect 211066 226335 211122 226344
rect 210516 226228 210568 226234
rect 210516 226170 210568 226176
rect 210528 225010 210556 226170
rect 210516 225004 210568 225010
rect 210516 224946 210568 224952
rect 210976 225004 211028 225010
rect 210976 224946 211028 224952
rect 209136 202224 209188 202230
rect 209136 202166 209188 202172
rect 209148 171737 209176 202166
rect 210422 175400 210478 175409
rect 210422 175335 210478 175344
rect 209134 171728 209190 171737
rect 209134 171663 209190 171672
rect 210436 155961 210464 175335
rect 210988 156058 211016 224946
rect 210516 156052 210568 156058
rect 210516 155994 210568 156000
rect 210976 156052 211028 156058
rect 210976 155994 211028 156000
rect 210422 155952 210478 155961
rect 210422 155887 210478 155896
rect 210436 151814 210464 155887
rect 210528 155417 210556 155994
rect 210514 155408 210570 155417
rect 210514 155343 210570 155352
rect 210436 151786 210648 151814
rect 209136 147008 209188 147014
rect 209136 146950 209188 146956
rect 209148 140978 209176 146950
rect 209872 145036 209924 145042
rect 209872 144978 209924 144984
rect 209148 140950 209254 140978
rect 209042 140584 209098 140593
rect 209884 140570 209912 144978
rect 210514 144120 210570 144129
rect 210514 144055 210570 144064
rect 210528 140964 210556 144055
rect 210620 140978 210648 151786
rect 211080 149054 211108 226335
rect 211802 192536 211858 192545
rect 211802 192471 211858 192480
rect 211158 153776 211214 153785
rect 211158 153711 211214 153720
rect 211068 149048 211120 149054
rect 211068 148990 211120 148996
rect 211080 148481 211108 148990
rect 211066 148472 211122 148481
rect 211066 148407 211122 148416
rect 211172 140978 211200 153711
rect 211816 152017 211844 192471
rect 212460 158817 212488 240887
rect 213184 240100 213236 240106
rect 213184 240042 213236 240048
rect 213196 216753 213224 240042
rect 213932 237386 213960 241604
rect 216324 241534 216352 241604
rect 215300 241528 215352 241534
rect 215300 241470 215352 241476
rect 216312 241528 216364 241534
rect 216312 241470 216364 241476
rect 213920 237380 213972 237386
rect 213920 237322 213972 237328
rect 213932 236026 213960 237322
rect 214656 236768 214708 236774
rect 214656 236710 214708 236716
rect 213920 236020 213972 236026
rect 213920 235962 213972 235968
rect 214564 236020 214616 236026
rect 214564 235962 214616 235968
rect 213182 216744 213238 216753
rect 213182 216679 213238 216688
rect 213184 189780 213236 189786
rect 213184 189722 213236 189728
rect 213196 177342 213224 189722
rect 214576 180198 214604 235962
rect 214668 229090 214696 236710
rect 214656 229084 214708 229090
rect 214656 229026 214708 229032
rect 214654 200696 214710 200705
rect 214654 200631 214710 200640
rect 214564 180192 214616 180198
rect 214564 180134 214616 180140
rect 213184 177336 213236 177342
rect 213184 177278 213236 177284
rect 211894 158808 211950 158817
rect 211894 158743 211950 158752
rect 212446 158808 212502 158817
rect 212446 158743 212502 158752
rect 211802 152008 211858 152017
rect 211802 151943 211858 151952
rect 211908 151065 211936 158743
rect 213196 151814 213224 177278
rect 214012 175976 214064 175982
rect 214012 175918 214064 175924
rect 214024 175302 214052 175918
rect 214012 175296 214064 175302
rect 214012 175238 214064 175244
rect 213012 151786 213224 151814
rect 214024 151814 214052 175238
rect 214668 157350 214696 200631
rect 214656 157344 214708 157350
rect 214656 157286 214708 157292
rect 214024 151786 214328 151814
rect 211894 151056 211950 151065
rect 211894 150991 211950 151000
rect 213012 147694 213040 151786
rect 213000 147688 213052 147694
rect 213000 147630 213052 147636
rect 212908 142860 212960 142866
rect 212908 142802 212960 142808
rect 212354 142488 212410 142497
rect 212354 142423 212410 142432
rect 210620 140950 211094 140978
rect 211172 140950 211646 140978
rect 212368 140964 212396 142423
rect 210148 140616 210200 140622
rect 210146 140584 210148 140593
rect 210200 140584 210202 140593
rect 209806 140554 210096 140570
rect 209806 140548 210108 140554
rect 209806 140542 210056 140548
rect 209042 140519 209098 140528
rect 210146 140519 210202 140528
rect 210056 140490 210108 140496
rect 205232 140428 205588 140434
rect 205180 140422 205588 140428
rect 212540 140480 212592 140486
rect 212920 140434 212948 142802
rect 213012 140978 213040 147630
rect 214012 147620 214064 147626
rect 214012 147562 214064 147568
rect 213012 140950 213486 140978
rect 214024 140964 214052 147562
rect 214300 140978 214328 151786
rect 215312 148345 215340 241470
rect 217322 231160 217378 231169
rect 217322 231095 217378 231104
rect 217336 217977 217364 231095
rect 217322 217968 217378 217977
rect 217322 217903 217378 217912
rect 217336 172553 217364 217903
rect 217322 172544 217378 172553
rect 217322 172479 217378 172488
rect 215392 170400 215444 170406
rect 215392 170342 215444 170348
rect 215404 161498 215432 170342
rect 216678 169008 216734 169017
rect 216678 168943 216734 168952
rect 215392 161492 215444 161498
rect 215392 161434 215444 161440
rect 215404 151814 215432 161434
rect 216692 151814 216720 168943
rect 215404 151786 216168 151814
rect 216692 151786 216996 151814
rect 215298 148336 215354 148345
rect 215298 148271 215354 148280
rect 215850 143712 215906 143721
rect 215850 143647 215906 143656
rect 214300 140950 214774 140978
rect 215864 140964 215892 143647
rect 216140 140978 216168 151786
rect 216772 149728 216824 149734
rect 216772 149670 216824 149676
rect 216784 140978 216812 149670
rect 216864 149116 216916 149122
rect 216864 149058 216916 149064
rect 216876 147626 216904 149058
rect 216864 147620 216916 147626
rect 216864 147562 216916 147568
rect 216968 142154 216996 151786
rect 217336 149122 217364 172479
rect 218716 171134 218744 241604
rect 221108 237726 221136 241604
rect 222108 238672 222160 238678
rect 222108 238614 222160 238620
rect 222120 237726 222148 238614
rect 221096 237720 221148 237726
rect 221096 237662 221148 237668
rect 222108 237720 222160 237726
rect 222108 237662 222160 237668
rect 219440 229764 219492 229770
rect 219440 229706 219492 229712
rect 218716 171106 218928 171134
rect 218796 160132 218848 160138
rect 218796 160074 218848 160080
rect 218060 155984 218112 155990
rect 218060 155926 218112 155932
rect 218072 153882 218100 155926
rect 218704 154624 218756 154630
rect 218704 154566 218756 154572
rect 218060 153876 218112 153882
rect 218060 153818 218112 153824
rect 217324 149116 217376 149122
rect 217324 149058 217376 149064
rect 218716 149054 218744 154566
rect 218520 149048 218572 149054
rect 218520 148990 218572 148996
rect 218704 149048 218756 149054
rect 218704 148990 218756 148996
rect 218244 142928 218296 142934
rect 218244 142870 218296 142876
rect 218256 142225 218284 142870
rect 218242 142216 218298 142225
rect 216968 142126 217364 142154
rect 218242 142151 218298 142160
rect 217336 140978 217364 142126
rect 216140 140950 216614 140978
rect 216784 140950 217166 140978
rect 217336 140950 217718 140978
rect 218256 140964 218284 142151
rect 218532 140978 218560 148990
rect 218808 146266 218836 160074
rect 218900 155990 218928 171106
rect 219452 167113 219480 229706
rect 220084 222896 220136 222902
rect 220084 222838 220136 222844
rect 220096 208321 220124 222838
rect 220082 208312 220138 208321
rect 220082 208247 220138 208256
rect 220084 176724 220136 176730
rect 220084 176666 220136 176672
rect 219438 167104 219494 167113
rect 219438 167039 219494 167048
rect 218888 155984 218940 155990
rect 218888 155926 218940 155932
rect 218796 146260 218848 146266
rect 218796 146202 218848 146208
rect 219532 143540 219584 143546
rect 219532 143482 219584 143488
rect 218532 140950 219006 140978
rect 219544 140964 219572 143482
rect 220096 142186 220124 176666
rect 221464 171828 221516 171834
rect 221464 171770 221516 171776
rect 220174 167104 220230 167113
rect 220174 167039 220230 167048
rect 220188 150521 220216 167039
rect 221004 158772 221056 158778
rect 221004 158714 221056 158720
rect 220820 151836 220872 151842
rect 220820 151778 220872 151784
rect 220832 151094 220860 151778
rect 220820 151088 220872 151094
rect 220820 151030 220872 151036
rect 220174 150512 220230 150521
rect 220174 150447 220230 150456
rect 220188 143546 220216 150447
rect 220176 143540 220228 143546
rect 220176 143482 220228 143488
rect 220084 142180 220136 142186
rect 220004 142128 220084 142154
rect 220004 142126 220136 142128
rect 220004 140978 220032 142126
rect 220084 142122 220136 142126
rect 221016 140978 221044 158714
rect 221476 146402 221504 171770
rect 222120 151842 222148 237662
rect 223500 229090 223528 241604
rect 225604 240168 225656 240174
rect 225604 240110 225656 240116
rect 224224 239420 224276 239426
rect 224224 239362 224276 239368
rect 223488 229084 223540 229090
rect 223488 229026 223540 229032
rect 223500 227798 223528 229026
rect 222936 227792 222988 227798
rect 222936 227734 222988 227740
rect 223488 227792 223540 227798
rect 223488 227734 223540 227740
rect 222844 220108 222896 220114
rect 222844 220050 222896 220056
rect 222384 212424 222436 212430
rect 222384 212366 222436 212372
rect 222200 168428 222252 168434
rect 222200 168370 222252 168376
rect 222108 151836 222160 151842
rect 222108 151778 222160 151784
rect 221464 146396 221516 146402
rect 221464 146338 221516 146344
rect 221096 146260 221148 146266
rect 221096 146202 221148 146208
rect 220004 140950 220110 140978
rect 220846 140950 221044 140978
rect 221108 140978 221136 146202
rect 221476 142154 221504 146338
rect 221476 142126 221596 142154
rect 221568 140978 221596 142126
rect 222212 141137 222240 168370
rect 222292 167680 222344 167686
rect 222292 167622 222344 167628
rect 222304 162926 222332 167622
rect 222292 162920 222344 162926
rect 222292 162862 222344 162868
rect 222198 141128 222254 141137
rect 222198 141063 222254 141072
rect 222304 140978 222332 162862
rect 222396 152522 222424 212366
rect 222856 168434 222884 220050
rect 222948 212430 222976 227734
rect 224236 217938 224264 239362
rect 224868 239012 224920 239018
rect 224868 238954 224920 238960
rect 224224 217932 224276 217938
rect 224224 217874 224276 217880
rect 222936 212424 222988 212430
rect 222936 212366 222988 212372
rect 222844 168428 222896 168434
rect 222844 168370 222896 168376
rect 224224 165708 224276 165714
rect 224224 165650 224276 165656
rect 223578 157448 223634 157457
rect 223578 157383 223634 157392
rect 222384 152516 222436 152522
rect 222384 152458 222436 152464
rect 222844 152516 222896 152522
rect 222844 152458 222896 152464
rect 222856 151978 222884 152458
rect 222844 151972 222896 151978
rect 222844 151914 222896 151920
rect 222856 144809 222884 151914
rect 222842 144800 222898 144809
rect 222842 144735 222898 144744
rect 222842 141536 222898 141545
rect 222842 141471 222898 141480
rect 221108 140950 221398 140978
rect 221568 140950 221950 140978
rect 222304 140950 222502 140978
rect 222856 140729 222884 141471
rect 223210 141128 223266 141137
rect 223210 141063 223266 141072
rect 223224 140842 223252 141063
rect 223592 140978 223620 157383
rect 223672 153944 223724 153950
rect 223672 153886 223724 153892
rect 223684 144090 223712 153886
rect 223672 144084 223724 144090
rect 223672 144026 223724 144032
rect 224236 142361 224264 165650
rect 224776 163532 224828 163538
rect 224776 163474 224828 163480
rect 224788 157457 224816 163474
rect 224774 157448 224830 157457
rect 224774 157383 224830 157392
rect 224498 144256 224554 144265
rect 224880 144226 224908 238954
rect 225616 231810 225644 240110
rect 225984 239018 226012 241604
rect 225972 239012 226024 239018
rect 225972 238954 226024 238960
rect 225604 231804 225656 231810
rect 225604 231746 225656 231752
rect 224960 180192 225012 180198
rect 224960 180134 225012 180140
rect 224972 154698 225000 180134
rect 224960 154692 225012 154698
rect 224960 154634 225012 154640
rect 224972 151814 225000 154634
rect 224972 151786 225092 151814
rect 224960 146328 225012 146334
rect 224960 146270 225012 146276
rect 224498 144191 224500 144200
rect 224552 144191 224554 144200
rect 224868 144220 224920 144226
rect 224500 144162 224552 144168
rect 224868 144162 224920 144168
rect 224500 144084 224552 144090
rect 224500 144026 224552 144032
rect 224222 142352 224278 142361
rect 224222 142287 224278 142296
rect 224236 142154 224264 142287
rect 224236 142126 224356 142154
rect 223592 140950 223790 140978
rect 224328 140964 224356 142126
rect 224512 140978 224540 144026
rect 224512 140950 224894 140978
rect 223394 140856 223450 140865
rect 223224 140828 223394 140842
rect 223238 140814 223394 140828
rect 223394 140791 223450 140800
rect 222842 140720 222898 140729
rect 222842 140655 222898 140664
rect 215390 140584 215446 140593
rect 215326 140542 215390 140570
rect 215390 140519 215446 140528
rect 215404 140486 215432 140519
rect 212592 140428 212948 140434
rect 212540 140422 212948 140428
rect 215392 140480 215444 140486
rect 215392 140422 215444 140428
rect 205192 140420 205588 140422
rect 212552 140420 212948 140422
rect 205192 140406 205574 140420
rect 212552 140406 212934 140420
rect 194966 140383 195022 140392
rect 193402 140176 193458 140185
rect 193402 140111 193404 140120
rect 193456 140111 193458 140120
rect 193404 140082 193456 140088
rect 193220 137964 193272 137970
rect 193220 137906 193272 137912
rect 193218 131880 193274 131889
rect 193218 131815 193274 131824
rect 193232 131481 193260 131815
rect 193218 131472 193274 131481
rect 193218 131407 193274 131416
rect 193232 104281 193260 131407
rect 224972 122834 225000 146270
rect 225064 129713 225092 151786
rect 225144 140480 225196 140486
rect 225144 140422 225196 140428
rect 225156 139466 225184 140422
rect 225144 139460 225196 139466
rect 225144 139402 225196 139408
rect 225050 129704 225106 129713
rect 225050 129639 225106 129648
rect 224972 122806 225092 122834
rect 225064 113801 225092 122806
rect 225142 114880 225198 114889
rect 225142 114815 225198 114824
rect 225050 113792 225106 113801
rect 225050 113727 225106 113736
rect 225050 109168 225106 109177
rect 224972 109126 225050 109154
rect 193218 104272 193274 104281
rect 193218 104207 193274 104216
rect 193126 102640 193182 102649
rect 193126 102575 193182 102584
rect 193126 92576 193182 92585
rect 193126 92511 193182 92520
rect 193036 83496 193088 83502
rect 193036 83438 193088 83444
rect 193140 76566 193168 92511
rect 193128 76560 193180 76566
rect 193128 76502 193180 76508
rect 193232 73817 193260 104207
rect 224040 93424 224092 93430
rect 199198 93392 199254 93401
rect 198950 93364 199198 93378
rect 198936 93350 199198 93364
rect 198936 92834 198964 93350
rect 208950 93392 209006 93401
rect 208702 93364 208950 93378
rect 199198 93327 199254 93336
rect 208688 93350 208950 93364
rect 208688 92834 208716 93350
rect 221950 93362 222148 93378
rect 224040 93366 224092 93372
rect 221950 93356 222160 93362
rect 221950 93350 222108 93356
rect 208950 93327 209006 93336
rect 222108 93298 222160 93304
rect 213274 93120 213330 93129
rect 213274 93055 213330 93064
rect 193324 92806 193614 92834
rect 193692 92806 194166 92834
rect 194718 92806 194824 92834
rect 193218 73808 193274 73817
rect 193218 73743 193274 73752
rect 193324 68950 193352 92806
rect 193692 84194 193720 92806
rect 194692 90976 194744 90982
rect 194692 90918 194744 90924
rect 194704 90574 194732 90918
rect 194692 90568 194744 90574
rect 194692 90510 194744 90516
rect 193416 84182 193720 84194
rect 193404 84176 193720 84182
rect 193456 84166 193720 84176
rect 193404 84118 193456 84124
rect 193416 83570 193444 84118
rect 193404 83564 193456 83570
rect 193404 83506 193456 83512
rect 193312 68944 193364 68950
rect 193312 68886 193364 68892
rect 193864 68944 193916 68950
rect 193864 68886 193916 68892
rect 193876 63510 193904 68886
rect 193864 63504 193916 63510
rect 193864 63446 193916 63452
rect 193876 28286 193904 63446
rect 194704 61946 194732 90510
rect 194796 62082 194824 92806
rect 195256 90574 195284 92820
rect 195992 91050 196020 92820
rect 196544 92449 196572 92820
rect 196530 92440 196586 92449
rect 196530 92375 196586 92384
rect 195980 91044 196032 91050
rect 195980 90986 196032 90992
rect 195244 90568 195296 90574
rect 195244 90510 195296 90516
rect 194784 62076 194836 62082
rect 194784 62018 194836 62024
rect 194692 61940 194744 61946
rect 194692 61882 194744 61888
rect 194704 60790 194732 61882
rect 194692 60784 194744 60790
rect 194692 60726 194744 60732
rect 194796 60722 194824 62018
rect 195244 60784 195296 60790
rect 195244 60726 195296 60732
rect 194784 60716 194836 60722
rect 194784 60658 194836 60664
rect 195256 33794 195284 60726
rect 195992 59294 196020 90986
rect 197096 86873 197124 92820
rect 197662 92806 198044 92834
rect 198752 92820 198964 92834
rect 198016 92449 198044 92806
rect 198002 92440 198058 92449
rect 198002 92375 198058 92384
rect 197082 86864 197138 86873
rect 197082 86799 197138 86808
rect 198016 66230 198044 92375
rect 198384 85474 198412 92820
rect 198752 92806 198950 92820
rect 199396 92806 199502 92834
rect 198372 85468 198424 85474
rect 198372 85410 198424 85416
rect 198004 66224 198056 66230
rect 198004 66166 198056 66172
rect 195980 59288 196032 59294
rect 195980 59230 196032 59236
rect 196624 59288 196676 59294
rect 196624 59230 196676 59236
rect 195244 33788 195296 33794
rect 195244 33730 195296 33736
rect 193864 28280 193916 28286
rect 193864 28222 193916 28228
rect 196636 8974 196664 59230
rect 198016 10334 198044 66166
rect 198752 58682 198780 92806
rect 199396 89622 199424 92806
rect 200224 91089 200252 92820
rect 200776 92177 200804 92820
rect 200868 92806 201342 92834
rect 201604 92806 201894 92834
rect 200762 92168 200818 92177
rect 200762 92103 200818 92112
rect 200210 91080 200266 91089
rect 200210 91015 200266 91024
rect 199384 89616 199436 89622
rect 199384 89558 199436 89564
rect 199396 60042 199424 89558
rect 200868 88482 200896 92806
rect 200946 91080 201002 91089
rect 200946 91015 201002 91024
rect 200132 88454 200896 88482
rect 200132 82754 200160 88454
rect 200960 84194 200988 91015
rect 200776 84166 200988 84194
rect 200120 82748 200172 82754
rect 200120 82690 200172 82696
rect 200776 66230 200804 84166
rect 201408 82748 201460 82754
rect 201408 82690 201460 82696
rect 201420 82142 201448 82690
rect 201408 82136 201460 82142
rect 201408 82078 201460 82084
rect 201604 80714 201632 92806
rect 202616 92410 202644 92820
rect 202892 92806 203182 92834
rect 202604 92404 202656 92410
rect 202604 92346 202656 92352
rect 201592 80708 201644 80714
rect 201592 80650 201644 80656
rect 201604 80102 201632 80650
rect 201592 80096 201644 80102
rect 201592 80038 201644 80044
rect 202144 80096 202196 80102
rect 202144 80038 202196 80044
rect 200764 66224 200816 66230
rect 200764 66166 200816 66172
rect 201408 66224 201460 66230
rect 201408 66166 201460 66172
rect 199384 60036 199436 60042
rect 199384 59978 199436 59984
rect 198740 58676 198792 58682
rect 198740 58618 198792 58624
rect 201420 13122 201448 66166
rect 202156 56574 202184 80038
rect 202892 77897 202920 92806
rect 203720 90545 203748 92820
rect 203706 90536 203762 90545
rect 203706 90471 203762 90480
rect 203720 88097 203748 90471
rect 204456 90409 204484 92820
rect 204442 90400 204498 90409
rect 204442 90335 204498 90344
rect 204456 89622 204484 90335
rect 204444 89616 204496 89622
rect 204444 89558 204496 89564
rect 203706 88088 203762 88097
rect 203706 88023 203762 88032
rect 205008 85542 205036 92820
rect 205560 92177 205588 92820
rect 206112 92449 206140 92820
rect 206098 92440 206154 92449
rect 206098 92375 206154 92384
rect 205546 92168 205602 92177
rect 205546 92103 205602 92112
rect 205560 88262 205588 92103
rect 206848 90273 206876 92820
rect 207400 92546 207428 92820
rect 207492 92806 207966 92834
rect 208412 92820 208716 92834
rect 208412 92806 208702 92820
rect 207388 92540 207440 92546
rect 207388 92482 207440 92488
rect 205638 90264 205694 90273
rect 205638 90199 205694 90208
rect 206834 90264 206890 90273
rect 206834 90199 206890 90208
rect 205548 88256 205600 88262
rect 205548 88198 205600 88204
rect 204996 85536 205048 85542
rect 204996 85478 205048 85484
rect 202878 77888 202934 77897
rect 202878 77823 202934 77832
rect 203522 77888 203578 77897
rect 203522 77823 203578 77832
rect 203536 77217 203564 77823
rect 203522 77208 203578 77217
rect 203522 77143 203578 77152
rect 205652 64802 205680 90199
rect 205732 89616 205784 89622
rect 205732 89558 205784 89564
rect 205744 86902 205772 89558
rect 207400 87650 207428 92482
rect 207388 87644 207440 87650
rect 207388 87586 207440 87592
rect 205732 86896 205784 86902
rect 205732 86838 205784 86844
rect 207492 84194 207520 92806
rect 207032 84166 207520 84194
rect 207032 73166 207060 84166
rect 207020 73160 207072 73166
rect 207020 73102 207072 73108
rect 207032 66162 207060 73102
rect 207020 66156 207072 66162
rect 207020 66098 207072 66104
rect 205640 64796 205692 64802
rect 205640 64738 205692 64744
rect 205652 63578 205680 64738
rect 205640 63572 205692 63578
rect 205640 63514 205692 63520
rect 206284 63572 206336 63578
rect 206284 63514 206336 63520
rect 202144 56568 202196 56574
rect 202144 56510 202196 56516
rect 206296 54534 206324 63514
rect 206284 54528 206336 54534
rect 206284 54470 206336 54476
rect 208412 37942 208440 92806
rect 209240 88233 209268 92820
rect 209226 88224 209282 88233
rect 209226 88159 209282 88168
rect 209792 60654 209820 92820
rect 210344 89729 210372 92820
rect 210712 92806 211094 92834
rect 210330 89720 210386 89729
rect 210330 89655 210386 89664
rect 210712 84194 210740 92806
rect 211632 89729 211660 92820
rect 211724 92806 212198 92834
rect 212552 92820 212934 92834
rect 212552 92806 212948 92820
rect 211618 89720 211674 89729
rect 211618 89655 211674 89664
rect 211724 84194 211752 92806
rect 209884 84166 210740 84194
rect 211172 84166 211752 84194
rect 209884 81433 209912 84166
rect 209870 81424 209926 81433
rect 209870 81359 209926 81368
rect 211066 81424 211122 81433
rect 211066 81359 211122 81368
rect 211080 80753 211108 81359
rect 211066 80744 211122 80753
rect 211066 80679 211122 80688
rect 209780 60648 209832 60654
rect 209780 60590 209832 60596
rect 211068 60648 211120 60654
rect 211068 60590 211120 60596
rect 211080 56574 211108 60590
rect 211172 59362 211200 84166
rect 212552 71777 212580 92806
rect 212920 92546 212948 92806
rect 212908 92540 212960 92546
rect 212908 92482 212960 92488
rect 213288 92410 213316 93055
rect 224052 92834 224080 93366
rect 213380 92806 213486 92834
rect 213276 92404 213328 92410
rect 213276 92346 213328 92352
rect 213380 89010 213408 92806
rect 213368 89004 213420 89010
rect 213368 88946 213420 88952
rect 213380 84194 213408 88946
rect 214024 88330 214052 92820
rect 214012 88324 214064 88330
rect 214012 88266 214064 88272
rect 214576 85542 214604 92820
rect 215312 90386 215340 92820
rect 215220 90358 215340 90386
rect 215404 92806 215878 92834
rect 215220 89593 215248 90358
rect 215298 90264 215354 90273
rect 215298 90199 215354 90208
rect 215206 89584 215262 89593
rect 215206 89519 215262 89528
rect 214564 85536 214616 85542
rect 214564 85478 214616 85484
rect 213196 84166 213408 84194
rect 213196 74526 213224 84166
rect 214564 82136 214616 82142
rect 214564 82078 214616 82084
rect 213184 74520 213236 74526
rect 213184 74462 213236 74468
rect 212538 71768 212594 71777
rect 212538 71703 212594 71712
rect 212552 70417 212580 71703
rect 212538 70408 212594 70417
rect 212538 70343 212594 70352
rect 213182 70408 213238 70417
rect 213182 70343 213238 70352
rect 213196 64190 213224 70343
rect 213184 64184 213236 64190
rect 213184 64126 213236 64132
rect 211160 59356 211212 59362
rect 211160 59298 211212 59304
rect 212448 59356 212500 59362
rect 212448 59298 212500 59304
rect 212460 57866 212488 59298
rect 212448 57860 212500 57866
rect 212448 57802 212500 57808
rect 211068 56568 211120 56574
rect 211068 56510 211120 56516
rect 208400 37936 208452 37942
rect 208400 37878 208452 37884
rect 201408 13116 201460 13122
rect 201408 13058 201460 13064
rect 198004 10328 198056 10334
rect 198004 10270 198056 10276
rect 196624 8968 196676 8974
rect 196624 8910 196676 8916
rect 191748 6180 191800 6186
rect 191748 6122 191800 6128
rect 150624 3664 150676 3670
rect 150624 3606 150676 3612
rect 152464 3664 152516 3670
rect 152464 3606 152516 3612
rect 148508 3596 148560 3602
rect 148508 3538 148560 3544
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 142804 3460 142856 3466
rect 142804 3402 142856 3408
rect 143552 480 143580 3470
rect 147140 480 147168 3470
rect 150636 480 150664 3606
rect 214576 3466 214604 82078
rect 215312 64870 215340 90199
rect 215404 82006 215432 92806
rect 216416 90273 216444 92820
rect 217152 92478 217180 92820
rect 217140 92472 217192 92478
rect 217140 92414 217192 92420
rect 217152 91050 217180 92414
rect 217140 91044 217192 91050
rect 217140 90986 217192 90992
rect 216402 90264 216458 90273
rect 216402 90199 216458 90208
rect 217704 89690 217732 92820
rect 217692 89684 217744 89690
rect 217692 89626 217744 89632
rect 218256 86970 218284 92820
rect 218822 92806 219296 92834
rect 219558 92806 219848 92834
rect 219162 91080 219218 91089
rect 219162 91015 219218 91024
rect 218244 86964 218296 86970
rect 218244 86906 218296 86912
rect 219176 85377 219204 91015
rect 219268 90386 219296 92806
rect 219438 90400 219494 90409
rect 219268 90358 219438 90386
rect 219438 90335 219494 90344
rect 219162 85368 219218 85377
rect 219162 85303 219218 85312
rect 219452 84194 219480 90335
rect 219820 89593 219848 92806
rect 220096 91089 220124 92820
rect 220082 91080 220138 91089
rect 220082 91015 220138 91024
rect 220648 89690 220676 92820
rect 221384 90982 221412 92820
rect 222212 92806 222502 92834
rect 222672 92806 223054 92834
rect 223790 92820 224080 92834
rect 223776 92806 224080 92820
rect 221372 90976 221424 90982
rect 221372 90918 221424 90924
rect 220636 89684 220688 89690
rect 220636 89626 220688 89632
rect 219806 89584 219862 89593
rect 219806 89519 219862 89528
rect 219820 84194 219848 89519
rect 219452 84166 219572 84194
rect 219820 84166 220124 84194
rect 215392 82000 215444 82006
rect 215392 81942 215444 81948
rect 216036 82000 216088 82006
rect 216036 81942 216088 81948
rect 215300 64864 215352 64870
rect 215300 64806 215352 64812
rect 215312 63578 215340 64806
rect 215300 63572 215352 63578
rect 215300 63514 215352 63520
rect 215944 63572 215996 63578
rect 215944 63514 215996 63520
rect 215956 29646 215984 63514
rect 216048 62014 216076 81942
rect 216036 62008 216088 62014
rect 216036 61950 216088 61956
rect 219544 57934 219572 84166
rect 220096 82793 220124 84166
rect 220082 82784 220138 82793
rect 220082 82719 220138 82728
rect 222212 69018 222240 92806
rect 222672 84194 222700 92806
rect 223776 90574 223804 92806
rect 224328 91089 224356 92820
rect 224880 92478 224908 92820
rect 224868 92472 224920 92478
rect 224868 92414 224920 92420
rect 224314 91080 224370 91089
rect 224314 91015 224370 91024
rect 223764 90568 223816 90574
rect 223764 90510 223816 90516
rect 224868 90568 224920 90574
rect 224868 90510 224920 90516
rect 222304 84166 222700 84194
rect 222304 69086 222332 84166
rect 222292 69080 222344 69086
rect 222292 69022 222344 69028
rect 222200 69012 222252 69018
rect 222200 68954 222252 68960
rect 222304 67561 222332 69022
rect 222844 69012 222896 69018
rect 222844 68954 222896 68960
rect 222290 67552 222346 67561
rect 222290 67487 222346 67496
rect 219532 57928 219584 57934
rect 219532 57870 219584 57876
rect 220084 57928 220136 57934
rect 220084 57870 220136 57876
rect 215944 29640 215996 29646
rect 215944 29582 215996 29588
rect 220096 7614 220124 57870
rect 222856 19990 222884 68954
rect 222844 19984 222896 19990
rect 222844 19926 222896 19932
rect 220084 7608 220136 7614
rect 220084 7550 220136 7556
rect 224880 4865 224908 90510
rect 224972 81394 225000 109126
rect 225050 109103 225106 109112
rect 225156 103514 225184 114815
rect 225064 103486 225184 103514
rect 225064 89457 225092 103486
rect 225142 94752 225198 94761
rect 225142 94687 225198 94696
rect 225156 93430 225184 94687
rect 225144 93424 225196 93430
rect 225144 93366 225196 93372
rect 225616 90982 225644 231746
rect 227720 206304 227772 206310
rect 227720 206246 227772 206252
rect 227732 205766 227760 206246
rect 227720 205760 227772 205766
rect 227720 205702 227772 205708
rect 227732 200114 227760 205702
rect 228376 202162 228404 241604
rect 230492 241590 230782 241618
rect 230492 238649 230520 241590
rect 230478 238640 230534 238649
rect 230478 238575 230534 238584
rect 229100 227044 229152 227050
rect 229100 226986 229152 226992
rect 229928 227044 229980 227050
rect 229928 226986 229980 226992
rect 228364 202156 228416 202162
rect 228364 202098 228416 202104
rect 227732 200086 227852 200114
rect 226340 186992 226392 186998
rect 226340 186934 226392 186940
rect 225696 142180 225748 142186
rect 225696 142122 225748 142128
rect 225708 112470 225736 142122
rect 226156 115932 226208 115938
rect 226156 115874 226208 115880
rect 226168 114889 226196 115874
rect 226154 114880 226210 114889
rect 226154 114815 226210 114824
rect 226352 113174 226380 186934
rect 226430 171728 226486 171737
rect 226430 171663 226486 171672
rect 226444 134745 226472 171663
rect 226524 161560 226576 161566
rect 226524 161502 226576 161508
rect 226430 134736 226486 134745
rect 226430 134671 226486 134680
rect 226536 129146 226564 161502
rect 227720 157412 227772 157418
rect 227720 157354 227772 157360
rect 226614 146568 226670 146577
rect 226614 146503 226670 146512
rect 226628 136649 226656 146503
rect 226708 139256 226760 139262
rect 226708 139198 226760 139204
rect 226720 139097 226748 139198
rect 226706 139088 226762 139097
rect 226706 139023 226762 139032
rect 226708 137964 226760 137970
rect 226708 137906 226760 137912
rect 226720 137193 226748 137906
rect 226706 137184 226762 137193
rect 226706 137119 226762 137128
rect 226614 136640 226670 136649
rect 226614 136575 226670 136584
rect 226706 135552 226762 135561
rect 226706 135487 226762 135496
rect 226720 135250 226748 135487
rect 226708 135244 226760 135250
rect 226708 135186 226760 135192
rect 226614 134736 226670 134745
rect 226614 134671 226670 134680
rect 226628 134570 226656 134671
rect 226616 134564 226668 134570
rect 226616 134506 226668 134512
rect 226616 133884 226668 133890
rect 226616 133826 226668 133832
rect 226628 132841 226656 133826
rect 226708 133680 226760 133686
rect 226706 133648 226708 133657
rect 226760 133648 226762 133657
rect 226706 133583 226762 133592
rect 226614 132832 226670 132841
rect 226614 132767 226670 132776
rect 226708 132456 226760 132462
rect 226708 132398 226760 132404
rect 226720 132025 226748 132398
rect 226706 132016 226762 132025
rect 226706 131951 226762 131960
rect 226708 131096 226760 131102
rect 226708 131038 226760 131044
rect 226720 130937 226748 131038
rect 226800 131028 226852 131034
rect 226800 130970 226852 130976
rect 226706 130928 226762 130937
rect 226706 130863 226762 130872
rect 226812 130121 226840 130970
rect 226798 130112 226854 130121
rect 226798 130047 226854 130056
rect 226536 129118 226748 129146
rect 226614 129024 226670 129033
rect 226614 128959 226670 128968
rect 226430 128480 226486 128489
rect 226430 128415 226486 128424
rect 226444 128382 226472 128415
rect 226432 128376 226484 128382
rect 226432 128318 226484 128324
rect 226628 124681 226656 128959
rect 226720 127634 226748 129118
rect 226708 127628 226760 127634
rect 226708 127570 226760 127576
rect 226720 127401 226748 127570
rect 226706 127392 226762 127401
rect 226706 127327 226762 127336
rect 226708 126948 226760 126954
rect 226708 126890 226760 126896
rect 226720 126585 226748 126890
rect 226706 126576 226762 126585
rect 226706 126511 226762 126520
rect 226614 124672 226670 124681
rect 226614 124607 226670 124616
rect 226708 124160 226760 124166
rect 226708 124102 226760 124108
rect 226720 123049 226748 124102
rect 227626 123856 227682 123865
rect 227732 123842 227760 157354
rect 227682 123814 227760 123842
rect 227626 123791 227682 123800
rect 226706 123040 226762 123049
rect 226706 122975 226762 122984
rect 226524 122800 226576 122806
rect 226524 122742 226576 122748
rect 226536 122233 226564 122742
rect 226522 122224 226578 122233
rect 226522 122159 226578 122168
rect 226708 121440 226760 121446
rect 226708 121382 226760 121388
rect 226720 120329 226748 121382
rect 226706 120320 226762 120329
rect 226706 120255 226762 120264
rect 226522 118416 226578 118425
rect 226522 118351 226578 118360
rect 226536 117434 226564 118351
rect 226614 117600 226670 117609
rect 226614 117535 226670 117544
rect 226524 117428 226576 117434
rect 226524 117370 226576 117376
rect 226628 117366 226656 117535
rect 226616 117360 226668 117366
rect 226616 117302 226668 117308
rect 227626 116784 227682 116793
rect 227682 116742 227760 116770
rect 227626 116719 227682 116728
rect 226708 116000 226760 116006
rect 226706 115968 226708 115977
rect 226760 115968 226762 115977
rect 226706 115903 226762 115912
rect 226430 114064 226486 114073
rect 226430 113999 226486 114008
rect 226444 113898 226472 113999
rect 226432 113892 226484 113898
rect 226432 113834 226484 113840
rect 226352 113146 226472 113174
rect 225696 112464 225748 112470
rect 225696 112406 225748 112412
rect 226338 112160 226394 112169
rect 226338 112095 226394 112104
rect 226352 111858 226380 112095
rect 226340 111852 226392 111858
rect 226340 111794 226392 111800
rect 226340 111104 226392 111110
rect 226340 111046 226392 111052
rect 226352 110537 226380 111046
rect 226338 110528 226394 110537
rect 226338 110463 226394 110472
rect 226338 105904 226394 105913
rect 226338 105839 226394 105848
rect 226352 105602 226380 105839
rect 226340 105596 226392 105602
rect 226340 105538 226392 105544
rect 225696 104168 225748 104174
rect 225696 104110 225748 104116
rect 225708 93362 225736 104110
rect 226340 102128 226392 102134
rect 226340 102070 226392 102076
rect 226352 101561 226380 102070
rect 226338 101552 226394 101561
rect 226338 101487 226394 101496
rect 226338 99512 226394 99521
rect 226338 99447 226394 99456
rect 226352 99414 226380 99447
rect 226340 99408 226392 99414
rect 226340 99350 226392 99356
rect 226444 95169 226472 113146
rect 226708 111580 226760 111586
rect 226708 111522 226760 111528
rect 226720 111353 226748 111522
rect 226706 111344 226762 111353
rect 226706 111279 226762 111288
rect 226524 108928 226576 108934
rect 226524 108870 226576 108876
rect 226536 108633 226564 108870
rect 226522 108624 226578 108633
rect 226522 108559 226578 108568
rect 226984 108316 227036 108322
rect 226984 108258 227036 108264
rect 226708 107636 226760 107642
rect 226708 107578 226760 107584
rect 226720 107001 226748 107578
rect 226706 106992 226762 107001
rect 226706 106927 226762 106936
rect 226706 105088 226762 105097
rect 226706 105023 226708 105032
rect 226760 105023 226762 105032
rect 226708 104994 226760 105000
rect 226706 104272 226762 104281
rect 226706 104207 226762 104216
rect 226720 103562 226748 104207
rect 226708 103556 226760 103562
rect 226708 103498 226760 103504
rect 226706 103456 226762 103465
rect 226706 103391 226762 103400
rect 226720 102814 226748 103391
rect 226708 102808 226760 102814
rect 226708 102750 226760 102756
rect 226706 102368 226762 102377
rect 226706 102303 226762 102312
rect 226720 102202 226748 102303
rect 226708 102196 226760 102202
rect 226708 102138 226760 102144
rect 226708 101448 226760 101454
rect 226708 101390 226760 101396
rect 226720 98841 226748 101390
rect 226706 98832 226762 98841
rect 226762 98790 226840 98818
rect 226706 98767 226762 98776
rect 226616 98660 226668 98666
rect 226616 98602 226668 98608
rect 226628 98025 226656 98602
rect 226614 98016 226670 98025
rect 226614 97951 226670 97960
rect 226430 95160 226486 95169
rect 226430 95095 226486 95104
rect 225696 93356 225748 93362
rect 225696 93298 225748 93304
rect 226628 92410 226656 97951
rect 226708 96620 226760 96626
rect 226708 96562 226760 96568
rect 226720 96121 226748 96562
rect 226706 96112 226762 96121
rect 226706 96047 226762 96056
rect 226812 93854 226840 98790
rect 226996 97209 227024 108258
rect 227168 97300 227220 97306
rect 227168 97242 227220 97248
rect 226982 97200 227038 97209
rect 226982 97135 227038 97144
rect 227074 95160 227130 95169
rect 227074 95095 227130 95104
rect 226720 93826 226840 93854
rect 226616 92404 226668 92410
rect 226616 92346 226668 92352
rect 225604 90976 225656 90982
rect 225604 90918 225656 90924
rect 225050 89448 225106 89457
rect 225050 89383 225106 89392
rect 226720 84153 226748 93826
rect 226706 84144 226762 84153
rect 226706 84079 226762 84088
rect 226984 83564 227036 83570
rect 226984 83506 227036 83512
rect 224960 81388 225012 81394
rect 224960 81330 225012 81336
rect 224866 4856 224922 4865
rect 224866 4791 224922 4800
rect 214564 3460 214616 3466
rect 214564 3402 214616 3408
rect 226996 3369 227024 83506
rect 227088 82890 227116 95095
rect 227180 93673 227208 97242
rect 227166 93664 227222 93673
rect 227166 93599 227222 93608
rect 227076 82884 227128 82890
rect 227076 82826 227128 82832
rect 227088 79966 227116 82826
rect 227076 79960 227128 79966
rect 227076 79902 227128 79908
rect 227732 67590 227760 116742
rect 227824 92478 227852 200086
rect 228364 177336 228416 177342
rect 228364 177278 228416 177284
rect 228376 172650 228404 177278
rect 228364 172644 228416 172650
rect 228364 172586 228416 172592
rect 228376 144974 228404 172586
rect 229112 162897 229140 226986
rect 229940 226370 229968 226986
rect 229928 226364 229980 226370
rect 229928 226306 229980 226312
rect 229098 162888 229154 162897
rect 229098 162823 229154 162832
rect 229112 161474 229140 162823
rect 230492 162081 230520 238575
rect 231858 228848 231914 228857
rect 231858 228783 231914 228792
rect 231872 227769 231900 228783
rect 233160 227769 233188 241604
rect 235552 239426 235580 241604
rect 235540 239420 235592 239426
rect 235540 239362 235592 239368
rect 237944 233238 237972 241604
rect 237380 233232 237432 233238
rect 237380 233174 237432 233180
rect 237932 233232 237984 233238
rect 237932 233174 237984 233180
rect 236642 232520 236698 232529
rect 236642 232455 236698 232464
rect 231858 227760 231914 227769
rect 231858 227695 231914 227704
rect 233146 227760 233202 227769
rect 233146 227695 233202 227704
rect 230572 171148 230624 171154
rect 230572 171090 230624 171096
rect 230478 162072 230534 162081
rect 230478 162007 230534 162016
rect 229112 161446 229232 161474
rect 229100 156052 229152 156058
rect 229100 155994 229152 156000
rect 228364 144968 228416 144974
rect 227994 144936 228050 144945
rect 228364 144910 228416 144916
rect 227994 144871 228050 144880
rect 227902 129296 227958 129305
rect 227902 129231 227958 129240
rect 227916 127702 227944 129231
rect 227904 127696 227956 127702
rect 227904 127638 227956 127644
rect 227902 126984 227958 126993
rect 228008 126970 228036 144871
rect 228376 139913 228404 144910
rect 228362 139904 228418 139913
rect 228362 139839 228418 139848
rect 227958 126942 228036 126970
rect 227902 126919 227958 126928
rect 227916 125769 227944 126919
rect 227902 125760 227958 125769
rect 227902 125695 227958 125704
rect 229112 108934 229140 155994
rect 229204 139262 229232 161446
rect 230478 158808 230534 158817
rect 230478 158743 230534 158752
rect 229192 139256 229244 139262
rect 229192 139198 229244 139204
rect 230388 116680 230440 116686
rect 230388 116622 230440 116628
rect 230400 116006 230428 116622
rect 229192 116000 229244 116006
rect 229192 115942 229244 115948
rect 230388 116000 230440 116006
rect 230388 115942 230440 115948
rect 229100 108928 229152 108934
rect 229100 108870 229152 108876
rect 229100 103556 229152 103562
rect 229100 103498 229152 103504
rect 227902 100736 227958 100745
rect 227902 100671 227958 100680
rect 227812 92472 227864 92478
rect 227812 92414 227864 92420
rect 227916 73098 227944 100671
rect 227996 95940 228048 95946
rect 227996 95882 228048 95888
rect 228008 95305 228036 95882
rect 227994 95296 228050 95305
rect 227994 95231 228050 95240
rect 228008 75857 228036 95231
rect 229112 82822 229140 103498
rect 229100 82816 229152 82822
rect 229100 82758 229152 82764
rect 229204 77246 229232 115942
rect 230492 111586 230520 158743
rect 230584 124166 230612 171090
rect 231124 160812 231176 160818
rect 231124 160754 231176 160760
rect 230664 150476 230716 150482
rect 230664 150418 230716 150424
rect 230676 131102 230704 150418
rect 231136 133686 231164 160754
rect 231124 133680 231176 133686
rect 231124 133622 231176 133628
rect 230664 131096 230716 131102
rect 230664 131038 230716 131044
rect 230572 124160 230624 124166
rect 230572 124102 230624 124108
rect 231124 117428 231176 117434
rect 231124 117370 231176 117376
rect 230480 111580 230532 111586
rect 230480 111522 230532 111528
rect 231136 110430 231164 117370
rect 231124 110424 231176 110430
rect 231124 110366 231176 110372
rect 230572 105052 230624 105058
rect 230572 104994 230624 105000
rect 230480 102808 230532 102814
rect 230480 102750 230532 102756
rect 229192 77240 229244 77246
rect 229192 77182 229244 77188
rect 230492 75886 230520 102750
rect 230584 78606 230612 104994
rect 230572 78600 230624 78606
rect 230572 78542 230624 78548
rect 230480 75880 230532 75886
rect 227994 75848 228050 75857
rect 230480 75822 230532 75828
rect 227994 75783 228050 75792
rect 231136 73137 231164 110366
rect 231872 77897 231900 227695
rect 236656 220833 236684 232455
rect 237392 229094 237420 233174
rect 237300 229066 237420 229094
rect 236642 220824 236698 220833
rect 236642 220759 236698 220768
rect 236000 210520 236052 210526
rect 236000 210462 236052 210468
rect 236012 210361 236040 210462
rect 235998 210352 236054 210361
rect 235998 210287 236054 210296
rect 232504 188352 232556 188358
rect 232504 188294 232556 188300
rect 232516 153105 232544 188294
rect 234620 178696 234672 178702
rect 234620 178638 234672 178644
rect 231950 153096 232006 153105
rect 231950 153031 232006 153040
rect 232502 153096 232558 153105
rect 232502 153031 232558 153040
rect 231964 151881 231992 153031
rect 231950 151872 232006 151881
rect 231950 151807 232006 151816
rect 231964 135250 231992 151807
rect 233238 150648 233294 150657
rect 233238 150583 233294 150592
rect 232502 142352 232558 142361
rect 232502 142287 232558 142296
rect 231952 135244 232004 135250
rect 231952 135186 232004 135192
rect 232516 120766 232544 142287
rect 233252 131034 233280 150583
rect 233884 147688 233936 147694
rect 233884 147630 233936 147636
rect 233240 131028 233292 131034
rect 233240 130970 233292 130976
rect 232504 120760 232556 120766
rect 232504 120702 232556 120708
rect 231952 111852 232004 111858
rect 231952 111794 232004 111800
rect 231858 77888 231914 77897
rect 231858 77823 231914 77832
rect 231122 73128 231178 73137
rect 227904 73092 227956 73098
rect 231122 73063 231178 73072
rect 227904 73034 227956 73040
rect 227916 71806 227944 73034
rect 227904 71800 227956 71806
rect 227904 71742 227956 71748
rect 228364 71800 228416 71806
rect 228364 71742 228416 71748
rect 227720 67584 227772 67590
rect 227720 67526 227772 67532
rect 228376 4826 228404 71742
rect 231964 71738 231992 111794
rect 232594 77888 232650 77897
rect 232594 77823 232650 77832
rect 231952 71732 232004 71738
rect 231952 71674 232004 71680
rect 232608 54534 232636 77823
rect 232504 54528 232556 54534
rect 232504 54470 232556 54476
rect 232596 54528 232648 54534
rect 232596 54470 232648 54476
rect 228364 4820 228416 4826
rect 228364 4762 228416 4768
rect 232516 3534 232544 54470
rect 233896 32434 233924 147630
rect 234632 137970 234660 178638
rect 236012 169833 236040 210287
rect 235998 169824 236054 169833
rect 235998 169759 236054 169768
rect 234712 145580 234764 145586
rect 234712 145522 234764 145528
rect 234620 137964 234672 137970
rect 234620 137906 234672 137912
rect 234724 121446 234752 145522
rect 236012 138961 236040 169759
rect 235998 138952 236054 138961
rect 235998 138887 236054 138896
rect 236012 138718 236040 138887
rect 236000 138712 236052 138718
rect 236000 138654 236052 138660
rect 235264 123480 235316 123486
rect 235264 123422 235316 123428
rect 234712 121440 234764 121446
rect 234712 121382 234764 121388
rect 235276 89010 235304 123422
rect 237300 98666 237328 229066
rect 238024 228404 238076 228410
rect 238024 228346 238076 228352
rect 237380 171828 237432 171834
rect 237380 171770 237432 171776
rect 237392 164393 237420 171770
rect 238036 167686 238064 228346
rect 239404 217320 239456 217326
rect 239404 217262 239456 217268
rect 238024 167680 238076 167686
rect 238024 167622 238076 167628
rect 237378 164384 237434 164393
rect 237378 164319 237434 164328
rect 237392 133890 237420 164319
rect 238116 144220 238168 144226
rect 238116 144162 238168 144168
rect 238022 140856 238078 140865
rect 238022 140791 238078 140800
rect 237380 133884 237432 133890
rect 237380 133826 237432 133832
rect 237380 102196 237432 102202
rect 237380 102138 237432 102144
rect 237288 98660 237340 98666
rect 237288 98602 237340 98608
rect 235264 89004 235316 89010
rect 235264 88946 235316 88952
rect 233884 32428 233936 32434
rect 233884 32370 233936 32376
rect 235276 24138 235304 88946
rect 237392 74458 237420 102138
rect 237380 74452 237432 74458
rect 237380 74394 237432 74400
rect 237392 73234 237420 74394
rect 237380 73228 237432 73234
rect 237380 73170 237432 73176
rect 235264 24132 235316 24138
rect 235264 24074 235316 24080
rect 238036 17270 238064 140791
rect 238128 124914 238156 144162
rect 238116 124908 238168 124914
rect 238116 124850 238168 124856
rect 239416 90409 239444 217262
rect 240230 154456 240286 154465
rect 240230 154391 240286 154400
rect 240244 153241 240272 154391
rect 240230 153232 240286 153241
rect 240230 153167 240286 153176
rect 240244 122806 240272 153167
rect 240336 149161 240364 241604
rect 242728 240009 242756 241604
rect 244922 241088 244978 241097
rect 244922 241023 244978 241032
rect 242254 240000 242310 240009
rect 242254 239935 242310 239944
rect 242714 240000 242770 240009
rect 242714 239935 242770 239944
rect 242164 232552 242216 232558
rect 242164 232494 242216 232500
rect 241426 224224 241482 224233
rect 241426 224159 241482 224168
rect 241440 178702 241468 224159
rect 241428 178696 241480 178702
rect 241428 178638 241480 178644
rect 241440 178090 241468 178638
rect 240784 178084 240836 178090
rect 240784 178026 240836 178032
rect 241428 178084 241480 178090
rect 241428 178026 241480 178032
rect 240796 154465 240824 178026
rect 240782 154456 240838 154465
rect 240782 154391 240838 154400
rect 240322 149152 240378 149161
rect 240322 149087 240378 149096
rect 240782 149152 240838 149161
rect 240782 149087 240838 149096
rect 240796 131782 240824 149087
rect 240876 137964 240928 137970
rect 240876 137906 240928 137912
rect 240784 131776 240836 131782
rect 240784 131718 240836 131724
rect 240232 122800 240284 122806
rect 240232 122742 240284 122748
rect 240784 120828 240836 120834
rect 240784 120770 240836 120776
rect 240796 105602 240824 120770
rect 240784 105596 240836 105602
rect 240784 105538 240836 105544
rect 239402 90400 239458 90409
rect 239402 90335 239458 90344
rect 238116 73228 238168 73234
rect 238116 73170 238168 73176
rect 238024 17264 238076 17270
rect 238024 17206 238076 17212
rect 238128 4894 238156 73170
rect 240140 58676 240192 58682
rect 240140 58618 240192 58624
rect 238116 4888 238168 4894
rect 238116 4830 238168 4836
rect 239312 4888 239364 4894
rect 239312 4830 239364 4836
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 226982 3360 227038 3369
rect 226982 3295 227038 3304
rect 239324 480 239352 4830
rect 240152 490 240180 58618
rect 240796 18698 240824 105538
rect 240888 60110 240916 137906
rect 241520 82884 241572 82890
rect 241520 82826 241572 82832
rect 240876 60104 240928 60110
rect 240876 60046 240928 60052
rect 240784 18692 240836 18698
rect 240784 18634 240836 18640
rect 241532 16574 241560 82826
rect 242176 82142 242204 232494
rect 242268 92546 242296 239935
rect 244936 217977 244964 241023
rect 244922 217968 244978 217977
rect 244922 217903 244978 217912
rect 244924 214600 244976 214606
rect 244924 214542 244976 214548
rect 243544 200796 243596 200802
rect 243544 200738 243596 200744
rect 243556 123486 243584 200738
rect 244936 195974 244964 214542
rect 244924 195968 244976 195974
rect 244924 195910 244976 195916
rect 243544 123480 243596 123486
rect 243544 123422 243596 123428
rect 244280 117360 244332 117366
rect 244280 117302 244332 117308
rect 242256 92540 242308 92546
rect 242256 92482 242308 92488
rect 242164 82136 242216 82142
rect 242164 82078 242216 82084
rect 242176 21418 242204 82078
rect 244292 70310 244320 117302
rect 244936 95946 244964 195910
rect 245120 146985 245148 241604
rect 247512 239465 247540 241604
rect 249064 240644 249116 240650
rect 249064 240586 249116 240592
rect 247498 239456 247554 239465
rect 247498 239391 247554 239400
rect 247774 238096 247830 238105
rect 247774 238031 247830 238040
rect 246394 236872 246450 236881
rect 246394 236807 246450 236816
rect 246304 231124 246356 231130
rect 246304 231066 246356 231072
rect 245106 146976 245162 146985
rect 245106 146911 245162 146920
rect 245016 143608 245068 143614
rect 245016 143550 245068 143556
rect 245028 116618 245056 143550
rect 245016 116612 245068 116618
rect 245016 116554 245068 116560
rect 246316 113174 246344 231066
rect 246408 199345 246436 236807
rect 247684 232620 247736 232626
rect 247684 232562 247736 232568
rect 246394 199336 246450 199345
rect 246394 199271 246450 199280
rect 247696 175302 247724 232562
rect 247788 216578 247816 238031
rect 247776 216572 247828 216578
rect 247776 216514 247828 216520
rect 249076 184210 249104 240586
rect 249154 239456 249210 239465
rect 249154 239391 249210 239400
rect 249168 217326 249196 239391
rect 249156 217320 249208 217326
rect 249156 217262 249208 217268
rect 249708 199436 249760 199442
rect 249708 199378 249760 199384
rect 249064 184204 249116 184210
rect 249064 184146 249116 184152
rect 247684 175296 247736 175302
rect 247684 175238 247736 175244
rect 246396 155984 246448 155990
rect 246396 155926 246448 155932
rect 246408 113830 246436 155926
rect 247696 137290 247724 175238
rect 249616 159452 249668 159458
rect 249616 159394 249668 159400
rect 249628 158710 249656 159394
rect 249616 158704 249668 158710
rect 249616 158646 249668 158652
rect 249064 144220 249116 144226
rect 249064 144162 249116 144168
rect 247684 137284 247736 137290
rect 247684 137226 247736 137232
rect 246396 113824 246448 113830
rect 246396 113766 246448 113772
rect 246316 113146 246436 113174
rect 245016 105596 245068 105602
rect 245016 105538 245068 105544
rect 244924 95940 244976 95946
rect 244924 95882 244976 95888
rect 245028 89690 245056 105538
rect 246408 91050 246436 113146
rect 246488 98796 246540 98802
rect 246488 98738 246540 98744
rect 246396 91044 246448 91050
rect 246396 90986 246448 90992
rect 245016 89684 245068 89690
rect 245016 89626 245068 89632
rect 246304 87644 246356 87650
rect 246304 87586 246356 87592
rect 244280 70304 244332 70310
rect 244280 70246 244332 70252
rect 244292 69902 244320 70246
rect 244280 69896 244332 69902
rect 244280 69838 244332 69844
rect 244924 69896 244976 69902
rect 244924 69838 244976 69844
rect 244280 60036 244332 60042
rect 244280 59978 244332 59984
rect 242164 21412 242216 21418
rect 242164 21354 242216 21360
rect 242992 18624 243044 18630
rect 242992 18566 243044 18572
rect 243004 16574 243032 18566
rect 241532 16546 241744 16574
rect 243004 16546 244136 16574
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 16546
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 242912 480 242940 3470
rect 244108 480 244136 16546
rect 244292 6914 244320 59978
rect 244936 15910 244964 69838
rect 244924 15904 244976 15910
rect 244924 15846 244976 15852
rect 244292 6886 245240 6914
rect 245212 480 245240 6886
rect 246316 2990 246344 87586
rect 246408 11762 246436 90986
rect 246500 85542 246528 98738
rect 247684 98660 247736 98666
rect 247684 98602 247736 98608
rect 247696 93158 247724 98602
rect 247684 93152 247736 93158
rect 247684 93094 247736 93100
rect 246488 85536 246540 85542
rect 246488 85478 246540 85484
rect 249076 75206 249104 144162
rect 249720 139466 249748 199378
rect 249812 160750 249840 241998
rect 250166 241975 250222 241984
rect 251836 241590 252310 241618
rect 250444 240780 250496 240786
rect 250444 240722 250496 240728
rect 249890 236600 249946 236609
rect 249890 236535 249946 236544
rect 249800 160744 249852 160750
rect 249800 160686 249852 160692
rect 249708 139460 249760 139466
rect 249708 139402 249760 139408
rect 249812 126954 249840 160686
rect 249904 160177 249932 236535
rect 249890 160168 249946 160177
rect 249890 160103 249946 160112
rect 249904 132462 249932 160103
rect 249892 132456 249944 132462
rect 249892 132398 249944 132404
rect 249800 126948 249852 126954
rect 249800 126890 249852 126896
rect 248420 75200 248472 75206
rect 248420 75142 248472 75148
rect 249064 75200 249116 75206
rect 249064 75142 249116 75148
rect 246396 11756 246448 11762
rect 246396 11698 246448 11704
rect 246396 3460 246448 3466
rect 246396 3402 246448 3408
rect 246304 2984 246356 2990
rect 246304 2926 246356 2932
rect 246408 480 246436 3402
rect 247592 2984 247644 2990
rect 247592 2926 247644 2932
rect 247604 480 247632 2926
rect 248432 490 248460 75142
rect 250456 66230 250484 240722
rect 251836 239873 251864 241590
rect 251822 239864 251878 239873
rect 251822 239799 251878 239808
rect 251836 238649 251864 239799
rect 252100 239216 252152 239222
rect 252100 239158 252152 239164
rect 251822 238640 251878 238649
rect 251822 238575 251878 238584
rect 251836 177342 251864 238575
rect 252112 232529 252140 239158
rect 252388 236774 252416 242286
rect 252468 239420 252520 239426
rect 252468 239362 252520 239368
rect 252376 236768 252428 236774
rect 252376 236710 252428 236716
rect 252098 232520 252154 232529
rect 252098 232455 252154 232464
rect 251824 177336 251876 177342
rect 251824 177278 251876 177284
rect 252480 149802 252508 239362
rect 252572 224262 252600 297622
rect 252834 297599 252890 297608
rect 252834 293448 252890 293457
rect 252834 293383 252890 293392
rect 252848 292574 252876 293383
rect 252664 292546 252876 292574
rect 252560 224256 252612 224262
rect 252560 224198 252612 224204
rect 252560 221468 252612 221474
rect 252560 221410 252612 221416
rect 252572 220969 252600 221410
rect 252558 220960 252614 220969
rect 252558 220895 252614 220904
rect 252468 149796 252520 149802
rect 252468 149738 252520 149744
rect 252480 149190 252508 149738
rect 252468 149184 252520 149190
rect 252468 149126 252520 149132
rect 252192 146940 252244 146946
rect 252192 146882 252244 146888
rect 252204 145625 252232 146882
rect 252190 145616 252246 145625
rect 252190 145551 252246 145560
rect 251180 139460 251232 139466
rect 251180 139402 251232 139408
rect 251088 126948 251140 126954
rect 251088 126890 251140 126896
rect 251100 126274 251128 126890
rect 251088 126268 251140 126274
rect 251088 126210 251140 126216
rect 250536 122120 250588 122126
rect 250536 122062 250588 122068
rect 250548 113898 250576 122062
rect 250536 113892 250588 113898
rect 250536 113834 250588 113840
rect 250444 66224 250496 66230
rect 250444 66166 250496 66172
rect 250548 49094 250576 113834
rect 250536 49088 250588 49094
rect 250536 49030 250588 49036
rect 249800 43444 249852 43450
rect 249800 43386 249852 43392
rect 249812 16574 249840 43386
rect 249812 16546 250024 16574
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 251192 3602 251220 139402
rect 252572 120834 252600 220895
rect 252664 220114 252692 292546
rect 252940 291938 252968 302206
rect 253400 301594 253428 304982
rect 253952 302234 253980 342858
rect 253952 302206 254256 302234
rect 253230 301566 253428 301594
rect 254124 301504 254176 301510
rect 254124 301446 254176 301452
rect 253938 300656 253994 300665
rect 253938 300591 253994 300600
rect 253020 299464 253072 299470
rect 253020 299406 253072 299412
rect 253032 298897 253060 299406
rect 253018 298888 253074 298897
rect 253018 298823 253074 298832
rect 253032 297673 253060 298823
rect 253018 297664 253074 297673
rect 253018 297599 253074 297608
rect 253952 296585 253980 300591
rect 254032 300144 254084 300150
rect 254032 300086 254084 300092
rect 253938 296576 253994 296585
rect 253938 296511 253994 296520
rect 254044 295633 254072 300086
rect 254030 295624 254086 295633
rect 254030 295559 254086 295568
rect 254136 293185 254164 301446
rect 254228 299849 254256 302206
rect 254582 301744 254638 301753
rect 254582 301679 254638 301688
rect 254214 299840 254270 299849
rect 254214 299775 254270 299784
rect 254122 293176 254178 293185
rect 254122 293111 254178 293120
rect 252756 291910 252968 291938
rect 252756 287054 252784 291910
rect 252756 287026 252876 287054
rect 252848 265577 252876 287026
rect 252834 265568 252890 265577
rect 252834 265503 252890 265512
rect 253846 265296 253902 265305
rect 253846 265231 253902 265240
rect 253860 264994 253888 265231
rect 253848 264988 253900 264994
rect 253848 264930 253900 264936
rect 252834 258768 252890 258777
rect 252834 258703 252890 258712
rect 252848 248414 252876 258703
rect 254596 255338 254624 301679
rect 255332 300393 255360 358702
rect 256804 356726 256832 497422
rect 256884 474020 256936 474026
rect 256884 473962 256936 473968
rect 256896 432682 256924 473962
rect 258092 472054 258120 549850
rect 258184 534818 258212 582354
rect 259552 577108 259604 577114
rect 259552 577050 259604 577056
rect 259460 564460 259512 564466
rect 259460 564402 259512 564408
rect 258356 545284 258408 545290
rect 258356 545226 258408 545232
rect 258172 534812 258224 534818
rect 258172 534754 258224 534760
rect 258264 527944 258316 527950
rect 258264 527886 258316 527892
rect 258170 475416 258226 475425
rect 258170 475351 258226 475360
rect 258080 472048 258132 472054
rect 258080 471990 258132 471996
rect 258092 454714 258120 471990
rect 258080 454708 258132 454714
rect 258080 454650 258132 454656
rect 258080 454096 258132 454102
rect 258080 454038 258132 454044
rect 257344 451376 257396 451382
rect 257344 451318 257396 451324
rect 256884 432676 256936 432682
rect 256884 432618 256936 432624
rect 256882 404016 256938 404025
rect 256882 403951 256938 403960
rect 256896 403034 256924 403951
rect 256884 403028 256936 403034
rect 256884 402970 256936 402976
rect 256896 383654 256924 402970
rect 256884 383648 256936 383654
rect 256884 383590 256936 383596
rect 256792 356720 256844 356726
rect 256792 356662 256844 356668
rect 256884 325032 256936 325038
rect 256884 324974 256936 324980
rect 255504 324964 255556 324970
rect 255504 324906 255556 324912
rect 255412 311160 255464 311166
rect 255412 311102 255464 311108
rect 255318 300384 255374 300393
rect 255318 300319 255374 300328
rect 255332 300218 255360 300319
rect 255320 300212 255372 300218
rect 255320 300154 255372 300160
rect 255318 297800 255374 297809
rect 255318 297735 255374 297744
rect 255332 296750 255360 297735
rect 255320 296744 255372 296750
rect 255320 296686 255372 296692
rect 255320 288312 255372 288318
rect 255320 288254 255372 288260
rect 255332 287609 255360 288254
rect 255318 287600 255374 287609
rect 255318 287535 255374 287544
rect 255424 287054 255452 311102
rect 255516 292574 255544 324906
rect 256792 318096 256844 318102
rect 256792 318038 256844 318044
rect 256700 315308 256752 315314
rect 256700 315250 256752 315256
rect 256712 314770 256740 315250
rect 256700 314764 256752 314770
rect 256700 314706 256752 314712
rect 255596 308440 255648 308446
rect 255596 308382 255648 308388
rect 255608 296177 255636 308382
rect 256804 302234 256832 318038
rect 256896 306374 256924 324974
rect 257356 309874 257384 451318
rect 257436 315308 257488 315314
rect 257436 315250 257488 315256
rect 257344 309868 257396 309874
rect 257344 309810 257396 309816
rect 256896 306346 257016 306374
rect 256804 302206 256924 302234
rect 256606 298208 256662 298217
rect 256606 298143 256608 298152
rect 256660 298143 256662 298152
rect 256608 298114 256660 298120
rect 255594 296168 255650 296177
rect 255594 296103 255650 296112
rect 256606 296168 256662 296177
rect 256606 296103 256662 296112
rect 256620 296070 256648 296103
rect 256608 296064 256660 296070
rect 256608 296006 256660 296012
rect 256608 295316 256660 295322
rect 256608 295258 256660 295264
rect 256330 294808 256386 294817
rect 256330 294743 256386 294752
rect 256344 294030 256372 294743
rect 256620 294409 256648 295258
rect 256606 294400 256662 294409
rect 256606 294335 256662 294344
rect 256332 294024 256384 294030
rect 256332 293966 256384 293972
rect 255964 293276 256016 293282
rect 255964 293218 256016 293224
rect 255976 292641 256004 293218
rect 256146 293176 256202 293185
rect 256146 293111 256148 293120
rect 256200 293111 256202 293120
rect 256148 293082 256200 293088
rect 255962 292632 256018 292641
rect 255516 292546 255728 292574
rect 255962 292567 256018 292576
rect 255700 291689 255728 292546
rect 256896 292194 256924 302206
rect 255964 292188 256016 292194
rect 255964 292130 256016 292136
rect 256884 292188 256936 292194
rect 256884 292130 256936 292136
rect 255976 291825 256004 292130
rect 255962 291816 256018 291825
rect 255962 291751 256018 291760
rect 255686 291680 255742 291689
rect 255686 291615 255742 291624
rect 256606 291136 256662 291145
rect 256988 291122 257016 306346
rect 257344 291848 257396 291854
rect 257344 291790 257396 291796
rect 256662 291094 257016 291122
rect 256606 291071 256662 291080
rect 255504 291032 255556 291038
rect 255504 290974 255556 290980
rect 255516 290057 255544 290974
rect 255502 290048 255558 290057
rect 255502 289983 255558 289992
rect 255504 289740 255556 289746
rect 255504 289682 255556 289688
rect 255516 289241 255544 289682
rect 255502 289232 255558 289241
rect 255502 289167 255558 289176
rect 255504 288380 255556 288386
rect 255504 288322 255556 288328
rect 255516 288017 255544 288322
rect 255502 288008 255558 288017
rect 255502 287943 255558 287952
rect 255332 287026 255452 287054
rect 255332 266121 255360 287026
rect 257356 286686 257384 291790
rect 257448 287065 257476 315250
rect 258092 305114 258120 454038
rect 258184 355434 258212 475351
rect 258276 468518 258304 527886
rect 258368 521665 258396 545226
rect 258354 521656 258410 521665
rect 258354 521591 258410 521600
rect 258264 468512 258316 468518
rect 258264 468454 258316 468460
rect 258276 412486 258304 468454
rect 258724 447500 258776 447506
rect 258724 447442 258776 447448
rect 258736 432614 258764 447442
rect 258724 432608 258776 432614
rect 258724 432550 258776 432556
rect 258264 412480 258316 412486
rect 258264 412422 258316 412428
rect 258908 398268 258960 398274
rect 258908 398210 258960 398216
rect 258920 395321 258948 398210
rect 258906 395312 258962 395321
rect 258906 395247 258962 395256
rect 258724 373380 258776 373386
rect 258724 373322 258776 373328
rect 258172 355428 258224 355434
rect 258172 355370 258224 355376
rect 258172 329860 258224 329866
rect 258172 329802 258224 329808
rect 258080 305108 258132 305114
rect 258080 305050 258132 305056
rect 258184 291038 258212 329802
rect 258736 325009 258764 373322
rect 259472 369170 259500 564402
rect 259564 539714 259592 577050
rect 260760 552702 260788 585142
rect 260748 552696 260800 552702
rect 260748 552638 260800 552644
rect 259644 550724 259696 550730
rect 259644 550666 259696 550672
rect 259552 539708 259604 539714
rect 259552 539650 259604 539656
rect 259550 526416 259606 526425
rect 259550 526351 259606 526360
rect 259460 369164 259512 369170
rect 259460 369106 259512 369112
rect 259564 354006 259592 526351
rect 259656 476814 259684 550666
rect 260840 536104 260892 536110
rect 260840 536046 260892 536052
rect 259644 476808 259696 476814
rect 259644 476750 259696 476756
rect 259656 464438 259684 476750
rect 259644 464432 259696 464438
rect 259644 464374 259696 464380
rect 259736 460964 259788 460970
rect 259736 460906 259788 460912
rect 259644 450492 259696 450498
rect 259644 450434 259696 450440
rect 259656 413846 259684 450434
rect 259748 435402 259776 460906
rect 260564 443692 260616 443698
rect 260564 443634 260616 443640
rect 260576 442270 260604 443634
rect 260564 442264 260616 442270
rect 260564 442206 260616 442212
rect 259736 435396 259788 435402
rect 259736 435338 259788 435344
rect 259644 413840 259696 413846
rect 259644 413782 259696 413788
rect 260104 411936 260156 411942
rect 260104 411878 260156 411884
rect 259644 407856 259696 407862
rect 259644 407798 259696 407804
rect 259656 390590 259684 407798
rect 259644 390584 259696 390590
rect 259644 390526 259696 390532
rect 260116 389298 260144 411878
rect 260104 389292 260156 389298
rect 260104 389234 260156 389240
rect 260104 363724 260156 363730
rect 260104 363666 260156 363672
rect 259552 354000 259604 354006
rect 259552 353942 259604 353948
rect 260116 331974 260144 363666
rect 260852 359514 260880 536046
rect 260932 530596 260984 530602
rect 260932 530538 260984 530544
rect 260944 387802 260972 530538
rect 261036 529145 261064 593370
rect 262404 589348 262456 589354
rect 262404 589290 262456 589296
rect 262220 579760 262272 579766
rect 262220 579702 262272 579708
rect 261022 529136 261078 529145
rect 261022 529071 261078 529080
rect 261022 452976 261078 452985
rect 261022 452911 261078 452920
rect 260932 387796 260984 387802
rect 260932 387738 260984 387744
rect 260840 359508 260892 359514
rect 260840 359450 260892 359456
rect 261036 337482 261064 452911
rect 261114 446448 261170 446457
rect 261114 446383 261170 446392
rect 261128 384849 261156 446383
rect 261114 384840 261170 384849
rect 261114 384775 261170 384784
rect 262232 358057 262260 579702
rect 262312 547936 262364 547942
rect 262312 547878 262364 547884
rect 262324 370705 262352 547878
rect 262416 501702 262444 589290
rect 262404 501696 262456 501702
rect 262404 501638 262456 501644
rect 262864 465724 262916 465730
rect 262864 465666 262916 465672
rect 262404 452668 262456 452674
rect 262404 452610 262456 452616
rect 262416 388385 262444 452610
rect 262876 442338 262904 465666
rect 262864 442332 262916 442338
rect 262864 442274 262916 442280
rect 263612 389065 263640 603094
rect 266372 585206 266400 697546
rect 266360 585200 266412 585206
rect 266360 585142 266412 585148
rect 266360 583772 266412 583778
rect 266360 583714 266412 583720
rect 263692 556232 263744 556238
rect 263692 556174 263744 556180
rect 263598 389056 263654 389065
rect 263598 388991 263654 389000
rect 262864 388476 262916 388482
rect 262864 388418 262916 388424
rect 262402 388376 262458 388385
rect 262402 388311 262458 388320
rect 262876 386374 262904 388418
rect 262864 386368 262916 386374
rect 262864 386310 262916 386316
rect 262310 370696 262366 370705
rect 262310 370631 262366 370640
rect 263704 367810 263732 556174
rect 265072 552696 265124 552702
rect 265072 552638 265124 552644
rect 264980 542496 265032 542502
rect 264980 542438 265032 542444
rect 263784 420232 263836 420238
rect 263784 420174 263836 420180
rect 264888 420232 264940 420238
rect 264888 420174 264940 420180
rect 263796 419558 263824 420174
rect 263784 419552 263836 419558
rect 263784 419494 263836 419500
rect 264244 391264 264296 391270
rect 264244 391206 264296 391212
rect 264256 378146 264284 391206
rect 264244 378140 264296 378146
rect 264244 378082 264296 378088
rect 263692 367804 263744 367810
rect 263692 367746 263744 367752
rect 262218 358048 262274 358057
rect 262218 357983 262274 357992
rect 262404 354068 262456 354074
rect 262404 354010 262456 354016
rect 261024 337476 261076 337482
rect 261024 337418 261076 337424
rect 260104 331968 260156 331974
rect 260104 331910 260156 331916
rect 259460 330540 259512 330546
rect 259460 330482 259512 330488
rect 258722 325000 258778 325009
rect 258722 324935 258778 324944
rect 258724 305108 258776 305114
rect 258724 305050 258776 305056
rect 258264 304836 258316 304842
rect 258264 304778 258316 304784
rect 258172 291032 258224 291038
rect 258172 290974 258224 290980
rect 258170 290864 258226 290873
rect 258170 290799 258226 290808
rect 257434 287056 257490 287065
rect 257434 286991 257490 287000
rect 255412 286680 255464 286686
rect 255410 286648 255412 286657
rect 257344 286680 257396 286686
rect 255464 286648 255466 286657
rect 257344 286622 257396 286628
rect 255410 286583 255466 286592
rect 257448 286521 257476 286991
rect 257434 286512 257490 286521
rect 257434 286447 257490 286456
rect 255504 286340 255556 286346
rect 255504 286282 255556 286288
rect 255516 286249 255544 286282
rect 255502 286240 255558 286249
rect 255502 286175 255558 286184
rect 256698 286104 256754 286113
rect 256698 286039 256754 286048
rect 255412 285660 255464 285666
rect 255412 285602 255464 285608
rect 255424 285433 255452 285602
rect 255410 285424 255466 285433
rect 255410 285359 255466 285368
rect 255412 284300 255464 284306
rect 255412 284242 255464 284248
rect 255424 284073 255452 284242
rect 255410 284064 255466 284073
rect 255410 283999 255466 284008
rect 255504 283416 255556 283422
rect 255504 283358 255556 283364
rect 255516 283257 255544 283358
rect 255502 283248 255558 283257
rect 255502 283183 255558 283192
rect 255504 282872 255556 282878
rect 255504 282814 255556 282820
rect 255410 282432 255466 282441
rect 255410 282367 255466 282376
rect 255424 281994 255452 282367
rect 255516 282033 255544 282814
rect 255502 282024 255558 282033
rect 255412 281988 255464 281994
rect 255502 281959 255558 281968
rect 255412 281930 255464 281936
rect 255504 281512 255556 281518
rect 255410 281480 255466 281489
rect 255504 281454 255556 281460
rect 255410 281415 255412 281424
rect 255464 281415 255466 281424
rect 255412 281386 255464 281392
rect 255516 280265 255544 281454
rect 255502 280256 255558 280265
rect 255502 280191 255558 280200
rect 255504 280152 255556 280158
rect 255504 280094 255556 280100
rect 255516 279041 255544 280094
rect 255502 279032 255558 279041
rect 255502 278967 255558 278976
rect 255412 278724 255464 278730
rect 255412 278666 255464 278672
rect 255424 277681 255452 278666
rect 255504 278656 255556 278662
rect 255504 278598 255556 278604
rect 255516 278497 255544 278598
rect 255502 278488 255558 278497
rect 255502 278423 255558 278432
rect 255410 277672 255466 277681
rect 255410 277607 255466 277616
rect 255502 277400 255558 277409
rect 255502 277335 255558 277344
rect 255596 277364 255648 277370
rect 255516 276865 255544 277335
rect 255596 277306 255648 277312
rect 255502 276856 255558 276865
rect 255502 276791 255558 276800
rect 255412 276684 255464 276690
rect 255412 276626 255464 276632
rect 255424 276049 255452 276626
rect 255608 276457 255636 277306
rect 255594 276448 255650 276457
rect 255594 276383 255650 276392
rect 255410 276040 255466 276049
rect 255410 275975 255466 275984
rect 255504 276004 255556 276010
rect 255504 275946 255556 275952
rect 255516 275097 255544 275946
rect 255502 275088 255558 275097
rect 255502 275023 255558 275032
rect 255412 274712 255464 274718
rect 255410 274680 255412 274689
rect 255464 274680 255466 274689
rect 255410 274615 255466 274624
rect 255504 274644 255556 274650
rect 255504 274586 255556 274592
rect 255412 274304 255464 274310
rect 255410 274272 255412 274281
rect 255464 274272 255466 274281
rect 255410 274207 255466 274216
rect 255516 273873 255544 274586
rect 255502 273864 255558 273873
rect 255502 273799 255558 273808
rect 255412 273216 255464 273222
rect 255412 273158 255464 273164
rect 255424 272513 255452 273158
rect 255410 272504 255466 272513
rect 255410 272439 255466 272448
rect 255410 272096 255466 272105
rect 255410 272031 255466 272040
rect 255424 271930 255452 272031
rect 255412 271924 255464 271930
rect 255412 271866 255464 271872
rect 255504 271856 255556 271862
rect 255504 271798 255556 271804
rect 255516 271289 255544 271798
rect 255502 271280 255558 271289
rect 255502 271215 255558 271224
rect 255412 270292 255464 270298
rect 255412 270234 255464 270240
rect 255424 269929 255452 270234
rect 255410 269920 255466 269929
rect 255410 269855 255466 269864
rect 255410 269512 255466 269521
rect 255410 269447 255466 269456
rect 255424 269210 255452 269447
rect 255412 269204 255464 269210
rect 255412 269146 255464 269152
rect 255412 268388 255464 268394
rect 255412 268330 255464 268336
rect 255424 268297 255452 268330
rect 255410 268288 255466 268297
rect 255410 268223 255466 268232
rect 255410 267880 255466 267889
rect 255410 267815 255466 267824
rect 255424 267782 255452 267815
rect 255412 267776 255464 267782
rect 255412 267718 255464 267724
rect 255410 266928 255466 266937
rect 255410 266863 255466 266872
rect 255424 266422 255452 266863
rect 255412 266416 255464 266422
rect 255412 266358 255464 266364
rect 255318 266112 255374 266121
rect 255318 266047 255374 266056
rect 255332 265674 255360 266047
rect 255320 265668 255372 265674
rect 255320 265610 255372 265616
rect 255502 264344 255558 264353
rect 255502 264279 255558 264288
rect 255412 264240 255464 264246
rect 255412 264182 255464 264188
rect 255424 263945 255452 264182
rect 255410 263936 255466 263945
rect 255410 263871 255466 263880
rect 255516 263634 255544 264279
rect 255504 263628 255556 263634
rect 255504 263570 255556 263576
rect 255412 263560 255464 263566
rect 255412 263502 255464 263508
rect 255502 263528 255558 263537
rect 255424 262313 255452 263502
rect 255502 263463 255558 263472
rect 255686 263528 255742 263537
rect 255686 263463 255742 263472
rect 255516 262886 255544 263463
rect 255504 262880 255556 262886
rect 255504 262822 255556 262828
rect 255700 262721 255728 263463
rect 255686 262712 255742 262721
rect 255686 262647 255742 262656
rect 255410 262304 255466 262313
rect 255410 262239 255466 262248
rect 255504 261520 255556 261526
rect 255504 261462 255556 261468
rect 255516 261361 255544 261462
rect 255502 261352 255558 261361
rect 255502 261287 255558 261296
rect 255410 260536 255466 260545
rect 255410 260471 255466 260480
rect 255424 260166 255452 260471
rect 255412 260160 255464 260166
rect 255412 260102 255464 260108
rect 256422 260128 256478 260137
rect 256422 260063 256478 260072
rect 255410 259720 255466 259729
rect 255410 259655 255466 259664
rect 255424 259486 255452 259655
rect 255412 259480 255464 259486
rect 255412 259422 255464 259428
rect 255596 259412 255648 259418
rect 255596 259354 255648 259360
rect 255502 259312 255558 259321
rect 255502 259247 255558 259256
rect 255516 258738 255544 259247
rect 255504 258732 255556 258738
rect 255504 258674 255556 258680
rect 255608 258369 255636 259354
rect 255594 258360 255650 258369
rect 255594 258295 255650 258304
rect 255410 257952 255466 257961
rect 255410 257887 255466 257896
rect 255424 256834 255452 257887
rect 255412 256828 255464 256834
rect 255412 256770 255464 256776
rect 255410 256320 255466 256329
rect 255410 256255 255466 256264
rect 255424 255406 255452 256255
rect 255412 255400 255464 255406
rect 255318 255368 255374 255377
rect 254584 255332 254636 255338
rect 255412 255342 255464 255348
rect 255318 255303 255374 255312
rect 255596 255332 255648 255338
rect 254584 255274 254636 255280
rect 254030 253736 254086 253745
rect 254030 253671 254086 253680
rect 253938 252512 253994 252521
rect 253938 252447 253994 252456
rect 252756 248386 252876 248414
rect 252756 222902 252784 248386
rect 252834 242856 252890 242865
rect 252834 242791 252890 242800
rect 252848 236881 252876 242791
rect 252926 242448 252982 242457
rect 252926 242383 252982 242392
rect 252940 242350 252968 242383
rect 252928 242344 252980 242350
rect 252928 242286 252980 242292
rect 253952 237969 253980 252447
rect 254044 239222 254072 253671
rect 254124 247104 254176 247110
rect 254124 247046 254176 247052
rect 254136 240650 254164 247046
rect 254676 246220 254728 246226
rect 254676 246162 254728 246168
rect 254582 241496 254638 241505
rect 254582 241431 254638 241440
rect 254596 240825 254624 241431
rect 254582 240816 254638 240825
rect 254582 240751 254638 240760
rect 254124 240644 254176 240650
rect 254124 240586 254176 240592
rect 254032 239216 254084 239222
rect 254032 239158 254084 239164
rect 253938 237960 253994 237969
rect 253938 237895 253994 237904
rect 252834 236872 252890 236881
rect 252834 236807 252890 236816
rect 253938 235784 253994 235793
rect 253938 235719 253994 235728
rect 253952 233073 253980 235719
rect 253938 233064 253994 233073
rect 253938 232999 253994 233008
rect 253204 224256 253256 224262
rect 253204 224198 253256 224204
rect 252744 222896 252796 222902
rect 252744 222838 252796 222844
rect 252652 220108 252704 220114
rect 252652 220050 252704 220056
rect 252560 120828 252612 120834
rect 252560 120770 252612 120776
rect 252560 112464 252612 112470
rect 252560 112406 252612 112412
rect 251272 49020 251324 49026
rect 251272 48962 251324 48968
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 251284 3482 251312 48962
rect 252572 6914 252600 112406
rect 253216 80714 253244 224198
rect 254596 89593 254624 240751
rect 254688 228993 254716 246162
rect 254674 228984 254730 228993
rect 254674 228919 254730 228928
rect 255332 225593 255360 255303
rect 255596 255274 255648 255280
rect 255502 254960 255558 254969
rect 255502 254895 255558 254904
rect 255412 254584 255464 254590
rect 255410 254552 255412 254561
rect 255464 254552 255466 254561
rect 255410 254487 255466 254496
rect 255516 253978 255544 254895
rect 255504 253972 255556 253978
rect 255504 253914 255556 253920
rect 255410 253328 255466 253337
rect 255410 253263 255466 253272
rect 255424 253230 255452 253263
rect 255412 253224 255464 253230
rect 255412 253166 255464 253172
rect 255410 251968 255466 251977
rect 255410 251903 255466 251912
rect 255504 251932 255556 251938
rect 255424 251870 255452 251903
rect 255504 251874 255556 251880
rect 255412 251864 255464 251870
rect 255412 251806 255464 251812
rect 255516 251569 255544 251874
rect 255502 251560 255558 251569
rect 255502 251495 255558 251504
rect 255502 251152 255558 251161
rect 255502 251087 255558 251096
rect 255410 250744 255466 250753
rect 255410 250679 255466 250688
rect 255424 249937 255452 250679
rect 255410 249928 255466 249937
rect 255410 249863 255466 249872
rect 255516 249830 255544 251087
rect 255504 249824 255556 249830
rect 255608 249801 255636 255274
rect 256436 253201 256464 260063
rect 256422 253192 256478 253201
rect 256422 253127 256478 253136
rect 255504 249766 255556 249772
rect 255594 249792 255650 249801
rect 255594 249727 255650 249736
rect 255502 249384 255558 249393
rect 255502 249319 255558 249328
rect 255410 248976 255466 248985
rect 255410 248911 255466 248920
rect 255424 248538 255452 248911
rect 255412 248532 255464 248538
rect 255412 248474 255464 248480
rect 255516 248470 255544 249319
rect 255504 248464 255556 248470
rect 255410 248432 255466 248441
rect 255504 248406 255556 248412
rect 255410 248367 255466 248376
rect 255424 235793 255452 248367
rect 255502 248160 255558 248169
rect 255502 248095 255558 248104
rect 255516 247722 255544 248095
rect 255504 247716 255556 247722
rect 255504 247658 255556 247664
rect 255502 247208 255558 247217
rect 255502 247143 255558 247152
rect 255516 246265 255544 247143
rect 255686 246800 255742 246809
rect 255686 246735 255742 246744
rect 255502 246256 255558 246265
rect 255502 246191 255558 246200
rect 255594 245984 255650 245993
rect 255594 245919 255650 245928
rect 255504 245608 255556 245614
rect 255502 245576 255504 245585
rect 255556 245576 255558 245585
rect 255502 245511 255558 245520
rect 255608 244934 255636 245919
rect 255700 245682 255728 246735
rect 255688 245676 255740 245682
rect 255688 245618 255740 245624
rect 255686 245168 255742 245177
rect 255686 245103 255742 245112
rect 255596 244928 255648 244934
rect 255596 244870 255648 244876
rect 255594 244760 255650 244769
rect 255594 244695 255650 244704
rect 255502 244216 255558 244225
rect 255502 244151 255558 244160
rect 255516 243574 255544 244151
rect 255504 243568 255556 243574
rect 255608 243545 255636 244695
rect 255504 243510 255556 243516
rect 255594 243536 255650 243545
rect 255594 243471 255650 243480
rect 255700 242894 255728 245103
rect 255778 243672 255834 243681
rect 255778 243607 255834 243616
rect 255688 242888 255740 242894
rect 255688 242830 255740 242836
rect 255504 242208 255556 242214
rect 255504 242150 255556 242156
rect 255594 242176 255650 242185
rect 255516 241777 255544 242150
rect 255594 242111 255650 242120
rect 255502 241768 255558 241777
rect 255502 241703 255558 241712
rect 255608 241466 255636 242111
rect 255792 241505 255820 243607
rect 255778 241496 255834 241505
rect 255596 241460 255648 241466
rect 255778 241431 255834 241440
rect 255596 241402 255648 241408
rect 255410 235784 255466 235793
rect 255410 235719 255466 235728
rect 256056 226840 256108 226846
rect 256056 226782 256108 226788
rect 256068 226370 256096 226782
rect 256056 226364 256108 226370
rect 256056 226306 256108 226312
rect 255318 225584 255374 225593
rect 255318 225519 255374 225528
rect 256068 220114 256096 226306
rect 256056 220108 256108 220114
rect 256056 220050 256108 220056
rect 256608 218748 256660 218754
rect 256608 218690 256660 218696
rect 255964 204944 256016 204950
rect 255964 204886 256016 204892
rect 255320 175296 255372 175302
rect 255320 175238 255372 175244
rect 255332 174593 255360 175238
rect 255318 174584 255374 174593
rect 255318 174519 255374 174528
rect 255320 137284 255372 137290
rect 255320 137226 255372 137232
rect 254582 89584 254638 89593
rect 254582 89519 254638 89528
rect 254596 89010 254624 89519
rect 254584 89004 254636 89010
rect 254584 88946 254636 88952
rect 253204 80708 253256 80714
rect 253204 80650 253256 80656
rect 253216 14482 253244 80650
rect 255332 16574 255360 137226
rect 255976 104174 256004 204886
rect 256620 175302 256648 218690
rect 256712 198694 256740 286039
rect 256790 269104 256846 269113
rect 256790 269039 256846 269048
rect 256804 234598 256832 269039
rect 256882 257544 256938 257553
rect 256882 257479 256938 257488
rect 256792 234592 256844 234598
rect 256792 234534 256844 234540
rect 256896 233209 256924 257479
rect 257526 246392 257582 246401
rect 257526 246327 257582 246336
rect 257540 238105 257568 246327
rect 258184 243506 258212 290799
rect 258276 275505 258304 304778
rect 258356 304292 258408 304298
rect 258356 304234 258408 304240
rect 258368 286346 258396 304234
rect 258736 302190 258764 305050
rect 258724 302184 258776 302190
rect 258724 302126 258776 302132
rect 258724 300960 258776 300966
rect 258724 300902 258776 300908
rect 258736 300150 258764 300902
rect 258724 300144 258776 300150
rect 258724 300086 258776 300092
rect 258538 299976 258594 299985
rect 258538 299911 258594 299920
rect 258552 296002 258580 299911
rect 258540 295996 258592 296002
rect 258540 295938 258592 295944
rect 258814 293856 258870 293865
rect 258814 293791 258870 293800
rect 258828 293282 258856 293791
rect 258816 293276 258868 293282
rect 258816 293218 258868 293224
rect 258632 292188 258684 292194
rect 258632 292130 258684 292136
rect 258356 286340 258408 286346
rect 258356 286282 258408 286288
rect 258446 278216 258502 278225
rect 258446 278151 258502 278160
rect 258262 275496 258318 275505
rect 258262 275431 258318 275440
rect 258356 266416 258408 266422
rect 258356 266358 258408 266364
rect 258368 246226 258396 266358
rect 258356 246220 258408 246226
rect 258356 246162 258408 246168
rect 258172 243500 258224 243506
rect 258172 243442 258224 243448
rect 258356 242888 258408 242894
rect 258356 242830 258408 242836
rect 257526 238096 257582 238105
rect 257526 238031 257582 238040
rect 257342 237416 257398 237425
rect 257342 237351 257398 237360
rect 256882 233200 256938 233209
rect 256882 233135 256938 233144
rect 257356 210458 257384 237351
rect 258262 236056 258318 236065
rect 258262 235991 258318 236000
rect 258276 222193 258304 235991
rect 258368 229770 258396 242830
rect 258460 237425 258488 278151
rect 258540 244928 258592 244934
rect 258540 244870 258592 244876
rect 258446 237416 258502 237425
rect 258446 237351 258502 237360
rect 258356 229764 258408 229770
rect 258356 229706 258408 229712
rect 258262 222184 258318 222193
rect 258262 222119 258318 222128
rect 258552 218754 258580 244870
rect 258540 218748 258592 218754
rect 258540 218690 258592 218696
rect 258644 212566 258672 292130
rect 259276 282192 259328 282198
rect 259276 282134 259328 282140
rect 259288 281081 259316 282134
rect 259368 281988 259420 281994
rect 259368 281930 259420 281936
rect 259380 281625 259408 281930
rect 259366 281616 259422 281625
rect 259366 281551 259422 281560
rect 259274 281072 259330 281081
rect 259274 281007 259330 281016
rect 259472 279449 259500 330482
rect 260840 326460 260892 326466
rect 260840 326402 260892 326408
rect 259552 309868 259604 309874
rect 259552 309810 259604 309816
rect 259458 279440 259514 279449
rect 259458 279375 259514 279384
rect 259458 278080 259514 278089
rect 259458 278015 259514 278024
rect 259472 273222 259500 278015
rect 259564 274310 259592 309810
rect 259736 306400 259788 306406
rect 259736 306342 259788 306348
rect 259642 292224 259698 292233
rect 259642 292159 259698 292168
rect 259552 274304 259604 274310
rect 259552 274246 259604 274252
rect 259460 273216 259512 273222
rect 259460 273158 259512 273164
rect 259368 271176 259420 271182
rect 259368 271118 259420 271124
rect 259380 270298 259408 271118
rect 259368 270292 259420 270298
rect 259368 270234 259420 270240
rect 259368 269136 259420 269142
rect 259368 269078 259420 269084
rect 259380 268705 259408 269078
rect 259366 268696 259422 268705
rect 259366 268631 259422 268640
rect 259564 258074 259592 274246
rect 259472 258046 259592 258074
rect 259276 242888 259328 242894
rect 259276 242830 259328 242836
rect 259288 242282 259316 242830
rect 259276 242276 259328 242282
rect 259276 242218 259328 242224
rect 258724 215960 258776 215966
rect 258724 215902 258776 215908
rect 258080 212560 258132 212566
rect 258080 212502 258132 212508
rect 258632 212560 258684 212566
rect 258632 212502 258684 212508
rect 257344 210452 257396 210458
rect 257344 210394 257396 210400
rect 256700 198688 256752 198694
rect 256700 198630 256752 198636
rect 256608 175296 256660 175302
rect 256608 175238 256660 175244
rect 256712 171834 256740 198630
rect 256700 171828 256752 171834
rect 256700 171770 256752 171776
rect 256056 149184 256108 149190
rect 256056 149126 256108 149132
rect 256068 135930 256096 149126
rect 256148 146396 256200 146402
rect 256148 146338 256200 146344
rect 256160 137290 256188 146338
rect 256148 137284 256200 137290
rect 256148 137226 256200 137232
rect 256056 135924 256108 135930
rect 256056 135866 256108 135872
rect 255964 104168 256016 104174
rect 255964 104110 256016 104116
rect 258092 94761 258120 212502
rect 258736 204377 258764 215902
rect 258170 204368 258226 204377
rect 258170 204303 258226 204312
rect 258722 204368 258778 204377
rect 258722 204303 258778 204312
rect 258078 94752 258134 94761
rect 258078 94687 258134 94696
rect 258184 91089 258212 204303
rect 259472 170406 259500 258046
rect 259552 247716 259604 247722
rect 259552 247658 259604 247664
rect 259564 238754 259592 247658
rect 259656 247110 259684 292159
rect 259748 283422 259776 306342
rect 260852 295225 260880 326402
rect 262220 323604 262272 323610
rect 262220 323546 262272 323552
rect 261024 320204 261076 320210
rect 261024 320146 261076 320152
rect 260932 313948 260984 313954
rect 260932 313890 260984 313896
rect 260838 295216 260894 295225
rect 260838 295151 260894 295160
rect 260748 293140 260800 293146
rect 260748 293082 260800 293088
rect 260760 291825 260788 293082
rect 260746 291816 260802 291825
rect 260746 291751 260802 291760
rect 260748 289808 260800 289814
rect 260746 289776 260748 289785
rect 260800 289776 260802 289785
rect 260746 289711 260802 289720
rect 260840 286340 260892 286346
rect 260840 286282 260892 286288
rect 259736 283416 259788 283422
rect 259736 283358 259788 283364
rect 259826 279848 259882 279857
rect 259826 279783 259882 279792
rect 259736 263628 259788 263634
rect 259736 263570 259788 263576
rect 259644 247104 259696 247110
rect 259644 247046 259696 247052
rect 259564 238726 259684 238754
rect 259552 235952 259604 235958
rect 259552 235894 259604 235900
rect 259460 170400 259512 170406
rect 259460 170342 259512 170348
rect 259564 156097 259592 235894
rect 259656 226846 259684 238726
rect 259748 236706 259776 263570
rect 259736 236700 259788 236706
rect 259736 236642 259788 236648
rect 259840 235958 259868 279783
rect 259828 235952 259880 235958
rect 259828 235894 259880 235900
rect 259644 226840 259696 226846
rect 259644 226782 259696 226788
rect 260852 164898 260880 286282
rect 260944 285666 260972 313890
rect 261036 291854 261064 320146
rect 261484 298172 261536 298178
rect 261484 298114 261536 298120
rect 261496 293894 261524 298114
rect 262232 293962 262260 323546
rect 262312 302320 262364 302326
rect 262312 302262 262364 302268
rect 261576 293956 261628 293962
rect 261576 293898 261628 293904
rect 262220 293956 262272 293962
rect 262220 293898 262272 293904
rect 261484 293888 261536 293894
rect 261484 293830 261536 293836
rect 261024 291848 261076 291854
rect 261024 291790 261076 291796
rect 260932 285660 260984 285666
rect 260932 285602 260984 285608
rect 261024 269816 261076 269822
rect 261024 269758 261076 269764
rect 261036 269210 261064 269758
rect 261024 269204 261076 269210
rect 261024 269146 261076 269152
rect 260930 266520 260986 266529
rect 260930 266455 260986 266464
rect 260944 235929 260972 266455
rect 261036 238746 261064 269146
rect 261496 239426 261524 293830
rect 261588 271862 261616 293898
rect 262218 291680 262274 291689
rect 262218 291615 262274 291624
rect 261576 271856 261628 271862
rect 261576 271798 261628 271804
rect 261484 239420 261536 239426
rect 261484 239362 261536 239368
rect 261024 238740 261076 238746
rect 261024 238682 261076 238688
rect 260930 235920 260986 235929
rect 260930 235855 260986 235864
rect 260930 205728 260986 205737
rect 260930 205663 260932 205672
rect 260984 205663 260986 205672
rect 260932 205634 260984 205640
rect 260840 164892 260892 164898
rect 260840 164834 260892 164840
rect 259550 156088 259606 156097
rect 259550 156023 259606 156032
rect 259368 145580 259420 145586
rect 259368 145522 259420 145528
rect 259380 143546 259408 145522
rect 259368 143540 259420 143546
rect 259368 143482 259420 143488
rect 259380 142866 259408 143482
rect 259368 142860 259420 142866
rect 259368 142802 259420 142808
rect 259564 142154 259592 156023
rect 260104 143540 260156 143546
rect 260104 143482 260156 143488
rect 259472 142126 259592 142154
rect 259472 129033 259500 142126
rect 259458 129024 259514 129033
rect 259458 128959 259514 128968
rect 258170 91080 258226 91089
rect 258170 91015 258226 91024
rect 258724 90364 258776 90370
rect 258724 90306 258776 90312
rect 258736 73234 258764 90306
rect 259460 83496 259512 83502
rect 259460 83438 259512 83444
rect 258724 73228 258776 73234
rect 258724 73170 258776 73176
rect 255332 16546 255912 16574
rect 253204 14476 253256 14482
rect 253204 14418 253256 14424
rect 252572 6886 253520 6914
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253492 480 253520 6886
rect 254674 4856 254730 4865
rect 254674 4791 254730 4800
rect 254688 480 254716 4791
rect 255884 480 255912 16546
rect 256700 15904 256752 15910
rect 256700 15846 256752 15852
rect 256712 490 256740 15846
rect 258736 8974 258764 73170
rect 258264 8968 258316 8974
rect 258264 8910 258316 8916
rect 258724 8968 258776 8974
rect 258724 8910 258776 8916
rect 256896 598 257108 626
rect 256896 490 256924 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 462 256924 490
rect 257080 480 257108 598
rect 258276 480 258304 8910
rect 259472 480 259500 83438
rect 260116 77994 260144 143482
rect 260944 89729 260972 205634
rect 262232 144226 262260 291615
rect 262324 232626 262352 302262
rect 262416 285025 262444 354010
rect 263784 321632 263836 321638
rect 263784 321574 263836 321580
rect 263600 316736 263652 316742
rect 263600 316678 263652 316684
rect 262496 312588 262548 312594
rect 262496 312530 262548 312536
rect 262508 289746 262536 312530
rect 262680 304292 262732 304298
rect 262680 304234 262732 304240
rect 262692 302326 262720 304234
rect 262680 302320 262732 302326
rect 262680 302262 262732 302268
rect 262496 289740 262548 289746
rect 262496 289682 262548 289688
rect 262402 285016 262458 285025
rect 262402 284951 262458 284960
rect 262416 284345 262444 284951
rect 262402 284336 262458 284345
rect 262402 284271 262458 284280
rect 263612 282878 263640 316678
rect 263692 314696 263744 314702
rect 263692 314638 263744 314644
rect 263600 282872 263652 282878
rect 263600 282814 263652 282820
rect 263704 281450 263732 314638
rect 263796 288318 263824 321574
rect 263784 288312 263836 288318
rect 263784 288254 263836 288260
rect 263966 284336 264022 284345
rect 263966 284271 264022 284280
rect 263692 281444 263744 281450
rect 263692 281386 263744 281392
rect 263600 280220 263652 280226
rect 263600 280162 263652 280168
rect 263612 278662 263640 280162
rect 263600 278656 263652 278662
rect 263600 278598 263652 278604
rect 262402 271552 262458 271561
rect 262402 271487 262458 271496
rect 262416 271153 262444 271487
rect 262402 271144 262458 271153
rect 262402 271079 262458 271088
rect 262312 232620 262364 232626
rect 262312 232562 262364 232568
rect 262416 230450 262444 271079
rect 263784 264104 263836 264110
rect 263784 264046 263836 264052
rect 263690 262984 263746 262993
rect 263690 262919 263746 262928
rect 263598 260128 263654 260137
rect 263598 260063 263654 260072
rect 263612 259486 263640 260063
rect 263600 259480 263652 259486
rect 263600 259422 263652 259428
rect 262770 257136 262826 257145
rect 262770 257071 262826 257080
rect 262784 256834 262812 257071
rect 262588 256828 262640 256834
rect 262588 256770 262640 256776
rect 262772 256828 262824 256834
rect 262772 256770 262824 256776
rect 262494 253328 262550 253337
rect 262494 253263 262550 253272
rect 262508 253230 262536 253263
rect 262496 253224 262548 253230
rect 262496 253166 262548 253172
rect 262600 238754 262628 256770
rect 263506 254280 263562 254289
rect 263506 254215 263562 254224
rect 263520 253858 263548 254215
rect 263612 254017 263640 259422
rect 263598 254008 263654 254017
rect 263598 253943 263654 253952
rect 263520 253830 263640 253858
rect 263612 246401 263640 253830
rect 263598 246392 263654 246401
rect 263598 246327 263654 246336
rect 262508 238726 262628 238754
rect 262404 230444 262456 230450
rect 262404 230386 262456 230392
rect 262312 168496 262364 168502
rect 262312 168438 262364 168444
rect 262220 144220 262272 144226
rect 262220 144162 262272 144168
rect 260930 89720 260986 89729
rect 260930 89655 260986 89664
rect 262218 79384 262274 79393
rect 262218 79319 262274 79328
rect 260104 77988 260156 77994
rect 260104 77930 260156 77936
rect 260840 49088 260892 49094
rect 260840 49030 260892 49036
rect 260852 16574 260880 49030
rect 260852 16546 261800 16574
rect 260656 3324 260708 3330
rect 260656 3266 260708 3272
rect 260668 480 260696 3266
rect 261772 480 261800 16546
rect 262232 626 262260 79319
rect 262324 3330 262352 168438
rect 262416 116686 262444 230386
rect 262508 226234 262536 238726
rect 262496 226228 262548 226234
rect 262496 226170 262548 226176
rect 263704 220794 263732 262919
rect 263796 228410 263824 264046
rect 263874 246256 263930 246265
rect 263874 246191 263930 246200
rect 263784 228404 263836 228410
rect 263784 228346 263836 228352
rect 263888 224233 263916 246191
rect 263874 224224 263930 224233
rect 263874 224159 263930 224168
rect 263692 220788 263744 220794
rect 263692 220730 263744 220736
rect 263600 208412 263652 208418
rect 263600 208354 263652 208360
rect 262680 169040 262732 169046
rect 262680 168982 262732 168988
rect 262692 168502 262720 168982
rect 262680 168496 262732 168502
rect 262680 168438 262732 168444
rect 262404 116680 262456 116686
rect 262404 116622 262456 116628
rect 262864 98728 262916 98734
rect 262864 98670 262916 98676
rect 262876 85474 262904 98670
rect 263612 97306 263640 208354
rect 263704 108322 263732 220730
rect 263980 208418 264008 284271
rect 264256 280226 264284 378082
rect 264900 330546 264928 420174
rect 264888 330540 264940 330546
rect 264888 330482 264940 330488
rect 264992 318073 265020 542438
rect 265084 471374 265112 552638
rect 265072 471368 265124 471374
rect 265072 471310 265124 471316
rect 265716 468580 265768 468586
rect 265716 468522 265768 468528
rect 265622 454200 265678 454209
rect 265622 454135 265678 454144
rect 265072 449268 265124 449274
rect 265072 449210 265124 449216
rect 265084 407862 265112 449210
rect 265164 416832 265216 416838
rect 265164 416774 265216 416780
rect 265072 407856 265124 407862
rect 265072 407798 265124 407804
rect 265176 383625 265204 416774
rect 265636 398138 265664 454135
rect 265728 453354 265756 468522
rect 265716 453348 265768 453354
rect 265716 453290 265768 453296
rect 265624 398132 265676 398138
rect 265624 398074 265676 398080
rect 265162 383616 265218 383625
rect 265162 383551 265218 383560
rect 265176 382401 265204 383551
rect 265162 382392 265218 382401
rect 265162 382327 265218 382336
rect 265072 380180 265124 380186
rect 265072 380122 265124 380128
rect 264978 318064 265034 318073
rect 264978 317999 265034 318008
rect 264980 316056 265032 316062
rect 264980 315998 265032 316004
rect 264992 283529 265020 315998
rect 264978 283520 265034 283529
rect 264978 283455 265034 283464
rect 265084 280809 265112 380122
rect 266372 336025 266400 583714
rect 268396 583098 268424 703054
rect 269120 703044 269172 703050
rect 269120 702986 269172 702992
rect 280804 703044 280856 703050
rect 280804 702986 280856 702992
rect 268384 583092 268436 583098
rect 268384 583034 268436 583040
rect 267740 576904 267792 576910
rect 267740 576846 267792 576852
rect 266452 560312 266504 560318
rect 266452 560254 266504 560260
rect 266358 336016 266414 336025
rect 266358 335951 266414 335960
rect 265254 322144 265310 322153
rect 265254 322079 265310 322088
rect 265070 280800 265126 280809
rect 265070 280735 265126 280744
rect 264244 280220 264296 280226
rect 264244 280162 264296 280168
rect 264978 279440 265034 279449
rect 264978 279375 265034 279384
rect 264334 278896 264390 278905
rect 264334 278831 264390 278840
rect 264348 264110 264376 278831
rect 264336 264104 264388 264110
rect 264336 264046 264388 264052
rect 264992 216646 265020 279375
rect 265084 277394 265112 280735
rect 265084 277366 265204 277394
rect 265072 265668 265124 265674
rect 265072 265610 265124 265616
rect 264980 216640 265032 216646
rect 264980 216582 265032 216588
rect 263968 208412 264020 208418
rect 263968 208354 264020 208360
rect 263692 108316 263744 108322
rect 263692 108258 263744 108264
rect 263600 97300 263652 97306
rect 263600 97242 263652 97248
rect 264992 96626 265020 216582
rect 265084 204950 265112 265610
rect 265176 222154 265204 277366
rect 265268 267209 265296 322079
rect 266464 319433 266492 560254
rect 266544 532092 266596 532098
rect 266544 532034 266596 532040
rect 266556 387734 266584 532034
rect 266636 432676 266688 432682
rect 266636 432618 266688 432624
rect 266544 387728 266596 387734
rect 266544 387670 266596 387676
rect 266544 378820 266596 378826
rect 266544 378762 266596 378768
rect 266450 319424 266506 319433
rect 266450 319359 266506 319368
rect 266450 316160 266506 316169
rect 266450 316095 266506 316104
rect 266360 302184 266412 302190
rect 266360 302126 266412 302132
rect 265254 267200 265310 267209
rect 265254 267135 265310 267144
rect 265624 267028 265676 267034
rect 265624 266970 265676 266976
rect 265636 265713 265664 266970
rect 265254 265704 265310 265713
rect 265254 265639 265310 265648
rect 265622 265704 265678 265713
rect 265622 265639 265678 265648
rect 265268 235890 265296 265639
rect 265256 235884 265308 235890
rect 265256 235826 265308 235832
rect 265164 222148 265216 222154
rect 265164 222090 265216 222096
rect 265072 204944 265124 204950
rect 265072 204886 265124 204892
rect 266372 140894 266400 302126
rect 266464 282713 266492 316095
rect 266556 284889 266584 378762
rect 266648 373318 266676 432618
rect 266728 387728 266780 387734
rect 266728 387670 266780 387676
rect 266740 387122 266768 387670
rect 266728 387116 266780 387122
rect 266728 387058 266780 387064
rect 266636 373312 266688 373318
rect 266636 373254 266688 373260
rect 266636 363656 266688 363662
rect 266636 363598 266688 363604
rect 266648 362914 266676 363598
rect 266636 362908 266688 362914
rect 266636 362850 266688 362856
rect 266648 361729 266676 362850
rect 266634 361720 266690 361729
rect 266634 361655 266690 361664
rect 267752 347070 267780 576846
rect 267924 568676 267976 568682
rect 267924 568618 267976 568624
rect 267832 542428 267884 542434
rect 267832 542370 267884 542376
rect 267844 389230 267872 542370
rect 267936 507142 267964 568618
rect 269132 549914 269160 702986
rect 278044 607232 278096 607238
rect 278044 607174 278096 607180
rect 271880 604512 271932 604518
rect 271880 604454 271932 604460
rect 270500 574116 270552 574122
rect 270500 574058 270552 574064
rect 269212 559020 269264 559026
rect 269212 558962 269264 558968
rect 269120 549908 269172 549914
rect 269120 549850 269172 549856
rect 267924 507136 267976 507142
rect 267924 507078 267976 507084
rect 267922 449984 267978 449993
rect 267922 449919 267978 449928
rect 267832 389224 267884 389230
rect 267832 389166 267884 389172
rect 267740 347064 267792 347070
rect 267740 347006 267792 347012
rect 267740 344344 267792 344350
rect 267740 344286 267792 344292
rect 266634 301064 266690 301073
rect 266634 300999 266690 301008
rect 266542 284880 266598 284889
rect 266542 284815 266598 284824
rect 266556 284374 266584 284815
rect 266544 284368 266596 284374
rect 266544 284310 266596 284316
rect 266450 282704 266506 282713
rect 266450 282639 266506 282648
rect 266542 263120 266598 263129
rect 266542 263055 266598 263064
rect 266452 260840 266504 260846
rect 266452 260782 266504 260788
rect 266464 260166 266492 260782
rect 266452 260160 266504 260166
rect 266452 260102 266504 260108
rect 266464 259729 266492 260102
rect 266450 259720 266506 259729
rect 266450 259655 266506 259664
rect 266452 258732 266504 258738
rect 266452 258674 266504 258680
rect 266464 258097 266492 258674
rect 266450 258088 266506 258097
rect 266450 258023 266506 258032
rect 266450 251968 266506 251977
rect 266450 251903 266452 251912
rect 266504 251903 266506 251912
rect 266452 251874 266504 251880
rect 266556 234530 266584 263055
rect 266648 240786 266676 300999
rect 267752 295322 267780 344286
rect 267830 320104 267886 320113
rect 267830 320039 267886 320048
rect 267844 309777 267872 320039
rect 267936 319462 267964 449919
rect 268384 398812 268436 398818
rect 268384 398754 268436 398760
rect 268396 376689 268424 398754
rect 268382 376680 268438 376689
rect 268382 376615 268438 376624
rect 269224 355366 269252 558962
rect 269488 553512 269540 553518
rect 269488 553454 269540 553460
rect 269394 461000 269450 461009
rect 269394 460935 269450 460944
rect 269304 442944 269356 442950
rect 269304 442886 269356 442892
rect 269316 442270 269344 442886
rect 269304 442264 269356 442270
rect 269304 442206 269356 442212
rect 269212 355360 269264 355366
rect 269212 355302 269264 355308
rect 269316 325694 269344 442206
rect 269408 371890 269436 460935
rect 269396 371884 269448 371890
rect 269396 371826 269448 371832
rect 269396 342304 269448 342310
rect 269396 342246 269448 342252
rect 269224 325666 269344 325694
rect 269224 322969 269252 325666
rect 269210 322960 269266 322969
rect 269210 322895 269266 322904
rect 267924 319456 267976 319462
rect 267922 319424 267924 319433
rect 267976 319424 267978 319433
rect 267922 319359 267978 319368
rect 267830 309768 267886 309777
rect 267830 309703 267886 309712
rect 267832 307080 267884 307086
rect 267832 307022 267884 307028
rect 267740 295316 267792 295322
rect 267740 295258 267792 295264
rect 267738 286512 267794 286521
rect 267738 286447 267794 286456
rect 266728 284368 266780 284374
rect 266728 284310 266780 284316
rect 266636 240780 266688 240786
rect 266636 240722 266688 240728
rect 266544 234524 266596 234530
rect 266544 234466 266596 234472
rect 266740 214577 266768 284310
rect 266726 214568 266782 214577
rect 266726 214503 266782 214512
rect 266740 200114 266768 214503
rect 266464 200086 266768 200114
rect 266360 140888 266412 140894
rect 266360 140830 266412 140836
rect 266464 102134 266492 200086
rect 267004 140888 267056 140894
rect 267004 140830 267056 140836
rect 266452 102128 266504 102134
rect 266452 102070 266504 102076
rect 264980 96620 265032 96626
rect 264980 96562 265032 96568
rect 264242 95840 264298 95849
rect 264242 95775 264298 95784
rect 262864 85468 262916 85474
rect 262864 85410 262916 85416
rect 264256 78674 264284 95775
rect 263600 78668 263652 78674
rect 263600 78610 263652 78616
rect 264244 78668 264296 78674
rect 264244 78610 264296 78616
rect 263612 16574 263640 78610
rect 266360 29640 266412 29646
rect 266360 29582 266412 29588
rect 266372 16574 266400 29582
rect 263612 16546 264192 16574
rect 266372 16546 266584 16574
rect 262312 3324 262364 3330
rect 262312 3266 262364 3272
rect 262232 598 262536 626
rect 262508 490 262536 598
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 265346 3360 265402 3369
rect 265346 3295 265402 3304
rect 265360 480 265388 3295
rect 266556 480 266584 16546
rect 267016 4146 267044 140830
rect 267752 131034 267780 286447
rect 267844 282198 267872 307022
rect 269118 303920 269174 303929
rect 269118 303855 269174 303864
rect 268108 302252 268160 302258
rect 268108 302194 268160 302200
rect 267924 296744 267976 296750
rect 267924 296686 267976 296692
rect 267832 282192 267884 282198
rect 267832 282134 267884 282140
rect 267832 269068 267884 269074
rect 267832 269010 267884 269016
rect 267844 267782 267872 269010
rect 267832 267776 267884 267782
rect 267832 267718 267884 267724
rect 267844 149054 267872 267718
rect 267936 231130 267964 296686
rect 268014 295216 268070 295225
rect 268014 295151 268070 295160
rect 268028 232558 268056 295151
rect 268120 288425 268148 302194
rect 268106 288416 268162 288425
rect 268106 288351 268162 288360
rect 268108 241460 268160 241466
rect 268108 241402 268160 241408
rect 268120 240553 268148 241402
rect 268106 240544 268162 240553
rect 268106 240479 268162 240488
rect 268016 232552 268068 232558
rect 268016 232494 268068 232500
rect 267924 231124 267976 231130
rect 267924 231066 267976 231072
rect 268384 230036 268436 230042
rect 268384 229978 268436 229984
rect 268396 200802 268424 229978
rect 268384 200796 268436 200802
rect 268384 200738 268436 200744
rect 267832 149048 267884 149054
rect 267832 148990 267884 148996
rect 267740 131028 267792 131034
rect 267740 130970 267792 130976
rect 267832 127696 267884 127702
rect 267832 127638 267884 127644
rect 267844 16574 267872 127638
rect 269132 112470 269160 303855
rect 269224 289814 269252 322895
rect 269212 289808 269264 289814
rect 269212 289750 269264 289756
rect 269210 288416 269266 288425
rect 269210 288351 269266 288360
rect 269224 159390 269252 288351
rect 269408 280158 269436 342246
rect 269500 312497 269528 553454
rect 270512 463010 270540 574058
rect 270592 532024 270644 532030
rect 270592 531966 270644 531972
rect 270604 473414 270632 531966
rect 270592 473408 270644 473414
rect 270592 473350 270644 473356
rect 270500 463004 270552 463010
rect 270500 462946 270552 462952
rect 270500 458856 270552 458862
rect 270500 458798 270552 458804
rect 269764 455456 269816 455462
rect 269764 455398 269816 455404
rect 269776 441697 269804 455398
rect 269762 441688 269818 441697
rect 269762 441623 269818 441632
rect 270408 371272 270460 371278
rect 270408 371214 270460 371220
rect 269486 312488 269542 312497
rect 269486 312423 269542 312432
rect 269396 280152 269448 280158
rect 269396 280094 269448 280100
rect 269302 269240 269358 269249
rect 269302 269175 269358 269184
rect 269316 207058 269344 269175
rect 270420 266422 270448 371214
rect 270512 307737 270540 458798
rect 270604 443018 270632 473350
rect 270868 454708 270920 454714
rect 270868 454650 270920 454656
rect 270682 451616 270738 451625
rect 270682 451551 270738 451560
rect 270592 443012 270644 443018
rect 270592 442954 270644 442960
rect 270696 350606 270724 451551
rect 270776 408536 270828 408542
rect 270776 408478 270828 408484
rect 270788 361554 270816 408478
rect 270776 361548 270828 361554
rect 270776 361490 270828 361496
rect 270788 360233 270816 361490
rect 270774 360224 270830 360233
rect 270774 360159 270830 360168
rect 270684 350600 270736 350606
rect 270684 350542 270736 350548
rect 270880 316034 270908 454650
rect 271892 385014 271920 604454
rect 271972 599072 272024 599078
rect 271972 599014 272024 599020
rect 271984 465118 272012 599014
rect 276112 599004 276164 599010
rect 276112 598946 276164 598952
rect 273260 597576 273312 597582
rect 273260 597518 273312 597524
rect 271972 465112 272024 465118
rect 271972 465054 272024 465060
rect 272524 465112 272576 465118
rect 272524 465054 272576 465060
rect 272064 442332 272116 442338
rect 272064 442274 272116 442280
rect 271972 432608 272024 432614
rect 271972 432550 272024 432556
rect 271880 385008 271932 385014
rect 271880 384950 271932 384956
rect 270960 350600 271012 350606
rect 270960 350542 271012 350548
rect 270788 316006 270908 316034
rect 270788 311953 270816 316006
rect 270774 311944 270830 311953
rect 270774 311879 270830 311888
rect 270498 307728 270554 307737
rect 270498 307663 270554 307672
rect 270590 299840 270646 299849
rect 270590 299775 270646 299784
rect 270498 273592 270554 273601
rect 270498 273527 270554 273536
rect 270408 266416 270460 266422
rect 270408 266358 270460 266364
rect 269394 265568 269450 265577
rect 269394 265503 269450 265512
rect 269408 212498 269436 265503
rect 269396 212492 269448 212498
rect 269396 212434 269448 212440
rect 269304 207052 269356 207058
rect 269304 206994 269356 207000
rect 269212 159384 269264 159390
rect 269212 159326 269264 159332
rect 269120 112464 269172 112470
rect 269120 112406 269172 112412
rect 269316 98802 269344 206994
rect 270512 162761 270540 273527
rect 270604 224262 270632 299775
rect 270684 274712 270736 274718
rect 270684 274654 270736 274660
rect 270592 224256 270644 224262
rect 270592 224198 270644 224204
rect 270696 206310 270724 274654
rect 270788 269074 270816 311879
rect 270972 273601 271000 350542
rect 270958 273592 271014 273601
rect 270958 273527 271014 273536
rect 271142 269104 271198 269113
rect 270776 269068 270828 269074
rect 271142 269039 271198 269048
rect 270776 269010 270828 269016
rect 271156 268394 271184 269039
rect 271144 268388 271196 268394
rect 271144 268330 271196 268336
rect 271788 268388 271840 268394
rect 271788 268330 271840 268336
rect 271800 267782 271828 268330
rect 271788 267776 271840 267782
rect 271788 267718 271840 267724
rect 270776 266416 270828 266422
rect 270776 266358 270828 266364
rect 270788 238678 270816 266358
rect 271880 253972 271932 253978
rect 271880 253914 271932 253920
rect 270776 238672 270828 238678
rect 270776 238614 270828 238620
rect 271892 226953 271920 253914
rect 271984 247722 272012 432550
rect 272076 299470 272104 442274
rect 272536 434790 272564 465054
rect 273272 452441 273300 597518
rect 274732 588600 274784 588606
rect 274732 588542 274784 588548
rect 273352 558952 273404 558958
rect 273352 558894 273404 558900
rect 273258 452432 273314 452441
rect 273258 452367 273314 452376
rect 273074 451344 273130 451353
rect 273074 451279 273130 451288
rect 273088 451194 273116 451279
rect 273088 451166 273300 451194
rect 272524 434784 272576 434790
rect 272524 434726 272576 434732
rect 272248 387116 272300 387122
rect 272248 387058 272300 387064
rect 272156 330540 272208 330546
rect 272156 330482 272208 330488
rect 272064 299464 272116 299470
rect 272064 299406 272116 299412
rect 272064 296064 272116 296070
rect 272064 296006 272116 296012
rect 271972 247716 272024 247722
rect 271972 247658 272024 247664
rect 271970 243536 272026 243545
rect 271970 243471 272026 243480
rect 271878 226944 271934 226953
rect 271878 226879 271934 226888
rect 271984 219434 272012 243471
rect 272076 230042 272104 296006
rect 272168 246265 272196 330482
rect 272260 274718 272288 387058
rect 272248 274712 272300 274718
rect 272248 274654 272300 274660
rect 273272 269822 273300 451166
rect 273364 380186 273392 558894
rect 274640 557592 274692 557598
rect 274640 557534 274692 557540
rect 273442 533352 273498 533361
rect 273442 533287 273498 533296
rect 273456 480254 273484 533287
rect 273456 480226 273576 480254
rect 273548 459649 273576 480226
rect 273534 459640 273590 459649
rect 273534 459575 273590 459584
rect 273442 452704 273498 452713
rect 273442 452639 273498 452648
rect 273352 380180 273404 380186
rect 273352 380122 273404 380128
rect 273352 379296 273404 379302
rect 273352 379238 273404 379244
rect 273364 271153 273392 379238
rect 273456 298081 273484 452639
rect 273548 426426 273576 459575
rect 273536 426420 273588 426426
rect 273536 426362 273588 426368
rect 273548 425746 273576 426362
rect 273536 425740 273588 425746
rect 273536 425682 273588 425688
rect 273536 407788 273588 407794
rect 273536 407730 273588 407736
rect 273548 379506 273576 407730
rect 273536 379500 273588 379506
rect 273536 379442 273588 379448
rect 273548 379302 273576 379442
rect 273536 379296 273588 379302
rect 273536 379238 273588 379244
rect 274652 333266 274680 557534
rect 274744 382265 274772 588542
rect 274824 584452 274876 584458
rect 274824 584394 274876 584400
rect 274836 398818 274864 584394
rect 274916 453348 274968 453354
rect 274916 453290 274968 453296
rect 274824 398812 274876 398818
rect 274824 398754 274876 398760
rect 274730 382256 274786 382265
rect 274730 382191 274786 382200
rect 274928 371278 274956 453290
rect 276020 449200 276072 449206
rect 276020 449142 276072 449148
rect 275008 398132 275060 398138
rect 275008 398074 275060 398080
rect 274916 371272 274968 371278
rect 274916 371214 274968 371220
rect 274732 361616 274784 361622
rect 274732 361558 274784 361564
rect 274640 333260 274692 333266
rect 274640 333202 274692 333208
rect 274640 300212 274692 300218
rect 274640 300154 274692 300160
rect 273442 298072 273498 298081
rect 273442 298007 273498 298016
rect 273456 296857 273484 298007
rect 273442 296848 273498 296857
rect 273442 296783 273498 296792
rect 273444 282192 273496 282198
rect 273444 282134 273496 282140
rect 273456 281625 273484 282134
rect 273442 281616 273498 281625
rect 273442 281551 273498 281560
rect 273350 271144 273406 271153
rect 273350 271079 273406 271088
rect 273260 269816 273312 269822
rect 273260 269758 273312 269764
rect 273260 264988 273312 264994
rect 273260 264930 273312 264936
rect 272340 254652 272392 254658
rect 272340 254594 272392 254600
rect 272352 253978 272380 254594
rect 272340 253972 272392 253978
rect 272340 253914 272392 253920
rect 272522 247480 272578 247489
rect 272522 247415 272578 247424
rect 272536 247081 272564 247415
rect 272522 247072 272578 247081
rect 272522 247007 272578 247016
rect 272154 246256 272210 246265
rect 272154 246191 272210 246200
rect 272064 230036 272116 230042
rect 272064 229978 272116 229984
rect 271892 219406 272012 219434
rect 271892 218006 271920 219406
rect 271880 218000 271932 218006
rect 271880 217942 271932 217948
rect 270684 206304 270736 206310
rect 270684 206246 270736 206252
rect 270498 162752 270554 162761
rect 270498 162687 270554 162696
rect 270500 113824 270552 113830
rect 270500 113766 270552 113772
rect 270408 104848 270460 104854
rect 270408 104790 270460 104796
rect 270420 103562 270448 104790
rect 270408 103556 270460 103562
rect 270408 103498 270460 103504
rect 269304 98796 269356 98802
rect 269304 98738 269356 98744
rect 269118 73808 269174 73817
rect 269118 73743 269174 73752
rect 269132 16574 269160 73743
rect 269764 17264 269816 17270
rect 269764 17206 269816 17212
rect 267844 16546 268424 16574
rect 269132 16546 269712 16574
rect 267004 4140 267056 4146
rect 267004 4082 267056 4088
rect 267740 4140 267792 4146
rect 267740 4082 267792 4088
rect 267752 480 267780 4082
rect 268396 490 268424 16546
rect 269684 2938 269712 16546
rect 269776 3126 269804 17206
rect 270420 15910 270448 103498
rect 270512 16574 270540 113766
rect 271892 99346 271920 217942
rect 272536 195974 272564 247007
rect 273272 215966 273300 264930
rect 273260 215960 273312 215966
rect 273260 215902 273312 215908
rect 273456 213217 273484 281551
rect 273534 276720 273590 276729
rect 273534 276655 273590 276664
rect 273442 213208 273498 213217
rect 273442 213143 273498 213152
rect 273456 200114 273484 213143
rect 273272 200086 273484 200114
rect 272524 195968 272576 195974
rect 272524 195910 272576 195916
rect 272536 195294 272564 195910
rect 272524 195288 272576 195294
rect 272524 195230 272576 195236
rect 273272 105602 273300 200086
rect 273548 153785 273576 276655
rect 273534 153776 273590 153785
rect 273534 153711 273590 153720
rect 273260 105596 273312 105602
rect 273260 105538 273312 105544
rect 274652 104854 274680 300154
rect 274744 263566 274772 361558
rect 274824 295316 274876 295322
rect 274824 295258 274876 295264
rect 274732 263560 274784 263566
rect 274732 263502 274784 263508
rect 274730 261080 274786 261089
rect 274730 261015 274786 261024
rect 274744 160818 274772 261015
rect 274836 221474 274864 295258
rect 275020 293865 275048 398074
rect 275006 293856 275062 293865
rect 275006 293791 275062 293800
rect 275020 292641 275048 293791
rect 275006 292632 275062 292641
rect 275006 292567 275062 292576
rect 275282 267200 275338 267209
rect 275282 267135 275338 267144
rect 275296 257009 275324 267135
rect 275282 257000 275338 257009
rect 275282 256935 275338 256944
rect 274916 250504 274968 250510
rect 274916 250446 274968 250452
rect 274928 249830 274956 250446
rect 274916 249824 274968 249830
rect 274916 249766 274968 249772
rect 274928 223582 274956 249766
rect 276032 238649 276060 449142
rect 276124 408542 276152 598946
rect 277492 571464 277544 571470
rect 277492 571406 277544 571412
rect 276204 546508 276256 546514
rect 276204 546450 276256 546456
rect 276112 408536 276164 408542
rect 276112 408478 276164 408484
rect 276112 405748 276164 405754
rect 276112 405690 276164 405696
rect 276124 368490 276152 405690
rect 276216 389162 276244 546450
rect 277400 538348 277452 538354
rect 277400 538290 277452 538296
rect 276296 435396 276348 435402
rect 276296 435338 276348 435344
rect 276204 389156 276256 389162
rect 276204 389098 276256 389104
rect 276112 368484 276164 368490
rect 276112 368426 276164 368432
rect 276124 281518 276152 368426
rect 276308 310554 276336 435338
rect 277412 348401 277440 538290
rect 277504 458833 277532 571406
rect 277584 553444 277636 553450
rect 277584 553386 277636 553392
rect 277490 458824 277546 458833
rect 277490 458759 277546 458768
rect 277596 458182 277624 553386
rect 278056 541686 278084 607174
rect 278780 575544 278832 575550
rect 278780 575486 278832 575492
rect 278044 541680 278096 541686
rect 278044 541622 278096 541628
rect 277676 478168 277728 478174
rect 277676 478110 277728 478116
rect 277584 458176 277636 458182
rect 277584 458118 277636 458124
rect 277492 455524 277544 455530
rect 277492 455466 277544 455472
rect 277398 348392 277454 348401
rect 277398 348327 277454 348336
rect 277398 317520 277454 317529
rect 277398 317455 277454 317464
rect 276296 310548 276348 310554
rect 276296 310490 276348 310496
rect 276202 292632 276258 292641
rect 276202 292567 276258 292576
rect 276112 281512 276164 281518
rect 276112 281454 276164 281460
rect 276112 276072 276164 276078
rect 276112 276014 276164 276020
rect 276018 238640 276074 238649
rect 276018 238575 276074 238584
rect 274916 223576 274968 223582
rect 274916 223518 274968 223524
rect 274824 221468 274876 221474
rect 274824 221410 274876 221416
rect 274732 160812 274784 160818
rect 274732 160754 274784 160760
rect 276020 137284 276072 137290
rect 276020 137226 276072 137232
rect 274640 104848 274692 104854
rect 274640 104790 274692 104796
rect 271880 99340 271932 99346
rect 271880 99282 271932 99288
rect 271892 98734 271920 99282
rect 271880 98728 271932 98734
rect 271880 98670 271932 98676
rect 273258 86184 273314 86193
rect 273258 86119 273314 86128
rect 270512 16546 270816 16574
rect 270408 15904 270460 15910
rect 270408 15846 270460 15852
rect 269764 3120 269816 3126
rect 269764 3062 269816 3068
rect 269684 2910 270080 2938
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 2910
rect 270788 490 270816 16546
rect 272432 3120 272484 3126
rect 272432 3062 272484 3068
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3062
rect 273272 490 273300 86119
rect 274824 8968 274876 8974
rect 274824 8910 274876 8916
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 8910
rect 276032 3602 276060 137226
rect 276124 131102 276152 276014
rect 276216 169046 276244 292567
rect 276308 276690 276336 310490
rect 277412 276729 277440 317455
rect 277398 276720 277454 276729
rect 276296 276684 276348 276690
rect 277398 276655 277454 276664
rect 276296 276626 276348 276632
rect 276308 276078 276336 276626
rect 276296 276072 276348 276078
rect 276296 276014 276348 276020
rect 277504 267034 277532 455466
rect 277688 451274 277716 478110
rect 278792 461650 278820 575486
rect 278872 539640 278924 539646
rect 278872 539582 278924 539588
rect 278780 461644 278832 461650
rect 278780 461586 278832 461592
rect 277766 458824 277822 458833
rect 277766 458759 277822 458768
rect 277596 451246 277716 451274
rect 277596 447098 277624 451246
rect 277584 447092 277636 447098
rect 277584 447034 277636 447040
rect 277676 381540 277728 381546
rect 277676 381482 277728 381488
rect 277582 306504 277638 306513
rect 277582 306439 277638 306448
rect 277492 267028 277544 267034
rect 277492 266970 277544 266976
rect 276294 264344 276350 264353
rect 276294 264279 276350 264288
rect 276308 263673 276336 264279
rect 276294 263664 276350 263673
rect 276294 263599 276350 263608
rect 276308 188358 276336 263599
rect 277400 263560 277452 263566
rect 277400 263502 277452 263508
rect 276296 188352 276348 188358
rect 276296 188294 276348 188300
rect 276204 169040 276256 169046
rect 276204 168982 276256 168988
rect 276112 131096 276164 131102
rect 276112 131038 276164 131044
rect 277412 101454 277440 263502
rect 277490 243672 277546 243681
rect 277490 243607 277546 243616
rect 277504 243574 277532 243607
rect 277492 243568 277544 243574
rect 277492 243510 277544 243516
rect 277596 145586 277624 306439
rect 277688 276010 277716 381482
rect 277780 317529 277808 458759
rect 278778 452840 278834 452849
rect 278778 452775 278834 452784
rect 277766 317520 277822 317529
rect 277766 317455 277822 317464
rect 277676 276004 277728 276010
rect 277676 275946 277728 275952
rect 278318 262168 278374 262177
rect 278318 262103 278374 262112
rect 278332 261526 278360 262103
rect 278320 261520 278372 261526
rect 278320 261462 278372 261468
rect 278332 261361 278360 261462
rect 278318 261352 278374 261361
rect 278318 261287 278374 261296
rect 278044 248532 278096 248538
rect 278044 248474 278096 248480
rect 278056 232558 278084 248474
rect 278792 242282 278820 452775
rect 278884 340105 278912 539582
rect 280816 536722 280844 702986
rect 283852 700330 283880 703520
rect 285588 702840 285640 702846
rect 285588 702782 285640 702788
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 283104 583024 283156 583030
rect 283104 582966 283156 582972
rect 282000 566500 282052 566506
rect 282000 566442 282052 566448
rect 282012 565962 282040 566442
rect 281540 565956 281592 565962
rect 281540 565898 281592 565904
rect 282000 565956 282052 565962
rect 282000 565898 282052 565904
rect 280804 536716 280856 536722
rect 280804 536658 280856 536664
rect 280344 533384 280396 533390
rect 280344 533326 280396 533332
rect 280252 529236 280304 529242
rect 280252 529178 280304 529184
rect 279424 464364 279476 464370
rect 279424 464306 279476 464312
rect 278964 393372 279016 393378
rect 278964 393314 279016 393320
rect 278976 348430 279004 393314
rect 279436 392630 279464 464306
rect 280158 463720 280214 463729
rect 280158 463655 280214 463664
rect 279424 392624 279476 392630
rect 279424 392566 279476 392572
rect 279424 375352 279476 375358
rect 279424 375294 279476 375300
rect 278964 348424 279016 348430
rect 278964 348366 279016 348372
rect 278870 340096 278926 340105
rect 278870 340031 278926 340040
rect 278870 296848 278926 296857
rect 278870 296783 278926 296792
rect 278780 242276 278832 242282
rect 278780 242218 278832 242224
rect 278044 232552 278096 232558
rect 278044 232494 278096 232500
rect 278056 219434 278084 232494
rect 278688 229628 278740 229634
rect 278688 229570 278740 229576
rect 278044 219428 278096 219434
rect 278044 219370 278096 219376
rect 277584 145580 277636 145586
rect 277584 145522 277636 145528
rect 277400 101448 277452 101454
rect 277400 101390 277452 101396
rect 278044 60104 278096 60110
rect 278044 60046 278096 60052
rect 276112 18692 276164 18698
rect 276112 18634 276164 18640
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276124 3482 276152 18634
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 277136 480 277164 3538
rect 278056 3398 278084 60046
rect 278700 57866 278728 229570
rect 278884 159390 278912 296783
rect 278976 277370 279004 348366
rect 278964 277364 279016 277370
rect 278964 277306 279016 277312
rect 279436 260846 279464 375294
rect 279424 260840 279476 260846
rect 279424 260782 279476 260788
rect 278964 255400 279016 255406
rect 278964 255342 279016 255348
rect 278976 209778 279004 255342
rect 280068 246356 280120 246362
rect 280068 246298 280120 246304
rect 280080 245682 280108 246298
rect 279424 245676 279476 245682
rect 279424 245618 279476 245624
rect 280068 245676 280120 245682
rect 280068 245618 280120 245624
rect 278964 209772 279016 209778
rect 278964 209714 279016 209720
rect 278872 159384 278924 159390
rect 278872 159326 278924 159332
rect 279436 124166 279464 245618
rect 280172 235793 280200 463655
rect 280264 387705 280292 529178
rect 280356 391270 280384 533326
rect 281448 418124 281500 418130
rect 281448 418066 281500 418072
rect 281460 417450 281488 418066
rect 280436 417444 280488 417450
rect 280436 417386 280488 417392
rect 281448 417444 281500 417450
rect 281448 417386 281500 417392
rect 280448 416809 280476 417386
rect 280434 416800 280490 416809
rect 280434 416735 280490 416744
rect 280436 400240 280488 400246
rect 280436 400182 280488 400188
rect 280344 391264 280396 391270
rect 280344 391206 280396 391212
rect 280250 387696 280306 387705
rect 280250 387631 280306 387640
rect 280344 383716 280396 383722
rect 280344 383658 280396 383664
rect 280250 369744 280306 369753
rect 280250 369679 280306 369688
rect 280264 254658 280292 369679
rect 280356 278730 280384 383658
rect 280448 352578 280476 400182
rect 281446 387696 281502 387705
rect 281446 387631 281502 387640
rect 281460 387122 281488 387631
rect 281448 387116 281500 387122
rect 281448 387058 281500 387064
rect 281552 380905 281580 565898
rect 282920 565888 282972 565894
rect 282920 565830 282972 565836
rect 281632 469872 281684 469878
rect 281632 469814 281684 469820
rect 281644 438190 281672 469814
rect 281632 438184 281684 438190
rect 281632 438126 281684 438132
rect 281538 380896 281594 380905
rect 281538 380831 281594 380840
rect 281552 375358 281580 380831
rect 281540 375352 281592 375358
rect 281540 375294 281592 375300
rect 280436 352572 280488 352578
rect 280436 352514 280488 352520
rect 280344 278724 280396 278730
rect 280344 278666 280396 278672
rect 280448 271182 280476 352514
rect 280526 325816 280582 325825
rect 280526 325751 280582 325760
rect 280540 325718 280568 325751
rect 280528 325712 280580 325718
rect 280528 325654 280580 325660
rect 281540 321564 281592 321570
rect 281540 321506 281592 321512
rect 281552 321366 281580 321506
rect 281540 321360 281592 321366
rect 281540 321302 281592 321308
rect 281552 288386 281580 321302
rect 281540 288380 281592 288386
rect 281540 288322 281592 288328
rect 281644 286385 281672 438126
rect 281816 422340 281868 422346
rect 281816 422282 281868 422288
rect 281724 382968 281776 382974
rect 281724 382910 281776 382916
rect 281630 286376 281686 286385
rect 281630 286311 281686 286320
rect 281538 283520 281594 283529
rect 281538 283455 281594 283464
rect 280436 271176 280488 271182
rect 280436 271118 280488 271124
rect 280436 267776 280488 267782
rect 280436 267718 280488 267724
rect 280342 256728 280398 256737
rect 280342 256663 280398 256672
rect 280252 254652 280304 254658
rect 280252 254594 280304 254600
rect 280252 243568 280304 243574
rect 280252 243510 280304 243516
rect 280158 235784 280214 235793
rect 280158 235719 280214 235728
rect 280172 235278 280200 235719
rect 280160 235272 280212 235278
rect 280160 235214 280212 235220
rect 280160 225072 280212 225078
rect 280160 225014 280212 225020
rect 279424 124160 279476 124166
rect 279424 124102 279476 124108
rect 280172 115938 280200 225014
rect 280160 115932 280212 115938
rect 280160 115874 280212 115880
rect 280264 86970 280292 243510
rect 280356 198014 280384 256663
rect 280448 226302 280476 267718
rect 280436 226296 280488 226302
rect 280436 226238 280488 226244
rect 280448 225078 280476 226238
rect 280436 225072 280488 225078
rect 280436 225014 280488 225020
rect 280344 198008 280396 198014
rect 280344 197950 280396 197956
rect 280252 86964 280304 86970
rect 280252 86906 280304 86912
rect 280160 79348 280212 79354
rect 280160 79290 280212 79296
rect 278688 57860 278740 57866
rect 278688 57802 278740 57808
rect 278700 57254 278728 57802
rect 278688 57248 278740 57254
rect 278688 57190 278740 57196
rect 278780 37936 278832 37942
rect 278780 37878 278832 37884
rect 278792 16574 278820 37878
rect 280172 16574 280200 79290
rect 281552 68950 281580 283455
rect 281736 274650 281764 382910
rect 281828 321366 281856 422282
rect 281816 321360 281868 321366
rect 281816 321302 281868 321308
rect 282932 313993 282960 565830
rect 283012 447092 283064 447098
rect 283012 447034 283064 447040
rect 282918 313984 282974 313993
rect 282918 313919 282974 313928
rect 281814 304192 281870 304201
rect 281814 304127 281870 304136
rect 281724 274644 281776 274650
rect 281724 274586 281776 274592
rect 281724 271924 281776 271930
rect 281724 271866 281776 271872
rect 281632 252816 281684 252822
rect 281632 252758 281684 252764
rect 281644 251870 281672 252758
rect 281632 251864 281684 251870
rect 281632 251806 281684 251812
rect 281644 126993 281672 251806
rect 281736 152425 281764 271866
rect 281828 203590 281856 304127
rect 282920 300144 282972 300150
rect 282920 300086 282972 300092
rect 282000 272536 282052 272542
rect 282000 272478 282052 272484
rect 282012 271930 282040 272478
rect 282000 271924 282052 271930
rect 282000 271866 282052 271872
rect 281816 203584 281868 203590
rect 281816 203526 281868 203532
rect 281722 152416 281778 152425
rect 281722 152351 281778 152360
rect 281630 126984 281686 126993
rect 281630 126919 281686 126928
rect 282932 102814 282960 300086
rect 283024 241466 283052 447034
rect 283116 386073 283144 582966
rect 284300 573368 284352 573374
rect 284300 573310 284352 573316
rect 283196 425740 283248 425746
rect 283196 425682 283248 425688
rect 283102 386064 283158 386073
rect 283102 385999 283158 386008
rect 283208 279449 283236 425682
rect 283194 279440 283250 279449
rect 283194 279375 283250 279384
rect 283104 256012 283156 256018
rect 283104 255954 283156 255960
rect 283116 255338 283144 255954
rect 283104 255332 283156 255338
rect 283104 255274 283156 255280
rect 283012 241460 283064 241466
rect 283012 241402 283064 241408
rect 283116 163538 283144 255274
rect 284312 244934 284340 573310
rect 284392 568608 284444 568614
rect 284392 568550 284444 568556
rect 284404 390561 284432 568550
rect 285600 536761 285628 702782
rect 289728 604512 289780 604518
rect 288622 604480 288678 604489
rect 288622 604415 288678 604424
rect 289726 604480 289728 604489
rect 289780 604480 289782 604489
rect 289726 604415 289782 604424
rect 285680 601792 285732 601798
rect 285680 601734 285732 601740
rect 285586 536752 285642 536761
rect 285586 536687 285642 536696
rect 285600 536081 285628 536687
rect 285586 536072 285642 536081
rect 285586 536007 285642 536016
rect 284484 472116 284536 472122
rect 284484 472058 284536 472064
rect 284390 390552 284446 390561
rect 284390 390487 284446 390496
rect 284404 389201 284432 390487
rect 284390 389192 284446 389201
rect 284390 389127 284446 389136
rect 284390 385656 284446 385665
rect 284390 385591 284446 385600
rect 284300 244928 284352 244934
rect 284300 244870 284352 244876
rect 284404 242214 284432 385591
rect 284496 365022 284524 472058
rect 285692 419490 285720 601734
rect 287060 595468 287112 595474
rect 287060 595410 287112 595416
rect 286324 571396 286376 571402
rect 286324 571338 286376 571344
rect 285956 436756 286008 436762
rect 285956 436698 286008 436704
rect 285772 427100 285824 427106
rect 285772 427042 285824 427048
rect 285784 426494 285812 427042
rect 285772 426488 285824 426494
rect 285772 426430 285824 426436
rect 285784 422294 285812 426430
rect 285784 422266 285904 422294
rect 285680 419484 285732 419490
rect 285680 419426 285732 419432
rect 284484 365016 284536 365022
rect 284484 364958 284536 364964
rect 284484 305040 284536 305046
rect 284484 304982 284536 304988
rect 284392 242208 284444 242214
rect 284392 242150 284444 242156
rect 283104 163532 283156 163538
rect 283104 163474 283156 163480
rect 284300 119400 284352 119406
rect 284300 119342 284352 119348
rect 282920 102808 282972 102814
rect 282920 102750 282972 102756
rect 281540 68944 281592 68950
rect 281540 68886 281592 68892
rect 281540 51740 281592 51746
rect 281540 51682 281592 51688
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 278320 4820 278372 4826
rect 278320 4762 278372 4768
rect 278044 3392 278096 3398
rect 278044 3334 278096 3340
rect 278332 480 278360 4762
rect 279068 490 279096 16546
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 16546
rect 281552 490 281580 51682
rect 283104 3392 283156 3398
rect 283104 3334 283156 3340
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 3334
rect 284312 480 284340 119342
rect 284404 88097 284432 242150
rect 284496 229634 284524 304982
rect 285770 302424 285826 302433
rect 285770 302359 285826 302368
rect 284942 298752 284998 298761
rect 284942 298687 284998 298696
rect 284484 229628 284536 229634
rect 284484 229570 284536 229576
rect 284956 133521 284984 298687
rect 285678 291816 285734 291825
rect 285678 291751 285734 291760
rect 284942 133512 284998 133521
rect 284942 133447 284998 133456
rect 285692 122126 285720 291751
rect 285680 122120 285732 122126
rect 285680 122062 285732 122068
rect 285680 116612 285732 116618
rect 285680 116554 285732 116560
rect 284390 88088 284446 88097
rect 284390 88023 284446 88032
rect 284392 21412 284444 21418
rect 284392 21354 284444 21360
rect 284404 16574 284432 21354
rect 285692 16574 285720 116554
rect 285784 107642 285812 302359
rect 285876 252822 285904 422266
rect 285968 264353 285996 436698
rect 286336 391270 286364 571338
rect 287072 452577 287100 595410
rect 287152 541680 287204 541686
rect 287152 541622 287204 541628
rect 287058 452568 287114 452577
rect 287058 452503 287114 452512
rect 287058 450528 287114 450537
rect 287058 450463 287114 450472
rect 286324 391264 286376 391270
rect 286324 391206 286376 391212
rect 285954 264344 286010 264353
rect 285954 264279 286010 264288
rect 285956 258120 286008 258126
rect 285956 258062 286008 258068
rect 285968 254590 285996 258062
rect 285956 254584 286008 254590
rect 285956 254526 286008 254532
rect 285864 252816 285916 252822
rect 285864 252758 285916 252764
rect 285968 144129 285996 254526
rect 287072 242865 287100 450463
rect 287164 402966 287192 541622
rect 287242 467936 287298 467945
rect 287242 467871 287298 467880
rect 287152 402960 287204 402966
rect 287152 402902 287204 402908
rect 287150 268424 287206 268433
rect 287150 268359 287206 268368
rect 287058 242856 287114 242865
rect 287058 242791 287114 242800
rect 285954 144120 286010 144129
rect 285954 144055 286010 144064
rect 285772 107636 285824 107642
rect 285772 107578 285824 107584
rect 286232 107636 286284 107642
rect 286232 107578 286284 107584
rect 286244 106962 286272 107578
rect 286232 106956 286284 106962
rect 286232 106898 286284 106904
rect 287164 62082 287192 268359
rect 287256 262886 287284 467871
rect 288438 459776 288494 459785
rect 288438 459711 288494 459720
rect 288348 456068 288400 456074
rect 288348 456010 288400 456016
rect 288360 455569 288388 456010
rect 287334 455560 287390 455569
rect 287334 455495 287390 455504
rect 288346 455560 288402 455569
rect 288346 455495 288402 455504
rect 287244 262880 287296 262886
rect 287244 262822 287296 262828
rect 287256 180130 287284 262822
rect 287348 258126 287376 455495
rect 287428 419484 287480 419490
rect 287428 419426 287480 419432
rect 287440 418305 287468 419426
rect 287426 418296 287482 418305
rect 287426 418231 287482 418240
rect 288452 264217 288480 459711
rect 288530 452568 288586 452577
rect 288530 452503 288586 452512
rect 288544 451314 288572 452503
rect 288532 451308 288584 451314
rect 288532 451250 288584 451256
rect 288544 267073 288572 451250
rect 288636 439550 288664 604415
rect 295340 598256 295392 598262
rect 295340 598198 295392 598204
rect 293960 596828 294012 596834
rect 293960 596770 294012 596776
rect 291200 592680 291252 592686
rect 291200 592622 291252 592628
rect 288716 579692 288768 579698
rect 288716 579634 288768 579640
rect 288624 439544 288676 439550
rect 288624 439486 288676 439492
rect 288530 267064 288586 267073
rect 288530 266999 288586 267008
rect 288438 264208 288494 264217
rect 288438 264143 288494 264152
rect 287336 258120 287388 258126
rect 287336 258062 287388 258068
rect 287244 180124 287296 180130
rect 287244 180066 287296 180072
rect 288452 158001 288480 264143
rect 288636 261497 288664 439486
rect 288728 411942 288756 579634
rect 289820 567860 289872 567866
rect 289820 567802 289872 567808
rect 289832 464370 289860 567802
rect 290004 466540 290056 466546
rect 290004 466482 290056 466488
rect 289820 464364 289872 464370
rect 289820 464306 289872 464312
rect 289818 456920 289874 456929
rect 289818 456855 289874 456864
rect 288716 411936 288768 411942
rect 288716 411878 288768 411884
rect 288716 295996 288768 296002
rect 288716 295938 288768 295944
rect 288622 261488 288678 261497
rect 288622 261423 288678 261432
rect 288530 250472 288586 250481
rect 288530 250407 288586 250416
rect 288544 224913 288572 250407
rect 288530 224904 288586 224913
rect 288530 224839 288586 224848
rect 288438 157992 288494 158001
rect 288438 157927 288494 157936
rect 288728 146946 288756 295938
rect 289832 245614 289860 456855
rect 289912 431248 289964 431254
rect 289912 431190 289964 431196
rect 289820 245608 289872 245614
rect 289820 245550 289872 245556
rect 289832 244322 289860 245550
rect 289820 244316 289872 244322
rect 289820 244258 289872 244264
rect 289924 229090 289952 431190
rect 290016 346458 290044 466482
rect 291212 375329 291240 592622
rect 291384 498840 291436 498846
rect 291384 498782 291436 498788
rect 291292 474768 291344 474774
rect 291292 474710 291344 474716
rect 291304 427106 291332 474710
rect 291292 427100 291344 427106
rect 291292 427042 291344 427048
rect 291292 403028 291344 403034
rect 291292 402970 291344 402976
rect 291198 375320 291254 375329
rect 291198 375255 291254 375264
rect 290004 346452 290056 346458
rect 290004 346394 290056 346400
rect 290016 345014 290044 346394
rect 290016 344986 290136 345014
rect 290004 294024 290056 294030
rect 290004 293966 290056 293972
rect 289912 229084 289964 229090
rect 289912 229026 289964 229032
rect 290016 151814 290044 293966
rect 290108 272542 290136 344986
rect 291198 301608 291254 301617
rect 291198 301543 291254 301552
rect 290096 272536 290148 272542
rect 290096 272478 290148 272484
rect 289832 151786 290044 151814
rect 289832 147801 289860 151786
rect 289818 147792 289874 147801
rect 289818 147727 289874 147736
rect 288716 146940 288768 146946
rect 288716 146882 288768 146888
rect 289084 140820 289136 140826
rect 289084 140762 289136 140768
rect 287704 140072 287756 140078
rect 287704 140014 287756 140020
rect 287152 62076 287204 62082
rect 287152 62018 287204 62024
rect 287060 24132 287112 24138
rect 287060 24074 287112 24080
rect 287072 16574 287100 24074
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 284956 490 284984 16546
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 16546
rect 287348 490 287376 16546
rect 287716 3534 287744 140014
rect 288440 71052 288492 71058
rect 288440 70994 288492 71000
rect 288348 62076 288400 62082
rect 288348 62018 288400 62024
rect 288360 61402 288388 62018
rect 288348 61396 288400 61402
rect 288348 61338 288400 61344
rect 288452 16574 288480 70994
rect 288452 16546 289032 16574
rect 287704 3528 287756 3534
rect 287704 3470 287756 3476
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 16546
rect 289096 2990 289124 140762
rect 289832 119406 289860 147727
rect 289820 119400 289872 119406
rect 289820 119342 289872 119348
rect 291212 90370 291240 301543
rect 291304 273222 291332 402970
rect 291396 388482 291424 498782
rect 292580 391264 292632 391270
rect 292580 391206 292632 391212
rect 291384 388476 291436 388482
rect 291384 388418 291436 388424
rect 291384 374740 291436 374746
rect 291384 374682 291436 374688
rect 291396 282198 291424 374682
rect 292592 367033 292620 391206
rect 292578 367024 292634 367033
rect 292578 366959 292634 366968
rect 293972 362914 294000 596770
rect 294050 470656 294106 470665
rect 294050 470591 294106 470600
rect 293960 362908 294012 362914
rect 293960 362850 294012 362856
rect 292672 345092 292724 345098
rect 292672 345034 292724 345040
rect 291384 282192 291436 282198
rect 291384 282134 291436 282140
rect 292580 280220 292632 280226
rect 292580 280162 292632 280168
rect 291292 273216 291344 273222
rect 291292 273158 291344 273164
rect 291304 272513 291332 273158
rect 291290 272504 291346 272513
rect 291290 272439 291346 272448
rect 291292 269136 291344 269142
rect 291292 269078 291344 269084
rect 291304 201482 291332 269078
rect 292592 231810 292620 280162
rect 292684 278089 292712 345034
rect 294064 320249 294092 470591
rect 295352 391338 295380 598198
rect 299492 592686 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 702982 332548 703520
rect 348804 703186 348832 703520
rect 348792 703180 348844 703186
rect 348792 703122 348844 703128
rect 332508 702976 332560 702982
rect 332508 702918 332560 702924
rect 364996 702778 365024 703520
rect 397472 702794 397500 703520
rect 413664 703118 413692 703520
rect 413652 703112 413704 703118
rect 413652 703054 413704 703060
rect 429856 703050 429884 703520
rect 429844 703044 429896 703050
rect 429844 702986 429896 702992
rect 462332 702846 462360 703520
rect 364984 702772 365036 702778
rect 364984 702714 365036 702720
rect 397380 702766 397500 702794
rect 462320 702840 462372 702846
rect 462320 702782 462372 702788
rect 397380 702710 397408 702766
rect 397368 702704 397420 702710
rect 397368 702646 397420 702652
rect 478524 702642 478552 703520
rect 494808 702914 494836 703520
rect 494796 702908 494848 702914
rect 494796 702850 494848 702856
rect 478512 702636 478564 702642
rect 478512 702578 478564 702584
rect 527192 702506 527220 703520
rect 543476 702574 543504 703520
rect 543464 702568 543516 702574
rect 543464 702510 543516 702516
rect 527180 702500 527232 702506
rect 527180 702442 527232 702448
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 582840 700324 582892 700330
rect 582840 700266 582892 700272
rect 582470 697232 582526 697241
rect 582470 697167 582526 697176
rect 582378 617536 582434 617545
rect 582378 617471 582434 617480
rect 582392 607170 582420 617471
rect 582380 607164 582432 607170
rect 582380 607106 582432 607112
rect 299480 592680 299532 592686
rect 299480 592622 299532 592628
rect 296720 591320 296772 591326
rect 296720 591262 296772 591268
rect 295430 536072 295486 536081
rect 295430 536007 295486 536016
rect 295340 391332 295392 391338
rect 295340 391274 295392 391280
rect 295444 371210 295472 536007
rect 295524 434784 295576 434790
rect 295524 434726 295576 434732
rect 295432 371204 295484 371210
rect 295432 371146 295484 371152
rect 294144 337408 294196 337414
rect 294144 337350 294196 337356
rect 294050 320240 294106 320249
rect 294050 320175 294106 320184
rect 294064 316034 294092 320175
rect 293972 316006 294092 316034
rect 292670 278080 292726 278089
rect 292670 278015 292726 278024
rect 292672 248464 292724 248470
rect 292672 248406 292724 248412
rect 292580 231804 292632 231810
rect 292580 231746 292632 231752
rect 292684 204270 292712 248406
rect 292672 204264 292724 204270
rect 292672 204206 292724 204212
rect 291292 201476 291344 201482
rect 291292 201418 291344 201424
rect 293972 199442 294000 316006
rect 294156 259418 294184 337350
rect 295536 315314 295564 434726
rect 296732 363730 296760 591262
rect 582378 591016 582434 591025
rect 582378 590951 582434 590960
rect 582392 584458 582420 590951
rect 582380 584452 582432 584458
rect 582380 584394 582432 584400
rect 302240 578264 302292 578270
rect 302240 578206 302292 578212
rect 298100 495508 298152 495514
rect 298100 495450 298152 495456
rect 296812 437504 296864 437510
rect 296812 437446 296864 437452
rect 296720 363724 296772 363730
rect 296720 363666 296772 363672
rect 295616 340944 295668 340950
rect 295616 340886 295668 340892
rect 295524 315308 295576 315314
rect 295524 315250 295576 315256
rect 295430 310584 295486 310593
rect 295430 310519 295486 310528
rect 295338 309224 295394 309233
rect 295338 309159 295394 309168
rect 294144 259412 294196 259418
rect 294144 259354 294196 259360
rect 294052 244316 294104 244322
rect 294052 244258 294104 244264
rect 293960 199436 294012 199442
rect 293960 199378 294012 199384
rect 294064 155961 294092 244258
rect 294050 155952 294106 155961
rect 294050 155887 294106 155896
rect 294694 155952 294750 155961
rect 294694 155887 294750 155896
rect 294708 155242 294736 155887
rect 294696 155236 294748 155242
rect 294696 155178 294748 155184
rect 295352 132494 295380 309159
rect 295444 189786 295472 310519
rect 295628 284306 295656 340886
rect 296720 313336 296772 313342
rect 296720 313278 296772 313284
rect 295616 284300 295668 284306
rect 295616 284242 295668 284248
rect 295432 189780 295484 189786
rect 295432 189722 295484 189728
rect 295352 132466 295472 132494
rect 295340 111852 295392 111858
rect 295340 111794 295392 111800
rect 295352 111110 295380 111794
rect 295340 111104 295392 111110
rect 295340 111046 295392 111052
rect 295444 111042 295472 132466
rect 295432 111036 295484 111042
rect 295432 110978 295484 110984
rect 295444 110498 295472 110978
rect 295432 110492 295484 110498
rect 295432 110434 295484 110440
rect 295984 110492 296036 110498
rect 295984 110434 296036 110440
rect 291200 90364 291252 90370
rect 291200 90306 291252 90312
rect 291842 82104 291898 82113
rect 291842 82039 291898 82048
rect 291200 28280 291252 28286
rect 291200 28222 291252 28228
rect 291212 16574 291240 28222
rect 291212 16546 291424 16574
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 289084 2984 289136 2990
rect 289084 2926 289136 2932
rect 290200 480 290228 3470
rect 291396 480 291424 16546
rect 291856 3369 291884 82039
rect 295340 77988 295392 77994
rect 295340 77930 295392 77936
rect 295352 16574 295380 77930
rect 295996 49706 296024 110434
rect 296732 56574 296760 313278
rect 296824 253201 296852 437446
rect 298112 420238 298140 495450
rect 299478 465216 299534 465225
rect 299478 465151 299534 465160
rect 298190 458280 298246 458289
rect 298190 458215 298246 458224
rect 298100 420232 298152 420238
rect 298100 420174 298152 420180
rect 298204 304298 298232 458215
rect 298284 450560 298336 450566
rect 298284 450502 298336 450508
rect 298296 331809 298324 450502
rect 298376 420980 298428 420986
rect 298376 420922 298428 420928
rect 298282 331800 298338 331809
rect 298282 331735 298338 331744
rect 298192 304292 298244 304298
rect 298192 304234 298244 304240
rect 296810 253192 296866 253201
rect 296810 253127 296866 253136
rect 298388 246362 298416 420922
rect 299492 298761 299520 465151
rect 299570 462360 299626 462369
rect 299570 462295 299626 462304
rect 299584 305697 299612 462295
rect 299662 307864 299718 307873
rect 299662 307799 299718 307808
rect 299570 305688 299626 305697
rect 299570 305623 299626 305632
rect 299478 298752 299534 298761
rect 299478 298687 299534 298696
rect 298376 246356 298428 246362
rect 298376 246298 298428 246304
rect 298744 135924 298796 135930
rect 298744 135866 298796 135872
rect 296720 56568 296772 56574
rect 296720 56510 296772 56516
rect 298008 56568 298060 56574
rect 298008 56510 298060 56516
rect 298020 55894 298048 56510
rect 298008 55888 298060 55894
rect 298008 55830 298060 55836
rect 295984 49700 296036 49706
rect 295984 49642 296036 49648
rect 296720 49700 296772 49706
rect 296720 49642 296772 49648
rect 296732 16574 296760 49642
rect 298100 42084 298152 42090
rect 298100 42026 298152 42032
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 291936 11756 291988 11762
rect 291936 11698 291988 11704
rect 291948 3534 291976 11698
rect 293684 6180 293736 6186
rect 293684 6122 293736 6128
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 291842 3360 291898 3369
rect 291842 3295 291898 3304
rect 292580 2984 292632 2990
rect 292580 2926 292632 2932
rect 292592 480 292620 2926
rect 293696 480 293724 6122
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 294892 480 294920 3470
rect 295628 490 295656 16546
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 16546
rect 298112 490 298140 42026
rect 298756 3466 298784 135866
rect 299480 128376 299532 128382
rect 299480 128318 299532 128324
rect 299492 3534 299520 128318
rect 299676 110430 299704 307799
rect 302252 205601 302280 578206
rect 582378 577688 582434 577697
rect 582378 577623 582434 577632
rect 582392 538218 582420 577623
rect 582484 566506 582512 697167
rect 582562 683904 582618 683913
rect 582562 683839 582618 683848
rect 582576 571334 582604 683839
rect 582654 644056 582710 644065
rect 582654 643991 582710 644000
rect 582668 603673 582696 643991
rect 582746 630864 582802 630873
rect 582746 630799 582802 630808
rect 582760 607889 582788 630799
rect 582852 609278 582880 700266
rect 582930 670712 582986 670721
rect 582930 670647 582986 670656
rect 582840 609272 582892 609278
rect 582840 609214 582892 609220
rect 582746 607880 582802 607889
rect 582746 607815 582802 607824
rect 582840 604512 582892 604518
rect 582840 604454 582892 604460
rect 582654 603664 582710 603673
rect 582654 603599 582710 603608
rect 582748 601724 582800 601730
rect 582748 601666 582800 601672
rect 582656 593428 582708 593434
rect 582656 593370 582708 593376
rect 582564 571328 582616 571334
rect 582564 571270 582616 571276
rect 582472 566500 582524 566506
rect 582472 566442 582524 566448
rect 582380 538212 582432 538218
rect 582380 538154 582432 538160
rect 582378 537840 582434 537849
rect 582378 537775 582434 537784
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 302332 456816 302384 456822
rect 302332 456758 302384 456764
rect 302344 293962 302372 456758
rect 580184 456074 580212 458079
rect 580172 456068 580224 456074
rect 580172 456010 580224 456016
rect 582392 419490 582420 537775
rect 582668 511329 582696 593370
rect 582760 524521 582788 601666
rect 582852 564369 582880 604454
rect 582838 564360 582894 564369
rect 582838 564295 582894 564304
rect 582944 538286 582972 670647
rect 582932 538280 582984 538286
rect 582932 538222 582984 538228
rect 582746 524512 582802 524521
rect 582746 524447 582802 524456
rect 582654 511320 582710 511329
rect 582654 511255 582710 511264
rect 582470 471472 582526 471481
rect 582470 471407 582526 471416
rect 582380 419484 582432 419490
rect 582380 419426 582432 419432
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 580276 391270 580304 418231
rect 582484 418130 582512 471407
rect 582656 451308 582708 451314
rect 582656 451250 582708 451256
rect 582564 427100 582616 427106
rect 582564 427042 582616 427048
rect 582472 418124 582524 418130
rect 582472 418066 582524 418072
rect 580264 391264 580316 391270
rect 580264 391206 580316 391212
rect 582380 387116 582432 387122
rect 582380 387058 582432 387064
rect 582392 378457 582420 387058
rect 582378 378448 582434 378457
rect 582378 378383 582434 378392
rect 582470 365120 582526 365129
rect 582470 365055 582526 365064
rect 580908 325712 580960 325718
rect 580908 325654 580960 325660
rect 580920 325281 580948 325654
rect 580906 325272 580962 325281
rect 580906 325207 580962 325216
rect 582378 302288 582434 302297
rect 582378 302223 582434 302232
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 304264 298172 304316 298178
rect 304264 298114 304316 298120
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 302332 293956 302384 293962
rect 302332 293898 302384 293904
rect 304276 250481 304304 298114
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580722 258904 580778 258913
rect 580722 258839 580778 258848
rect 580736 256018 580764 258839
rect 580724 256012 580776 256018
rect 580724 255954 580776 255960
rect 304262 250472 304318 250481
rect 304262 250407 304318 250416
rect 580264 235272 580316 235278
rect 580264 235214 580316 235220
rect 580172 232552 580224 232558
rect 580172 232494 580224 232500
rect 580184 232393 580212 232494
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580276 219065 580304 235214
rect 580356 220108 580408 220114
rect 580356 220050 580408 220056
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 580368 205737 580396 220050
rect 580354 205728 580410 205737
rect 580354 205663 580410 205672
rect 302238 205592 302294 205601
rect 302238 205527 302294 205536
rect 579988 195288 580040 195294
rect 579988 195230 580040 195236
rect 580000 192545 580028 195230
rect 579986 192536 580042 192545
rect 579986 192471 580042 192480
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178702 580212 179143
rect 580172 178696 580224 178702
rect 580172 178638 580224 178644
rect 320180 172576 320232 172582
rect 320180 172518 320232 172524
rect 303620 167068 303672 167074
rect 303620 167010 303672 167016
rect 302240 151836 302292 151842
rect 302240 151778 302292 151784
rect 299664 110424 299716 110430
rect 299664 110366 299716 110372
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 298744 3460 298796 3466
rect 298744 3402 298796 3408
rect 299664 3120 299716 3126
rect 299664 3062 299716 3068
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3062
rect 300780 480 300808 3470
rect 301962 3360 302018 3369
rect 301962 3295 302018 3304
rect 301976 480 302004 3295
rect 302252 3126 302280 151778
rect 302332 19984 302384 19990
rect 302332 19926 302384 19932
rect 302344 16574 302372 19926
rect 303632 16574 303660 167010
rect 309784 134564 309836 134570
rect 309784 134506 309836 134512
rect 305644 124908 305696 124914
rect 305644 124850 305696 124856
rect 302344 16546 303200 16574
rect 303632 16546 303936 16574
rect 302240 3120 302292 3126
rect 302240 3062 302292 3068
rect 303172 480 303200 16546
rect 303908 490 303936 16546
rect 305656 5574 305684 124850
rect 307024 110424 307076 110430
rect 307024 110366 307076 110372
rect 306378 40624 306434 40633
rect 306378 40559 306434 40568
rect 305644 5568 305696 5574
rect 305644 5510 305696 5516
rect 305552 3460 305604 3466
rect 305552 3402 305604 3408
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3402
rect 306392 490 306420 40559
rect 307036 2990 307064 110366
rect 309140 39364 309192 39370
rect 309140 39306 309192 39312
rect 309048 5568 309100 5574
rect 309048 5510 309100 5516
rect 307024 2984 307076 2990
rect 307024 2926 307076 2932
rect 307944 2984 307996 2990
rect 307944 2926 307996 2932
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 2926
rect 309060 480 309088 5510
rect 309152 3534 309180 39306
rect 309796 4214 309824 134506
rect 317418 133104 317474 133113
rect 317418 133039 317474 133048
rect 313280 120760 313332 120766
rect 313280 120702 313332 120708
rect 310518 84824 310574 84833
rect 310518 84759 310574 84768
rect 310532 16574 310560 84759
rect 311900 33788 311952 33794
rect 311900 33730 311952 33736
rect 311912 16574 311940 33730
rect 313292 16574 313320 120702
rect 316040 32428 316092 32434
rect 316040 32370 316092 32376
rect 316052 16574 316080 32370
rect 317432 16574 317460 133039
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 309784 4208 309836 4214
rect 309784 4150 309836 4156
rect 309140 3528 309192 3534
rect 309140 3470 309192 3476
rect 310244 3528 310296 3534
rect 310244 3470 310296 3476
rect 310256 480 310284 3470
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 315028 4208 315080 4214
rect 315028 4150 315080 4156
rect 315040 480 315068 4150
rect 316236 480 316264 16546
rect 317328 4208 317380 4214
rect 317328 4150 317380 4156
rect 317340 480 317368 4150
rect 318076 490 318104 16546
rect 320192 3534 320220 172518
rect 338764 159384 338816 159390
rect 338764 159326 338816 159332
rect 327080 146940 327132 146946
rect 327080 146882 327132 146888
rect 323582 142216 323638 142225
rect 323582 142151 323638 142160
rect 321652 102808 321704 102814
rect 321652 102750 321704 102756
rect 320272 66904 320324 66910
rect 320272 66846 320324 66852
rect 320284 16574 320312 66846
rect 320284 16546 320496 16574
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 320180 3528 320232 3534
rect 320180 3470 320232 3476
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3470
rect 320468 490 320496 16546
rect 321560 14476 321612 14482
rect 321560 14418 321612 14424
rect 321572 3482 321600 14418
rect 321664 4214 321692 102750
rect 322940 55888 322992 55894
rect 322940 55830 322992 55836
rect 322204 26920 322256 26926
rect 322204 26862 322256 26868
rect 321652 4208 321704 4214
rect 321652 4150 321704 4156
rect 321572 3454 322152 3482
rect 322216 3466 322244 26862
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 3454
rect 322204 3460 322256 3466
rect 322204 3402 322256 3408
rect 322952 490 322980 55830
rect 323596 4962 323624 142151
rect 324320 111104 324372 111110
rect 324320 111046 324372 111052
rect 323584 4956 323636 4962
rect 323584 4898 323636 4904
rect 324332 3534 324360 111046
rect 324412 54528 324464 54534
rect 324412 54470 324464 54476
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 54470
rect 327092 16574 327120 146882
rect 335452 131776 335504 131782
rect 335452 131718 335504 131724
rect 327724 99408 327776 99414
rect 327724 99350 327776 99356
rect 327092 16546 327672 16574
rect 326804 4956 326856 4962
rect 326804 4898 326856 4904
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326816 480 326844 4898
rect 327644 3210 327672 16546
rect 327736 3330 327764 99350
rect 331220 93152 331272 93158
rect 331220 93094 331272 93100
rect 330392 15904 330444 15910
rect 330392 15846 330444 15852
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 327724 3324 327776 3330
rect 327724 3266 327776 3272
rect 327644 3182 328040 3210
rect 328012 480 328040 3182
rect 329208 480 329236 3402
rect 330404 480 330432 15846
rect 331232 490 331260 93094
rect 334622 91760 334678 91769
rect 334622 91695 334678 91704
rect 333980 64184 334032 64190
rect 333980 64126 334032 64132
rect 333992 6914 334020 64126
rect 334636 16574 334664 91695
rect 335360 50380 335412 50386
rect 335360 50322 335412 50328
rect 334636 16546 334756 16574
rect 333992 6886 334664 6914
rect 333888 4140 333940 4146
rect 333888 4082 333940 4088
rect 332692 3324 332744 3330
rect 332692 3266 332744 3272
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 3266
rect 333900 480 333928 4082
rect 334636 490 334664 6886
rect 334728 3466 334756 16546
rect 335372 3482 335400 50322
rect 335464 4146 335492 131718
rect 338120 76560 338172 76566
rect 338120 76502 338172 76508
rect 338132 16574 338160 76502
rect 338132 16546 338712 16574
rect 337476 4208 337528 4214
rect 337476 4150 337528 4156
rect 335452 4140 335504 4146
rect 335452 4082 335504 4088
rect 334716 3460 334768 3466
rect 335372 3454 336320 3482
rect 334716 3402 334768 3408
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3454
rect 337488 480 337516 4150
rect 338684 480 338712 16546
rect 338776 3330 338804 159326
rect 349804 144968 349856 144974
rect 349804 144910 349856 144916
rect 340880 127628 340932 127634
rect 340880 127570 340932 127576
rect 339500 69080 339552 69086
rect 339500 69022 339552 69028
rect 338764 3324 338816 3330
rect 338764 3266 338816 3272
rect 339512 490 339540 69022
rect 340892 4214 340920 127570
rect 342904 106956 342956 106962
rect 342904 106898 342956 106904
rect 342916 16574 342944 106898
rect 345020 61396 345072 61402
rect 345020 61338 345072 61344
rect 345032 16574 345060 61338
rect 342916 16546 343036 16574
rect 345032 16546 345336 16574
rect 340972 13116 341024 13122
rect 340972 13058 341024 13064
rect 340880 4208 340932 4214
rect 340880 4150 340932 4156
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 13058
rect 342904 10328 342956 10334
rect 342904 10270 342956 10276
rect 342168 3324 342220 3330
rect 342168 3266 342220 3272
rect 342180 480 342208 3266
rect 342916 490 342944 10270
rect 343008 4826 343036 16546
rect 342996 4820 343048 4826
rect 342996 4762 343048 4768
rect 344560 3460 344612 3466
rect 344560 3402 344612 3408
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3402
rect 345308 490 345336 16546
rect 346400 7608 346452 7614
rect 346400 7550 346452 7556
rect 346412 3398 346440 7550
rect 349816 5574 349844 144910
rect 351920 126268 351972 126274
rect 351920 126210 351972 126216
rect 349804 5568 349856 5574
rect 349804 5510 349856 5516
rect 350540 5568 350592 5574
rect 350540 5510 350592 5516
rect 346952 4820 347004 4826
rect 346952 4762 347004 4768
rect 346400 3392 346452 3398
rect 346400 3334 346452 3340
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 4762
rect 350552 3482 350580 5510
rect 350460 3454 350580 3482
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 348056 3324 348108 3330
rect 348056 3266 348108 3272
rect 348068 480 348096 3266
rect 349264 480 349292 3334
rect 350460 480 350488 3454
rect 351932 3330 351960 126210
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99346 580212 99447
rect 580172 99340 580224 99346
rect 580172 99282 580224 99288
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 353300 57248 353352 57254
rect 353300 57190 353352 57196
rect 351920 3324 351972 3330
rect 351920 3266 351972 3272
rect 353312 2922 353340 57190
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 582392 3482 582420 302223
rect 582484 252521 582512 365055
rect 582576 351937 582604 427042
rect 582668 404977 582696 451250
rect 582746 431624 582802 431633
rect 582746 431559 582802 431568
rect 582654 404968 582710 404977
rect 582654 404903 582710 404912
rect 582760 390561 582788 431559
rect 582746 390552 582802 390561
rect 582746 390487 582802 390496
rect 582562 351928 582618 351937
rect 582562 351863 582618 351872
rect 582654 312080 582710 312089
rect 582654 312015 582710 312024
rect 582562 289912 582618 289921
rect 582562 289847 582618 289856
rect 582470 252512 582526 252521
rect 582470 252447 582526 252456
rect 582472 248464 582524 248470
rect 582472 248406 582524 248412
rect 582484 245585 582512 248406
rect 582470 245576 582526 245585
rect 582470 245511 582526 245520
rect 582472 196648 582524 196654
rect 582472 196590 582524 196596
rect 582208 3454 582420 3482
rect 581000 3324 581052 3330
rect 581000 3266 581052 3272
rect 351644 2916 351696 2922
rect 351644 2858 351696 2864
rect 353300 2916 353352 2922
rect 353300 2858 353352 2864
rect 351656 480 351684 2858
rect 581012 480 581040 3266
rect 582208 480 582236 3454
rect 582484 3210 582512 196590
rect 582576 3330 582604 289847
rect 582668 250510 582696 312015
rect 582656 250504 582708 250510
rect 582656 250446 582708 250452
rect 582654 236056 582710 236065
rect 582654 235991 582710 236000
rect 582668 152697 582696 235991
rect 583024 175296 583076 175302
rect 583024 175238 583076 175244
rect 582838 165880 582894 165889
rect 582838 165815 582894 165824
rect 582654 152688 582710 152697
rect 582654 152623 582710 152632
rect 582748 149116 582800 149122
rect 582748 149058 582800 149064
rect 582656 138712 582708 138718
rect 582656 138654 582708 138660
rect 582668 19825 582696 138654
rect 582760 59673 582788 149058
rect 582852 124166 582880 165815
rect 582930 150512 582986 150521
rect 582930 150447 582986 150456
rect 582840 124160 582892 124166
rect 582840 124102 582892 124108
rect 582944 112849 582972 150447
rect 583036 139369 583064 175238
rect 583116 155236 583168 155242
rect 583116 155178 583168 155184
rect 583022 139360 583078 139369
rect 583022 139295 583078 139304
rect 583128 126041 583156 155178
rect 583114 126032 583170 126041
rect 583114 125967 583170 125976
rect 582930 112840 582986 112849
rect 582930 112775 582986 112784
rect 583024 89004 583076 89010
rect 583024 88946 583076 88952
rect 582838 87544 582894 87553
rect 582838 87479 582894 87488
rect 582746 59664 582802 59673
rect 582746 59599 582802 59608
rect 582654 19816 582710 19825
rect 582654 19751 582710 19760
rect 582852 6633 582880 87479
rect 582930 80744 582986 80753
rect 582930 80679 582986 80688
rect 582944 33153 582972 80679
rect 583036 73001 583064 88946
rect 583022 72992 583078 73001
rect 583022 72927 583078 72936
rect 582930 33144 582986 33153
rect 582930 33079 582986 33088
rect 582838 6624 582894 6633
rect 582838 6559 582894 6568
rect 582564 3324 582616 3330
rect 582564 3266 582616 3272
rect 582484 3182 583432 3210
rect 583404 480 583432 3182
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 3330 579944 3386 580000
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3422 501744 3478 501800
rect 3330 475632 3386 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 2778 410488 2834 410544
rect 3422 397432 3478 397488
rect 3422 380840 3478 380896
rect 3514 371320 3570 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 11058 333240 11114 333296
rect 4066 319232 4122 319288
rect 3422 306176 3478 306232
rect 5538 306448 5594 306504
rect 4158 294480 4214 294536
rect 3514 293120 3570 293176
rect 3514 267144 3570 267200
rect 3422 254088 3478 254144
rect 3422 241068 3424 241088
rect 3424 241068 3476 241088
rect 3476 241068 3478 241088
rect 3422 241032 3478 241068
rect 2778 215872 2834 215928
rect 3974 214940 4030 214976
rect 3974 214920 3976 214940
rect 3976 214920 4028 214940
rect 4028 214920 4030 214940
rect 3330 201864 3386 201920
rect 3422 188808 3478 188864
rect 2870 162868 2872 162888
rect 2872 162868 2924 162888
rect 2924 162868 2926 162888
rect 2870 162832 2926 162868
rect 3146 149776 3202 149832
rect 2870 136720 2926 136776
rect 3422 134816 3478 134872
rect 2870 110608 2926 110664
rect 3054 97552 3110 97608
rect 3514 84632 3570 84688
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 3422 58520 3478 58576
rect 3514 45464 3570 45520
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 12438 300056 12494 300112
rect 11150 298696 11206 298752
rect 24858 346976 24914 347032
rect 20718 338680 20774 338736
rect 17958 335416 18014 335472
rect 16578 331744 16634 331800
rect 19338 155216 19394 155272
rect 22742 334056 22798 334112
rect 22098 324400 22154 324456
rect 30378 330384 30434 330440
rect 27618 327664 27674 327720
rect 28998 322088 29054 322144
rect 31758 233824 31814 233880
rect 37278 318824 37334 318880
rect 36542 295976 36598 296032
rect 35898 30912 35954 30968
rect 26514 6160 26570 6216
rect 40038 323584 40094 323640
rect 39946 260072 40002 260128
rect 39854 255856 39910 255912
rect 42798 188264 42854 188320
rect 50986 440816 51042 440872
rect 48134 386960 48190 387016
rect 48134 264968 48190 265024
rect 46846 255856 46902 255912
rect 46938 43424 46994 43480
rect 50894 289040 50950 289096
rect 50802 267960 50858 268016
rect 50710 264968 50766 265024
rect 52274 434696 52330 434752
rect 52274 308352 52330 308408
rect 50894 150456 50950 150512
rect 53470 270680 53526 270736
rect 52274 149640 52330 149696
rect 57702 533296 57758 533352
rect 56506 425040 56562 425096
rect 55034 262792 55090 262848
rect 53562 141344 53618 141400
rect 53470 139440 53526 139496
rect 50986 88168 51042 88224
rect 54942 143520 54998 143576
rect 53746 139440 53802 139496
rect 55034 138080 55090 138136
rect 57794 389136 57850 389192
rect 57794 275168 57850 275224
rect 59174 284552 59230 284608
rect 58990 230424 59046 230480
rect 59266 283192 59322 283248
rect 59174 250008 59230 250064
rect 59082 153176 59138 153232
rect 61842 519424 61898 519480
rect 60462 241304 60518 241360
rect 60738 266464 60794 266520
rect 63130 439456 63186 439512
rect 63130 425040 63186 425096
rect 61934 282104 61990 282160
rect 61750 159296 61806 159352
rect 61750 158752 61806 158808
rect 56414 90888 56470 90944
rect 56598 80688 56654 80744
rect 53838 44784 53894 44840
rect 55218 28192 55274 28248
rect 59266 70216 59322 70272
rect 61934 158752 61990 158808
rect 64694 529080 64750 529136
rect 63406 391448 63462 391504
rect 63314 272040 63370 272096
rect 63222 179424 63278 179480
rect 66902 579944 66958 580000
rect 66166 575864 66222 575920
rect 67454 581032 67510 581088
rect 67362 575048 67418 575104
rect 65982 569880 66038 569936
rect 65890 563352 65946 563408
rect 65982 548256 66038 548312
rect 65890 535336 65946 535392
rect 66810 573144 66866 573200
rect 67546 577224 67602 577280
rect 67454 572600 67510 572656
rect 67454 570152 67510 570208
rect 66902 567432 66958 567488
rect 66442 564848 66498 564904
rect 66810 560632 66866 560688
rect 66810 559272 66866 559328
rect 66810 557912 66866 557968
rect 66534 555192 66590 555248
rect 66902 553560 66958 553616
rect 66166 546760 66222 546816
rect 67362 545400 67418 545456
rect 66810 544040 66866 544096
rect 66258 543360 66314 543416
rect 66258 541320 66314 541376
rect 66258 539960 66314 540016
rect 67362 538736 67418 538792
rect 66166 462848 66222 462904
rect 67454 451832 67510 451888
rect 66074 435240 66130 435296
rect 65982 432520 66038 432576
rect 65890 414024 65946 414080
rect 66810 433336 66866 433392
rect 66166 430344 66222 430400
rect 66074 403688 66130 403744
rect 65982 397296 66038 397352
rect 65982 393388 65984 393408
rect 65984 393388 66036 393408
rect 66036 393388 66038 393408
rect 65982 393352 66038 393388
rect 65982 375944 66038 376000
rect 63314 160656 63370 160712
rect 63222 124344 63278 124400
rect 64510 138216 64566 138272
rect 65890 283192 65946 283248
rect 65890 275984 65946 276040
rect 66626 429276 66682 429312
rect 66626 429256 66628 429276
rect 66628 429256 66680 429276
rect 66680 429256 66682 429276
rect 66810 427352 66866 427408
rect 66626 425176 66682 425232
rect 66810 424088 66866 424144
rect 66258 423272 66314 423328
rect 67178 422184 67234 422240
rect 66902 421096 66958 421152
rect 66626 418920 66682 418976
rect 66994 418124 67050 418160
rect 66994 418104 66996 418124
rect 66996 418104 67048 418124
rect 67048 418104 67050 418124
rect 66810 415928 66866 415984
rect 66810 414840 66866 414896
rect 66626 412936 66682 412992
rect 66902 411848 66958 411904
rect 66810 410760 66866 410816
rect 66810 408856 66866 408912
rect 66902 407768 66958 407824
rect 66810 406680 66866 406736
rect 66810 404504 66866 404560
rect 66810 401512 66866 401568
rect 66810 399608 66866 399664
rect 66534 398520 66590 398576
rect 67086 397468 67088 397488
rect 67088 397468 67140 397488
rect 67140 397468 67142 397488
rect 67086 397432 67142 397468
rect 66810 392264 66866 392320
rect 67362 420008 67418 420064
rect 72974 699760 73030 699816
rect 75918 599256 75974 599312
rect 73526 582528 73582 582584
rect 75366 580896 75422 580952
rect 82726 582664 82782 582720
rect 88982 603200 89038 603256
rect 94870 583344 94926 583400
rect 93766 581168 93822 581224
rect 70950 580760 71006 580816
rect 79966 580760 80022 580816
rect 84658 580760 84714 580816
rect 89258 580760 89314 580816
rect 67730 575864 67786 575920
rect 67638 566616 67694 566672
rect 67638 556552 67694 556608
rect 95238 563624 95294 563680
rect 95146 558832 95148 558852
rect 95148 558832 95200 558852
rect 95200 558832 95202 558852
rect 95146 558796 95202 558832
rect 94686 558592 94742 558648
rect 67822 552200 67878 552256
rect 69662 539008 69718 539064
rect 69662 536152 69718 536208
rect 68926 535472 68982 535528
rect 67730 529216 67786 529272
rect 68926 467880 68982 467936
rect 67546 431432 67602 431488
rect 67454 417016 67510 417072
rect 70858 448604 70860 448624
rect 70860 448604 70912 448624
rect 70912 448604 70914 448624
rect 70858 448568 70914 448604
rect 69662 438776 69718 438832
rect 68374 434696 68430 434752
rect 69294 434288 69350 434344
rect 73066 539552 73122 539608
rect 72422 535472 72478 535528
rect 76746 539552 76802 539608
rect 75734 460944 75790 461000
rect 74538 460128 74594 460184
rect 73158 454688 73214 454744
rect 74446 452920 74502 452976
rect 67730 428168 67786 428224
rect 67638 409672 67694 409728
rect 67270 405592 67326 405648
rect 67362 400424 67418 400480
rect 67270 395292 67272 395312
rect 67272 395292 67324 395312
rect 67324 395292 67326 395312
rect 67270 395256 67326 395292
rect 67822 402600 67878 402656
rect 67454 397432 67510 397488
rect 67270 386280 67326 386336
rect 67546 396344 67602 396400
rect 67730 394440 67786 394496
rect 67454 383560 67510 383616
rect 67822 377984 67878 378040
rect 67638 357312 67694 357368
rect 66258 282920 66314 282976
rect 66810 278840 66866 278896
rect 66166 272584 66222 272640
rect 66718 268232 66774 268288
rect 66258 264988 66314 265024
rect 66258 264968 66260 264988
rect 66260 264968 66312 264988
rect 66312 264968 66314 264988
rect 66258 264152 66314 264208
rect 66258 263336 66314 263392
rect 66350 262792 66406 262848
rect 66258 262520 66314 262576
rect 66258 261704 66314 261760
rect 66350 260888 66406 260944
rect 66626 258440 66682 258496
rect 66258 257624 66314 257680
rect 66718 255176 66774 255232
rect 66166 252728 66222 252784
rect 66626 252728 66682 252784
rect 65982 238584 66038 238640
rect 65982 133592 66038 133648
rect 66626 251912 66682 251968
rect 66258 251132 66260 251152
rect 66260 251132 66312 251152
rect 66312 251132 66314 251152
rect 66258 251096 66314 251132
rect 66626 247832 66682 247888
rect 66534 243752 66590 243808
rect 66902 276392 66958 276448
rect 66902 275576 66958 275632
rect 66902 273944 66958 274000
rect 66902 272312 66958 272368
rect 66902 270680 66958 270736
rect 66902 269864 66958 269920
rect 66902 266600 66958 266656
rect 66994 260072 67050 260128
rect 67270 260072 67326 260128
rect 66902 256012 66958 256048
rect 66902 255992 66904 256012
rect 66904 255992 66956 256012
rect 66956 255992 66958 256012
rect 66902 254360 66958 254416
rect 66902 253544 66958 253600
rect 80058 538328 80114 538384
rect 81990 538736 82046 538792
rect 74814 433608 74870 433664
rect 75458 436056 75514 436112
rect 76194 433608 76250 433664
rect 80058 457408 80114 457464
rect 84014 538056 84070 538112
rect 84290 533296 84346 533352
rect 88338 535472 88394 535528
rect 85762 530576 85818 530632
rect 80334 436464 80390 436520
rect 80058 436192 80114 436248
rect 80978 434016 81034 434072
rect 77482 433744 77538 433800
rect 78218 433744 78274 433800
rect 78126 433608 78182 433664
rect 81898 433608 81954 433664
rect 82910 433608 82966 433664
rect 88982 482840 89038 482896
rect 88982 481616 89038 481672
rect 83738 440816 83794 440872
rect 83830 433608 83886 433664
rect 84566 433608 84622 433664
rect 85854 433744 85910 433800
rect 88430 436328 88486 436384
rect 93398 536696 93454 536752
rect 89350 436736 89406 436792
rect 89902 436192 89958 436248
rect 94594 538872 94650 538928
rect 94778 540232 94834 540288
rect 95882 582528 95938 582584
rect 95422 565800 95478 565856
rect 95330 555464 95386 555520
rect 96894 578856 96950 578912
rect 98642 583344 98698 583400
rect 97906 577496 97962 577552
rect 97906 576680 97962 576736
rect 97906 575048 97962 575104
rect 97538 573416 97594 573472
rect 97262 572600 97318 572656
rect 97722 571396 97778 571432
rect 97722 571376 97724 571396
rect 97724 571376 97776 571396
rect 97776 571376 97778 571396
rect 97906 570016 97962 570072
rect 96710 569064 96766 569120
rect 97906 569064 97962 569120
rect 97906 567196 97908 567216
rect 97908 567196 97960 567216
rect 97960 567196 97962 567216
rect 97906 567160 97962 567196
rect 97906 562536 97962 562592
rect 96802 561040 96858 561096
rect 97906 561040 97962 561096
rect 96710 556824 96766 556880
rect 96618 552064 96674 552120
rect 96894 559544 96950 559600
rect 97906 556844 97962 556880
rect 97906 556824 97908 556844
rect 97908 556824 97960 556844
rect 97960 556824 97962 556844
rect 96986 554104 97042 554160
rect 96894 541728 96950 541784
rect 96710 526360 96766 526416
rect 95330 520920 95386 520976
rect 95238 512624 95294 512680
rect 94594 500112 94650 500168
rect 95698 434288 95754 434344
rect 96710 436056 96766 436112
rect 92754 434152 92810 434208
rect 97906 552744 97962 552800
rect 97814 552064 97870 552120
rect 97078 545672 97134 545728
rect 97538 544312 97594 544368
rect 97538 542952 97594 543008
rect 97906 541728 97962 541784
rect 101402 551928 101458 551984
rect 106922 581168 106978 581224
rect 98366 438096 98422 438152
rect 96986 436056 97042 436112
rect 100206 434288 100262 434344
rect 106278 450472 106334 450528
rect 104898 434560 104954 434616
rect 109038 474000 109094 474056
rect 109682 474000 109738 474056
rect 107658 436056 107714 436112
rect 133694 598168 133750 598224
rect 119342 582664 119398 582720
rect 116122 553968 116178 554024
rect 113822 449792 113878 449848
rect 101218 433744 101274 433800
rect 85946 433608 86002 433664
rect 87234 433608 87290 433664
rect 89994 433608 90050 433664
rect 90730 433608 90786 433664
rect 91558 433608 91614 433664
rect 93030 433608 93086 433664
rect 98458 433608 98514 433664
rect 99838 433608 99894 433664
rect 100666 433608 100722 433664
rect 106738 433608 106794 433664
rect 109498 433608 109554 433664
rect 111706 433608 111762 433664
rect 113270 425992 113326 426048
rect 113178 420824 113234 420880
rect 113086 407108 113142 407144
rect 113086 407088 113088 407108
rect 113088 407088 113140 407108
rect 113140 407088 113142 407108
rect 72422 390904 72478 390960
rect 84382 390904 84438 390960
rect 80150 390768 80206 390824
rect 80978 390768 81034 390824
rect 83186 390768 83242 390824
rect 70398 369008 70454 369064
rect 72422 385056 72478 385112
rect 71686 384920 71742 384976
rect 71686 369008 71742 369064
rect 67914 280472 67970 280528
rect 67546 279656 67602 279712
rect 67546 278024 67602 278080
rect 67454 263336 67510 263392
rect 67362 256808 67418 256864
rect 66902 248648 66958 248704
rect 66902 242936 66958 242992
rect 66902 242120 66958 242176
rect 67822 249464 67878 249520
rect 67362 247016 67418 247072
rect 67454 246200 67510 246256
rect 67638 240080 67694 240136
rect 67454 234504 67510 234560
rect 66902 131960 66958 132016
rect 66810 131144 66866 131200
rect 66810 130600 66866 130656
rect 66718 129784 66774 129840
rect 66810 128968 66866 129024
rect 66810 126792 66866 126848
rect 66074 125976 66130 126032
rect 66810 124344 66866 124400
rect 66994 123800 67050 123856
rect 66902 122984 66958 123040
rect 66350 122168 66406 122224
rect 66810 121372 66866 121408
rect 66810 121352 66812 121372
rect 66812 121352 66864 121372
rect 66864 121352 66866 121372
rect 66902 120536 66958 120592
rect 66810 120028 66812 120048
rect 66812 120028 66864 120048
rect 66864 120028 66866 120048
rect 66810 119992 66866 120028
rect 66902 119176 66958 119232
rect 66626 117544 66682 117600
rect 66626 116184 66682 116240
rect 66810 115368 66866 115424
rect 66902 114552 66958 114608
rect 66810 113736 66866 113792
rect 66902 113192 66958 113248
rect 66810 112376 66866 112432
rect 66810 111560 66866 111616
rect 66902 110744 66958 110800
rect 66902 110200 66958 110256
rect 66074 108568 66130 108624
rect 65890 103128 65946 103184
rect 64694 85448 64750 85504
rect 66810 107752 66866 107808
rect 66810 106936 66866 106992
rect 66626 106392 66682 106448
rect 66626 105596 66682 105632
rect 66626 105576 66628 105596
rect 66628 105576 66680 105596
rect 66680 105576 66682 105596
rect 66810 104796 66812 104816
rect 66812 104796 66864 104816
rect 66864 104796 66866 104816
rect 66810 104760 66866 104796
rect 67270 103944 67326 104000
rect 66442 102584 66498 102640
rect 66718 101768 66774 101824
rect 66810 100952 66866 101008
rect 66810 99628 66812 99648
rect 66812 99628 66864 99648
rect 66864 99628 66866 99648
rect 66810 99592 66866 99628
rect 66810 98776 66866 98832
rect 67546 149116 67602 149152
rect 67546 149096 67548 149116
rect 67548 149096 67600 149116
rect 67600 149096 67602 149116
rect 68466 285912 68522 285968
rect 68558 282140 68560 282160
rect 68560 282140 68612 282160
rect 68612 282140 68614 282160
rect 68558 282104 68614 282140
rect 68190 258712 68246 258768
rect 69202 304136 69258 304192
rect 71042 313928 71098 313984
rect 70306 307672 70362 307728
rect 69662 303592 69718 303648
rect 69202 283736 69258 283792
rect 70076 283736 70132 283792
rect 70214 283464 70270 283520
rect 73066 387640 73122 387696
rect 77206 390360 77262 390416
rect 77206 388728 77262 388784
rect 77390 388456 77446 388512
rect 71962 283736 72018 283792
rect 77206 321408 77262 321464
rect 75918 321000 75974 321056
rect 77206 321000 77262 321056
rect 72836 283736 72892 283792
rect 74630 285504 74686 285560
rect 80242 388456 80298 388512
rect 80150 375944 80206 376000
rect 78586 313928 78642 313984
rect 77298 306584 77354 306640
rect 75458 292576 75514 292632
rect 75274 284416 75330 284472
rect 74630 284280 74686 284336
rect 75458 285504 75514 285560
rect 76562 303592 76618 303648
rect 82174 390496 82230 390552
rect 81438 388456 81494 388512
rect 80886 385600 80942 385656
rect 83554 387232 83610 387288
rect 82726 339516 82782 339552
rect 82726 339496 82728 339516
rect 82728 339496 82780 339516
rect 82780 339496 82782 339516
rect 82726 316648 82782 316704
rect 79966 311072 80022 311128
rect 78218 284416 78274 284472
rect 79322 287000 79378 287056
rect 79322 285912 79378 285968
rect 82634 300192 82690 300248
rect 80886 289856 80942 289912
rect 80426 285776 80482 285832
rect 83094 285912 83150 285968
rect 82634 285776 82690 285832
rect 85026 388320 85082 388376
rect 86866 387096 86922 387152
rect 87142 390904 87198 390960
rect 87878 390904 87934 390960
rect 86958 376488 87014 376544
rect 84106 370504 84162 370560
rect 84014 304136 84070 304192
rect 84106 285912 84162 285968
rect 89626 385736 89682 385792
rect 88430 379344 88486 379400
rect 87602 317328 87658 317384
rect 88246 317328 88302 317384
rect 87602 316104 87658 316160
rect 86866 313928 86922 313984
rect 86774 304272 86830 304328
rect 85854 287136 85910 287192
rect 84658 285504 84714 285560
rect 86774 287136 86830 287192
rect 86866 283600 86922 283656
rect 88246 308488 88302 308544
rect 91282 384240 91338 384296
rect 90362 329840 90418 329896
rect 89718 311208 89774 311264
rect 88982 287680 89038 287736
rect 90270 286048 90326 286104
rect 89810 283464 89866 283520
rect 91006 312432 91062 312488
rect 91006 286048 91062 286104
rect 92018 390360 92074 390416
rect 99654 390904 99710 390960
rect 104254 390904 104310 390960
rect 93766 382880 93822 382936
rect 92478 311888 92534 311944
rect 91374 307672 91430 307728
rect 95146 313928 95202 313984
rect 94502 311072 94558 311128
rect 91282 285504 91338 285560
rect 93950 285640 94006 285696
rect 94042 283464 94098 283520
rect 94686 283464 94742 283520
rect 96986 390360 97042 390416
rect 99286 389136 99342 389192
rect 103794 390768 103850 390824
rect 97538 387776 97594 387832
rect 99286 382064 99342 382120
rect 99286 370640 99342 370696
rect 95330 306992 95386 307048
rect 95238 288496 95294 288552
rect 70950 283192 71006 283248
rect 71962 283192 72018 283248
rect 73250 283192 73306 283248
rect 97906 284824 97962 284880
rect 98090 284416 98146 284472
rect 83462 283056 83518 283112
rect 88614 283056 88670 283112
rect 92386 283056 92442 283112
rect 95330 282920 95386 282976
rect 69018 282684 69020 282704
rect 69020 282684 69072 282704
rect 69072 282684 69074 282704
rect 69018 282648 69074 282684
rect 68926 281152 68982 281208
rect 100758 388592 100814 388648
rect 101954 385736 102010 385792
rect 101402 304136 101458 304192
rect 100022 289856 100078 289912
rect 99102 284552 99158 284608
rect 98090 267824 98146 267880
rect 98918 283328 98974 283384
rect 98918 282784 98974 282840
rect 99102 279520 99158 279576
rect 99470 270408 99526 270464
rect 99010 267996 99012 268016
rect 99012 267996 99064 268016
rect 99064 267996 99066 268016
rect 99010 267960 99066 267996
rect 69018 244296 69074 244352
rect 69846 241712 69902 241768
rect 70950 241712 71006 241768
rect 68834 241440 68890 241496
rect 68834 240080 68890 240136
rect 67914 236544 67970 236600
rect 69386 239944 69442 240000
rect 67822 136040 67878 136096
rect 67730 127608 67786 127664
rect 68558 128152 68614 128208
rect 67822 118360 67878 118416
rect 69662 134680 69718 134736
rect 71318 241440 71374 241496
rect 70398 146376 70454 146432
rect 70214 137944 70270 138000
rect 70306 134836 70362 134872
rect 70306 134816 70308 134836
rect 70308 134816 70360 134836
rect 70360 134816 70362 134836
rect 72606 239808 72662 239864
rect 72882 145016 72938 145072
rect 71410 141344 71466 141400
rect 70490 139576 70546 139632
rect 72330 137400 72386 137456
rect 74630 241168 74686 241224
rect 73802 239944 73858 240000
rect 73250 227568 73306 227624
rect 73158 138352 73214 138408
rect 73066 135088 73122 135144
rect 74814 238856 74870 238912
rect 74814 235864 74870 235920
rect 76562 238584 76618 238640
rect 76010 238312 76066 238368
rect 75182 163376 75238 163432
rect 74722 162016 74778 162072
rect 73802 142296 73858 142352
rect 74262 137264 74318 137320
rect 77942 236000 77998 236056
rect 77574 233144 77630 233200
rect 76654 165688 76710 165744
rect 76010 142432 76066 142488
rect 76654 136584 76710 136640
rect 79322 238720 79378 238776
rect 78034 138624 78090 138680
rect 80610 237224 80666 237280
rect 79414 236680 79470 236736
rect 80610 236000 80666 236056
rect 81806 241304 81862 241360
rect 82726 241576 82782 241632
rect 79966 141480 80022 141536
rect 79322 137400 79378 137456
rect 79046 136856 79102 136912
rect 80610 141344 80666 141400
rect 83278 235320 83334 235376
rect 85578 239944 85634 240000
rect 85578 238720 85634 238776
rect 86682 240080 86738 240136
rect 82818 217912 82874 217968
rect 85486 227704 85542 227760
rect 81438 152360 81494 152416
rect 81898 136720 81954 136776
rect 81070 136176 81126 136232
rect 82082 136856 82138 136912
rect 82818 151816 82874 151872
rect 88430 239400 88486 239456
rect 89626 239400 89682 239456
rect 86314 175752 86370 175808
rect 86314 175344 86370 175400
rect 86222 172488 86278 172544
rect 83462 142568 83518 142624
rect 86314 151816 86370 151872
rect 86314 145016 86370 145072
rect 86866 144744 86922 144800
rect 86866 140120 86922 140176
rect 86314 139984 86370 140040
rect 87050 137536 87106 137592
rect 87050 135904 87106 135960
rect 87602 148280 87658 148336
rect 87694 137264 87750 137320
rect 90362 241712 90418 241768
rect 92386 240760 92442 240816
rect 91006 238584 91062 238640
rect 90362 236544 90418 236600
rect 91098 238448 91154 238504
rect 91098 237360 91154 237416
rect 92294 236680 92350 236736
rect 89718 167048 89774 167104
rect 88522 137944 88578 138000
rect 92386 236544 92442 236600
rect 93490 240080 93546 240136
rect 95698 239944 95754 240000
rect 97078 240080 97134 240136
rect 95882 239944 95938 240000
rect 93674 176724 93730 176760
rect 93674 176704 93676 176724
rect 93676 176704 93728 176724
rect 93728 176704 93730 176724
rect 92754 157392 92810 157448
rect 93766 138216 93822 138272
rect 93950 145560 94006 145616
rect 94686 138080 94742 138136
rect 95146 136720 95202 136776
rect 94686 131824 94742 131880
rect 67454 100136 67510 100192
rect 66810 94968 66866 95024
rect 67178 93336 67234 93392
rect 67362 97960 67418 98016
rect 67362 97144 67418 97200
rect 67546 97144 67602 97200
rect 67546 95784 67602 95840
rect 66166 78512 66222 78568
rect 68558 92656 68614 92712
rect 94778 98504 94834 98560
rect 69018 92520 69074 92576
rect 68558 86672 68614 86728
rect 66258 55800 66314 55856
rect 69018 82048 69074 82104
rect 69708 92520 69764 92576
rect 71180 92656 71236 92712
rect 70398 73752 70454 73808
rect 72836 92656 72892 92712
rect 71778 88168 71834 88224
rect 73342 92384 73398 92440
rect 73710 92248 73766 92304
rect 74814 92112 74870 92168
rect 74354 90888 74410 90944
rect 72606 88168 72662 88224
rect 72606 86808 72662 86864
rect 76378 86536 76434 86592
rect 74538 72392 74594 72448
rect 78034 88032 78090 88088
rect 79322 79328 79378 79384
rect 81530 89392 81586 89448
rect 82634 91160 82690 91216
rect 83002 89664 83058 89720
rect 82082 88168 82138 88224
rect 83462 91160 83518 91216
rect 84658 89528 84714 89584
rect 84842 89528 84898 89584
rect 84106 87896 84162 87952
rect 87234 89528 87290 89584
rect 91006 92384 91062 92440
rect 90362 83408 90418 83464
rect 89902 82728 89958 82784
rect 85670 26832 85726 26888
rect 91834 92384 91890 92440
rect 92754 92248 92810 92304
rect 92386 91976 92442 92032
rect 91282 85312 91338 85368
rect 92478 71032 92534 71088
rect 93858 68176 93914 68232
rect 94778 89800 94834 89856
rect 95422 127608 95478 127664
rect 95330 120264 95386 120320
rect 95238 89392 95294 89448
rect 95146 77152 95202 77208
rect 95974 139440 96030 139496
rect 96618 130872 96674 130928
rect 95974 126384 96030 126440
rect 96066 120300 96068 120320
rect 96068 120300 96120 120320
rect 96120 120300 96122 120320
rect 96066 120264 96122 120300
rect 95974 86536 96030 86592
rect 97170 123256 97226 123312
rect 97078 120808 97134 120864
rect 99286 261432 99342 261488
rect 98090 260888 98146 260944
rect 98642 258440 98698 258496
rect 98182 242528 98238 242584
rect 97538 144744 97594 144800
rect 97906 133864 97962 133920
rect 97906 132232 97962 132288
rect 97538 131416 97594 131472
rect 97722 130872 97778 130928
rect 97538 130056 97594 130112
rect 97906 128424 97962 128480
rect 97630 127064 97686 127120
rect 97906 126248 97962 126304
rect 97814 125432 97870 125488
rect 97906 124616 97962 124672
rect 97906 124108 97908 124128
rect 97908 124108 97960 124128
rect 97960 124108 97962 124128
rect 97906 124072 97962 124108
rect 97354 122440 97410 122496
rect 97906 121624 97962 121680
rect 97906 119448 97962 119504
rect 97906 118652 97962 118688
rect 97906 118632 97908 118652
rect 97908 118632 97960 118652
rect 97960 118632 97962 118652
rect 97906 117000 97962 117056
rect 97354 116456 97410 116512
rect 97906 115640 97962 115696
rect 97814 114824 97870 114880
rect 97262 114008 97318 114064
rect 96710 111868 96712 111888
rect 96712 111868 96764 111888
rect 96764 111868 96766 111888
rect 96710 111832 96766 111868
rect 96802 111016 96858 111072
rect 96710 96600 96766 96656
rect 96618 83408 96674 83464
rect 97538 113464 97594 113520
rect 97906 112648 97962 112704
rect 97354 111832 97410 111888
rect 97814 110200 97870 110256
rect 97906 109656 97962 109712
rect 97906 108024 97962 108080
rect 97906 107208 97962 107264
rect 97906 106664 97962 106720
rect 97906 104236 97962 104272
rect 97906 104216 97908 104236
rect 97908 104216 97960 104236
rect 97960 104216 97962 104236
rect 99378 249192 99434 249248
rect 98642 103536 98698 103592
rect 97906 103436 97908 103456
rect 97908 103436 97960 103456
rect 97960 103436 97962 103456
rect 97906 103400 97962 103436
rect 97906 102856 97962 102912
rect 97906 102076 97908 102096
rect 97908 102076 97960 102096
rect 97960 102076 97962 102096
rect 97906 102040 97962 102076
rect 97906 101224 97962 101280
rect 97538 100408 97594 100464
rect 97906 99592 97962 99648
rect 97906 98232 97962 98288
rect 97906 95260 97962 95296
rect 97906 95240 97908 95260
rect 97908 95240 97960 95260
rect 97960 95240 97962 95260
rect 97538 94424 97594 94480
rect 97906 93608 97962 93664
rect 97354 92792 97410 92848
rect 94502 67496 94558 67552
rect 98182 15816 98238 15872
rect 98826 214512 98882 214568
rect 100206 283056 100262 283112
rect 100758 281832 100814 281888
rect 100850 280200 100906 280256
rect 100758 279384 100814 279440
rect 101494 282648 101550 282704
rect 101402 278568 101458 278624
rect 100758 276120 100814 276176
rect 100758 275304 100814 275360
rect 100942 274488 100998 274544
rect 100850 273672 100906 273728
rect 100758 272856 100814 272912
rect 101954 276936 102010 276992
rect 101494 272448 101550 272504
rect 100850 272040 100906 272096
rect 101218 271224 101274 271280
rect 104162 385600 104218 385656
rect 103426 382880 103482 382936
rect 102138 287136 102194 287192
rect 100758 270408 100814 270464
rect 100758 268776 100814 268832
rect 100758 267144 100814 267200
rect 100758 266328 100814 266384
rect 100942 264696 100998 264752
rect 100758 263880 100814 263936
rect 100666 262248 100722 262304
rect 100574 258032 100630 258088
rect 100850 260616 100906 260672
rect 100758 259800 100814 259856
rect 100942 260072 100998 260128
rect 100758 258984 100814 259040
rect 101678 258168 101734 258224
rect 102046 257372 102102 257408
rect 102046 257352 102048 257372
rect 102048 257352 102100 257372
rect 102100 257352 102102 257372
rect 100758 256536 100814 256592
rect 100850 255720 100906 255776
rect 100758 254088 100814 254144
rect 100758 250824 100814 250880
rect 100942 252456 100998 252512
rect 100942 251096 100998 251152
rect 101494 250008 101550 250064
rect 100850 248376 100906 248432
rect 101034 245928 101090 245984
rect 100850 245148 100852 245168
rect 100852 245148 100904 245168
rect 100904 245148 100906 245168
rect 100850 245112 100906 245148
rect 100942 244296 100998 244352
rect 100850 243500 100906 243536
rect 100850 243480 100852 243500
rect 100852 243480 100904 243500
rect 100904 243480 100906 243500
rect 100850 242664 100906 242720
rect 100758 237360 100814 237416
rect 100758 124788 100760 124808
rect 100760 124788 100812 124808
rect 100812 124788 100814 124808
rect 100758 124752 100814 124788
rect 100022 102176 100078 102232
rect 98918 99048 98974 99104
rect 98826 87896 98882 87952
rect 101586 246744 101642 246800
rect 101586 148280 101642 148336
rect 101402 85176 101458 85232
rect 98918 84088 98974 84144
rect 102874 241440 102930 241496
rect 102138 152360 102194 152416
rect 102874 151816 102930 151872
rect 102782 147872 102838 147928
rect 101678 93064 101734 93120
rect 102230 124752 102286 124808
rect 102782 117816 102838 117872
rect 102322 93200 102378 93256
rect 105266 390904 105322 390960
rect 105910 390904 105966 390960
rect 105726 389000 105782 389056
rect 111982 390904 112038 390960
rect 112902 391040 112958 391096
rect 112902 390768 112958 390824
rect 106094 389000 106150 389056
rect 104806 370504 104862 370560
rect 105542 302368 105598 302424
rect 104438 285776 104494 285832
rect 104254 253272 104310 253328
rect 104162 233144 104218 233200
rect 106094 382200 106150 382256
rect 106094 378664 106150 378720
rect 106002 278704 106058 278760
rect 106186 320592 106242 320648
rect 106094 266328 106150 266384
rect 105634 241848 105690 241904
rect 105542 239944 105598 240000
rect 104254 223488 104310 223544
rect 106738 389272 106794 389328
rect 108302 389816 108358 389872
rect 107658 372544 107714 372600
rect 106370 276936 106426 276992
rect 102322 86672 102378 86728
rect 104990 204312 105046 204368
rect 105542 162832 105598 162888
rect 105542 132504 105598 132560
rect 105542 128968 105598 129024
rect 104990 111832 105046 111888
rect 107566 287680 107622 287736
rect 108394 380704 108450 380760
rect 108394 379480 108450 379536
rect 108946 379480 109002 379536
rect 108302 269320 108358 269376
rect 108394 254360 108450 254416
rect 108302 238040 108358 238096
rect 107014 90344 107070 90400
rect 107014 88032 107070 88088
rect 106278 71732 106334 71768
rect 106278 71712 106280 71732
rect 106280 71712 106332 71732
rect 106332 71712 106334 71732
rect 108394 236000 108450 236056
rect 108394 233144 108450 233200
rect 109038 361528 109094 361584
rect 109038 360168 109094 360224
rect 109682 360168 109738 360224
rect 109038 236000 109094 236056
rect 112626 280744 112682 280800
rect 112442 266328 112498 266384
rect 110602 238312 110658 238368
rect 110418 235184 110474 235240
rect 108394 90480 108450 90536
rect 110510 232600 110566 232656
rect 111062 232464 111118 232520
rect 113822 424904 113878 424960
rect 113362 418920 113418 418976
rect 113270 385736 113326 385792
rect 114650 420008 114706 420064
rect 114558 417832 114614 417888
rect 114466 406408 114522 406464
rect 113454 402328 113510 402384
rect 115202 516704 115258 516760
rect 115202 463528 115258 463584
rect 114834 430072 114890 430128
rect 114742 413888 114798 413944
rect 115754 433336 115810 433392
rect 115846 432248 115902 432304
rect 115570 431160 115626 431216
rect 115754 429256 115810 429312
rect 115846 428168 115902 428224
rect 115846 425992 115902 426048
rect 115846 424088 115902 424144
rect 115846 423000 115902 423056
rect 115202 421912 115258 421968
rect 115846 418920 115902 418976
rect 115846 416780 115848 416800
rect 115848 416780 115900 416800
rect 115900 416780 115902 416800
rect 115846 416744 115902 416780
rect 115846 415656 115902 415712
rect 115846 414840 115902 414896
rect 115754 412664 115810 412720
rect 115018 411576 115074 411632
rect 115570 410488 115626 410544
rect 115846 409672 115902 409728
rect 115846 408584 115902 408640
rect 115202 406408 115258 406464
rect 115110 396344 115166 396400
rect 114834 382880 114890 382936
rect 115846 405628 115848 405648
rect 115848 405628 115900 405648
rect 115900 405628 115902 405648
rect 115846 405592 115902 405628
rect 115846 404504 115902 404560
rect 115846 403416 115902 403472
rect 115754 401240 115810 401296
rect 115570 400424 115626 400480
rect 115846 399336 115902 399392
rect 115846 398284 115848 398304
rect 115848 398284 115900 398304
rect 115900 398284 115902 398304
rect 115846 398248 115902 398284
rect 115570 397160 115626 397216
rect 115846 395256 115902 395312
rect 115846 394168 115902 394224
rect 115846 393080 115902 393136
rect 115846 392012 115902 392048
rect 115846 391992 115848 392012
rect 115848 391992 115900 392012
rect 115900 391992 115902 392012
rect 118606 456864 118662 456920
rect 116582 449792 116638 449848
rect 118606 436736 118662 436792
rect 119342 452784 119398 452840
rect 119342 438096 119398 438152
rect 118790 436736 118846 436792
rect 116122 385600 116178 385656
rect 115938 301416 115994 301472
rect 114466 271088 114522 271144
rect 113914 247560 113970 247616
rect 113822 244840 113878 244896
rect 112626 239400 112682 239456
rect 113914 237224 113970 237280
rect 115202 235320 115258 235376
rect 113178 92248 113234 92304
rect 115386 231104 115442 231160
rect 115294 138624 115350 138680
rect 115202 88168 115258 88224
rect 118698 389816 118754 389872
rect 117962 387096 118018 387152
rect 117318 378664 117374 378720
rect 116030 232600 116086 232656
rect 120078 380840 120134 380896
rect 117962 235320 118018 235376
rect 116766 234504 116822 234560
rect 117318 206216 117374 206272
rect 122102 376624 122158 376680
rect 119342 228248 119398 228304
rect 120078 185544 120134 185600
rect 120722 83952 120778 84008
rect 123574 409128 123630 409184
rect 123574 389136 123630 389192
rect 123482 378664 123538 378720
rect 123666 379344 123722 379400
rect 122102 251096 122158 251152
rect 122194 235864 122250 235920
rect 122930 89528 122986 89584
rect 124218 237904 124274 237960
rect 123574 192480 123630 192536
rect 124954 309712 125010 309768
rect 129002 383560 129058 383616
rect 129002 337320 129058 337376
rect 126242 335960 126298 336016
rect 125046 291760 125102 291816
rect 124954 153176 125010 153232
rect 124954 124072 125010 124128
rect 126426 296112 126482 296168
rect 130382 324944 130438 325000
rect 129186 317464 129242 317520
rect 129002 128968 129058 129024
rect 127622 119312 127678 119368
rect 127622 117952 127678 118008
rect 126978 95784 127034 95840
rect 126334 79328 126390 79384
rect 127622 68176 127678 68232
rect 130474 322904 130530 322960
rect 130474 276664 130530 276720
rect 133786 530576 133842 530632
rect 133142 327800 133198 327856
rect 133142 264968 133198 265024
rect 133142 236544 133198 236600
rect 135902 538192 135958 538248
rect 134706 334600 134762 334656
rect 135902 331880 135958 331936
rect 134706 153176 134762 153232
rect 137834 392536 137890 392592
rect 137466 366988 137522 367024
rect 137466 366968 137468 366988
rect 137468 366968 137520 366988
rect 137520 366968 137522 366988
rect 137742 366968 137798 367024
rect 137282 365608 137338 365664
rect 137282 328616 137338 328672
rect 137466 278704 137522 278760
rect 137926 333376 137982 333432
rect 140594 489912 140650 489968
rect 139398 386280 139454 386336
rect 142618 593272 142674 593328
rect 141974 384920 142030 384976
rect 141974 384376 142030 384432
rect 140594 321408 140650 321464
rect 140042 313248 140098 313304
rect 138662 307808 138718 307864
rect 138662 294480 138718 294536
rect 137834 233824 137890 233880
rect 138662 227568 138718 227624
rect 141422 304136 141478 304192
rect 140134 262792 140190 262848
rect 140226 261432 140282 261488
rect 140134 160112 140190 160168
rect 143446 593272 143502 593328
rect 143262 433200 143318 433256
rect 142250 375264 142306 375320
rect 142802 375264 142858 375320
rect 143630 537376 143686 537432
rect 143354 429256 143410 429312
rect 142802 347656 142858 347712
rect 143262 347656 143318 347712
rect 142802 346976 142858 347032
rect 142894 326304 142950 326360
rect 142802 301688 142858 301744
rect 141606 262520 141662 262576
rect 145562 527720 145618 527776
rect 144642 413888 144698 413944
rect 144182 326440 144238 326496
rect 144274 314744 144330 314800
rect 143446 282784 143502 282840
rect 143446 282104 143502 282160
rect 142986 280472 143042 280528
rect 142986 169768 143042 169824
rect 146206 463664 146262 463720
rect 145562 392536 145618 392592
rect 144826 376488 144882 376544
rect 144642 238584 144698 238640
rect 144642 238040 144698 238096
rect 144182 117952 144238 118008
rect 145654 305632 145710 305688
rect 145562 296112 145618 296168
rect 145562 295296 145618 295352
rect 145562 271224 145618 271280
rect 147586 454008 147642 454064
rect 145654 156032 145710 156088
rect 147218 313928 147274 313984
rect 147034 310664 147090 310720
rect 147126 265512 147182 265568
rect 148966 400152 149022 400208
rect 148506 338816 148562 338872
rect 150346 515344 150402 515400
rect 150254 369688 150310 369744
rect 151082 476176 151138 476232
rect 151634 476176 151690 476232
rect 150438 333376 150494 333432
rect 150438 332560 150494 332616
rect 149794 328480 149850 328536
rect 149702 318008 149758 318064
rect 149702 306584 149758 306640
rect 149794 271088 149850 271144
rect 151266 465704 151322 465760
rect 151174 456048 151230 456104
rect 150530 299376 150586 299432
rect 150530 298696 150586 298752
rect 152462 533296 152518 533352
rect 151726 409128 151782 409184
rect 151082 267008 151138 267064
rect 151174 264152 151230 264208
rect 151174 258712 151230 258768
rect 151266 136176 151322 136232
rect 152922 460128 152978 460184
rect 152922 377984 152978 378040
rect 152922 377304 152978 377360
rect 153934 466520 153990 466576
rect 153934 436736 153990 436792
rect 154394 417424 154450 417480
rect 152646 285640 152702 285696
rect 155222 466520 155278 466576
rect 155682 439456 155738 439512
rect 155590 419600 155646 419656
rect 155682 390904 155738 390960
rect 154394 389816 154450 389872
rect 154486 378800 154542 378856
rect 155774 380160 155830 380216
rect 155222 357312 155278 357368
rect 153842 347656 153898 347712
rect 153198 338000 153254 338056
rect 154026 334736 154082 334792
rect 153842 310392 153898 310448
rect 154026 320728 154082 320784
rect 153934 278024 153990 278080
rect 153842 208256 153898 208312
rect 153842 185544 153898 185600
rect 152646 137808 152702 137864
rect 154026 276664 154082 276720
rect 154026 268368 154082 268424
rect 155222 261432 155278 261488
rect 153934 164328 153990 164384
rect 153934 144880 153990 144936
rect 155958 394712 156014 394768
rect 157154 481752 157210 481808
rect 156602 390904 156658 390960
rect 155406 260072 155462 260128
rect 155314 233144 155370 233200
rect 155406 226888 155462 226944
rect 155406 153720 155462 153776
rect 158626 498752 158682 498808
rect 158534 461488 158590 461544
rect 158442 390632 158498 390688
rect 157982 368328 158038 368384
rect 156602 251912 156658 251968
rect 156050 242120 156106 242176
rect 155958 137944 156014 138000
rect 156418 137944 156474 138000
rect 156418 137264 156474 137320
rect 158718 471144 158774 471200
rect 158626 338680 158682 338736
rect 158534 303456 158590 303512
rect 160834 581032 160890 581088
rect 159362 471144 159418 471200
rect 160742 382880 160798 382936
rect 160006 301552 160062 301608
rect 157982 274760 158038 274816
rect 157338 160656 157394 160712
rect 157338 160248 157394 160304
rect 158074 160248 158130 160304
rect 159362 246200 159418 246256
rect 158626 92112 158682 92168
rect 160282 282920 160338 282976
rect 160098 281424 160154 281480
rect 160098 280744 160154 280800
rect 159546 145016 159602 145072
rect 162582 401648 162638 401704
rect 162122 384240 162178 384296
rect 161294 383696 161350 383752
rect 162122 377304 162178 377360
rect 163502 483656 163558 483712
rect 162122 327120 162178 327176
rect 162122 284824 162178 284880
rect 160190 136040 160246 136096
rect 163502 401648 163558 401704
rect 164054 326984 164110 327040
rect 163686 303456 163742 303512
rect 164974 567840 165030 567896
rect 164330 371864 164386 371920
rect 164146 305632 164202 305688
rect 162766 93200 162822 93256
rect 164146 251912 164202 251968
rect 164146 220768 164202 220824
rect 164146 133048 164202 133104
rect 164146 94424 164202 94480
rect 163594 71032 163650 71088
rect 164330 261432 164386 261488
rect 165526 469240 165582 469296
rect 166354 451152 166410 451208
rect 166354 450472 166410 450528
rect 165526 320728 165582 320784
rect 166262 301688 166318 301744
rect 165526 261432 165582 261488
rect 166906 344256 166962 344312
rect 166814 287680 166870 287736
rect 166814 280064 166870 280120
rect 166814 279384 166870 279440
rect 166814 249056 166870 249112
rect 166262 230424 166318 230480
rect 166814 230424 166870 230480
rect 166814 162016 166870 162072
rect 167642 386008 167698 386064
rect 168194 423680 168250 423736
rect 168102 331744 168158 331800
rect 167090 280064 167146 280120
rect 171046 601976 171102 602032
rect 169574 475496 169630 475552
rect 169022 333240 169078 333296
rect 168470 297336 168526 297392
rect 168378 282104 168434 282160
rect 168194 260752 168250 260808
rect 168470 250416 168526 250472
rect 168470 230288 168526 230344
rect 170494 541048 170550 541104
rect 170402 382064 170458 382120
rect 169666 341400 169722 341456
rect 169206 269048 169262 269104
rect 169758 264832 169814 264888
rect 169206 251096 169262 251152
rect 169574 251132 169576 251152
rect 169576 251132 169628 251152
rect 169628 251132 169630 251152
rect 169574 251096 169630 251132
rect 169666 230288 169722 230344
rect 169666 224848 169722 224904
rect 169298 150592 169354 150648
rect 169114 145560 169170 145616
rect 169206 137264 169262 137320
rect 169298 124752 169354 124808
rect 173162 553968 173218 554024
rect 173254 523640 173310 523696
rect 173622 489096 173678 489152
rect 173162 469240 173218 469296
rect 172518 453872 172574 453928
rect 172518 438096 172574 438152
rect 171046 383424 171102 383480
rect 171046 346976 171102 347032
rect 170310 264832 170366 264888
rect 170770 254224 170826 254280
rect 171046 246200 171102 246256
rect 171782 258848 171838 258904
rect 175186 608640 175242 608696
rect 173530 388864 173586 388920
rect 173530 387640 173586 387696
rect 173254 379344 173310 379400
rect 173254 346432 173310 346488
rect 172058 242120 172114 242176
rect 171874 233144 171930 233200
rect 173806 387640 173862 387696
rect 172518 239400 172574 239456
rect 171966 116456 172022 116512
rect 171874 102176 171930 102232
rect 172426 102176 172482 102232
rect 172426 95784 172482 95840
rect 174634 366288 174690 366344
rect 174542 321544 174598 321600
rect 173346 233008 173402 233064
rect 173254 148008 173310 148064
rect 173254 141480 173310 141536
rect 173806 95240 173862 95296
rect 173162 73752 173218 73808
rect 175094 322224 175150 322280
rect 175186 321544 175242 321600
rect 176106 453736 176162 453792
rect 176014 444216 176070 444272
rect 176014 323620 176016 323640
rect 176016 323620 176068 323640
rect 176068 323620 176070 323640
rect 176014 323584 176070 323620
rect 175922 315288 175978 315344
rect 175278 289720 175334 289776
rect 175278 289040 175334 289096
rect 178774 599528 178830 599584
rect 177394 468424 177450 468480
rect 177578 468424 177634 468480
rect 176658 452512 176714 452568
rect 177302 452512 177358 452568
rect 176658 451832 176714 451888
rect 177302 427080 177358 427136
rect 176658 366968 176714 367024
rect 176106 289720 176162 289776
rect 174726 234096 174782 234152
rect 175186 234504 175242 234560
rect 175186 234096 175242 234152
rect 176106 267008 176162 267064
rect 175186 92384 175242 92440
rect 177578 419600 177634 419656
rect 177394 366968 177450 367024
rect 177578 340856 177634 340912
rect 177578 338816 177634 338872
rect 176750 306448 176806 306504
rect 177302 257352 177358 257408
rect 177394 228928 177450 228984
rect 177394 227704 177450 227760
rect 177394 155352 177450 155408
rect 177486 145696 177542 145752
rect 178038 435240 178094 435296
rect 178038 387504 178094 387560
rect 178038 386960 178094 387016
rect 178038 341400 178094 341456
rect 178038 337864 178094 337920
rect 178038 337320 178094 337376
rect 178130 337184 178186 337240
rect 178590 334600 178646 334656
rect 178774 387504 178830 387560
rect 180706 604560 180762 604616
rect 180430 474136 180486 474192
rect 180430 403552 180486 403608
rect 180614 400152 180670 400208
rect 180614 393352 180670 393408
rect 181534 533976 181590 534032
rect 180154 390904 180210 390960
rect 180062 387504 180118 387560
rect 180706 393080 180762 393136
rect 180614 387504 180670 387560
rect 180706 383696 180762 383752
rect 180706 383560 180762 383616
rect 180154 380704 180210 380760
rect 181534 384920 181590 384976
rect 181902 454688 181958 454744
rect 181902 400152 181958 400208
rect 181994 393896 182050 393952
rect 186962 600616 187018 600672
rect 186226 595448 186282 595504
rect 182914 536016 182970 536072
rect 183466 485016 183522 485072
rect 183374 446528 183430 446584
rect 182822 390768 182878 390824
rect 181994 389136 182050 389192
rect 181810 381928 181866 381984
rect 181994 375128 182050 375184
rect 180706 374040 180762 374096
rect 180706 373904 180762 373960
rect 179326 343032 179382 343088
rect 178774 322088 178830 322144
rect 178682 319368 178738 319424
rect 177946 227704 178002 227760
rect 179326 302232 179382 302288
rect 179326 302096 179382 302152
rect 179326 287680 179382 287736
rect 178958 271224 179014 271280
rect 180706 364384 180762 364440
rect 180706 364248 180762 364304
rect 180706 354864 180762 354920
rect 180614 354592 180670 354648
rect 180614 346976 180670 347032
rect 180614 341400 180670 341456
rect 180062 300056 180118 300112
rect 180062 295976 180118 296032
rect 180062 253952 180118 254008
rect 179418 247560 179474 247616
rect 178866 236680 178922 236736
rect 178866 156168 178922 156224
rect 178038 81368 178094 81424
rect 179326 81368 179382 81424
rect 180614 253952 180670 254008
rect 180246 231240 180302 231296
rect 180890 234096 180946 234152
rect 180338 224168 180394 224224
rect 180246 199280 180302 199336
rect 180062 80688 180118 80744
rect 181994 247696 182050 247752
rect 182822 373904 182878 373960
rect 182086 234096 182142 234152
rect 181994 162152 182050 162208
rect 181534 146512 181590 146568
rect 184202 459856 184258 459912
rect 183466 312432 183522 312488
rect 184754 452376 184810 452432
rect 184202 309168 184258 309224
rect 184662 305224 184718 305280
rect 184938 403552 184994 403608
rect 184846 366968 184902 367024
rect 184846 366288 184902 366344
rect 183282 242800 183338 242856
rect 184202 242664 184258 242720
rect 184202 241576 184258 241632
rect 182178 144744 182234 144800
rect 182178 135904 182234 135960
rect 182822 133048 182878 133104
rect 183466 144744 183522 144800
rect 183466 143656 183522 143712
rect 181442 82048 181498 82104
rect 184754 264172 184810 264208
rect 184754 264152 184756 264172
rect 184756 264152 184808 264172
rect 184808 264152 184810 264172
rect 188250 596808 188306 596864
rect 188250 596264 188306 596320
rect 191654 607824 191710 607880
rect 189722 605920 189778 605976
rect 188434 604424 188490 604480
rect 191010 597896 191066 597952
rect 188434 539280 188490 539336
rect 187606 530712 187662 530768
rect 186226 452512 186282 452568
rect 186318 451424 186374 451480
rect 186042 382064 186098 382120
rect 187514 469784 187570 469840
rect 187146 452376 187202 452432
rect 187146 451424 187202 451480
rect 186778 393896 186834 393952
rect 186962 384240 187018 384296
rect 186410 380296 186466 380352
rect 186962 376488 187018 376544
rect 186410 375264 186466 375320
rect 185582 306448 185638 306504
rect 186226 315288 186282 315344
rect 184938 242664 184994 242720
rect 184386 235184 184442 235240
rect 184478 151000 184534 151056
rect 184294 150456 184350 150512
rect 184754 126248 184810 126304
rect 184754 125704 184810 125760
rect 185766 267008 185822 267064
rect 186226 235864 186282 235920
rect 185582 206216 185638 206272
rect 185766 162016 185822 162072
rect 185766 144064 185822 144120
rect 185582 143520 185638 143576
rect 184846 92112 184902 92168
rect 185674 92248 185730 92304
rect 187698 468016 187754 468072
rect 187606 465704 187662 465760
rect 187790 467880 187846 467936
rect 187790 461624 187846 461680
rect 187698 459584 187754 459640
rect 187698 456048 187754 456104
rect 189722 567432 189778 567488
rect 189814 553424 189870 553480
rect 189078 536152 189134 536208
rect 189078 530576 189134 530632
rect 188434 460128 188490 460184
rect 188434 452648 188490 452704
rect 188434 438776 188490 438832
rect 187698 389136 187754 389192
rect 188434 409128 188490 409184
rect 188526 389816 188582 389872
rect 188434 386144 188490 386200
rect 188526 383560 188582 383616
rect 188802 384376 188858 384432
rect 187698 378664 187754 378720
rect 187698 377984 187754 378040
rect 187698 370504 187754 370560
rect 187054 257216 187110 257272
rect 187054 244568 187110 244624
rect 186962 222128 187018 222184
rect 186962 217912 187018 217968
rect 186318 216688 186374 216744
rect 186962 216688 187018 216744
rect 188894 345616 188950 345672
rect 188802 333240 188858 333296
rect 188342 313928 188398 313984
rect 187698 310528 187754 310584
rect 187698 309712 187754 309768
rect 188342 307944 188398 308000
rect 188342 306312 188398 306368
rect 188342 305088 188398 305144
rect 187698 301144 187754 301200
rect 189814 471824 189870 471880
rect 191102 594904 191158 594960
rect 190550 588104 190606 588160
rect 190458 586508 190460 586528
rect 190460 586508 190512 586528
rect 190512 586508 190514 586528
rect 190458 586472 190514 586508
rect 191010 585112 191066 585168
rect 190918 578992 190974 579048
rect 190826 574504 190882 574560
rect 190826 572192 190882 572248
rect 196714 604424 196770 604480
rect 191746 603608 191802 603664
rect 191654 597216 191710 597272
rect 191378 596284 191434 596320
rect 191378 596264 191380 596284
rect 191380 596264 191432 596284
rect 191432 596264 191434 596284
rect 191286 593952 191342 594008
rect 191194 593272 191250 593328
rect 191378 592068 191434 592104
rect 191378 592048 191380 592068
rect 191380 592048 191432 592068
rect 191432 592048 191434 592068
rect 191286 591232 191342 591288
rect 191378 589348 191434 589384
rect 191378 589328 191380 589348
rect 191380 589328 191432 589348
rect 191432 589328 191434 589348
rect 194138 601840 194194 601896
rect 194138 600888 194194 600944
rect 192574 600752 192630 600808
rect 192666 599392 192722 599448
rect 198554 599392 198610 599448
rect 201130 601976 201186 602032
rect 199842 600616 199898 600672
rect 204810 601840 204866 601896
rect 204258 600752 204314 600808
rect 202418 600616 202474 600672
rect 193126 599052 193182 599108
rect 204442 599120 204498 599176
rect 207662 610000 207718 610056
rect 205638 599528 205694 599584
rect 206834 599528 206890 599584
rect 208398 608776 208454 608832
rect 209410 607280 209466 607336
rect 209962 600752 210018 600808
rect 212446 599392 212502 599448
rect 213274 599120 213330 599176
rect 215298 600344 215354 600400
rect 216402 600344 216458 600400
rect 218242 600344 218298 600400
rect 222106 605920 222162 605976
rect 219346 600344 219402 600400
rect 222934 600480 222990 600536
rect 227718 619656 227774 619712
rect 226430 608640 226486 608696
rect 226338 603064 226394 603120
rect 225786 600344 225842 600400
rect 226338 599392 226394 599448
rect 230110 603200 230166 603256
rect 230110 601840 230166 601896
rect 231766 600480 231822 600536
rect 193034 593408 193090 593464
rect 191746 586064 191802 586120
rect 191746 583888 191802 583944
rect 191286 582664 191342 582720
rect 191194 581712 191250 581768
rect 191746 581168 191802 581224
rect 191562 579672 191618 579728
rect 191562 578856 191618 578912
rect 191654 578312 191710 578368
rect 191746 578040 191802 578096
rect 191654 576136 191710 576192
rect 191746 575592 191802 575648
rect 191746 572756 191802 572792
rect 191746 572736 191748 572756
rect 191748 572736 191800 572756
rect 191800 572736 191802 572756
rect 191746 570832 191802 570888
rect 191746 570016 191802 570072
rect 191102 567840 191158 567896
rect 191378 567196 191380 567216
rect 191380 567196 191432 567216
rect 191432 567196 191434 567216
rect 191378 567160 191434 567196
rect 191286 565120 191342 565176
rect 191746 564984 191802 565040
rect 191746 563660 191748 563680
rect 191748 563660 191800 563680
rect 191800 563660 191802 563680
rect 191746 563624 191802 563660
rect 190918 562128 190974 562184
rect 190826 560904 190882 560960
rect 191746 559136 191802 559192
rect 191746 557776 191802 557832
rect 191746 556416 191802 556472
rect 191470 554920 191526 554976
rect 191102 552608 191158 552664
rect 191746 550704 191802 550760
rect 191654 549752 191710 549808
rect 190642 548256 190698 548312
rect 191746 549364 191802 549400
rect 191746 549344 191748 549364
rect 191748 549344 191800 549364
rect 191800 549344 191802 549364
rect 191562 547032 191618 547088
rect 191654 546524 191656 546544
rect 191656 546524 191708 546544
rect 191708 546524 191710 546544
rect 191654 546488 191710 546524
rect 191654 545264 191710 545320
rect 191010 544176 191066 544232
rect 191562 544040 191618 544096
rect 191654 540540 191656 540560
rect 191656 540540 191708 540560
rect 191708 540540 191710 540560
rect 191654 540504 191710 540540
rect 191654 456184 191710 456240
rect 191562 456048 191618 456104
rect 190458 449112 190514 449168
rect 191562 447752 191618 447808
rect 191562 446392 191618 446448
rect 191562 445052 191618 445088
rect 191562 445032 191564 445052
rect 191564 445032 191616 445052
rect 191616 445032 191618 445052
rect 191378 442040 191434 442096
rect 190642 440680 190698 440736
rect 190642 437960 190698 438016
rect 191654 439320 191710 439376
rect 191562 436736 191618 436792
rect 191654 436600 191710 436656
rect 191562 435240 191618 435296
rect 191470 433880 191526 433936
rect 191654 432248 191710 432304
rect 194598 598984 194654 599040
rect 197174 598984 197230 599040
rect 201590 598984 201646 599040
rect 203062 598984 203118 599040
rect 207110 598984 207166 599040
rect 210790 598984 210846 599040
rect 219714 598984 219770 599040
rect 220910 598984 220966 599040
rect 231214 599120 231270 599176
rect 234066 604560 234122 604616
rect 236366 599392 236422 599448
rect 236826 599120 236882 599176
rect 239218 601704 239274 601760
rect 240046 599120 240102 599176
rect 244186 600616 244242 600672
rect 243910 599120 243966 599176
rect 246210 600480 246266 600536
rect 246762 600480 246818 600536
rect 248326 599528 248382 599584
rect 249338 599256 249394 599312
rect 250074 600344 250130 600400
rect 223854 598984 223910 599040
rect 224222 598984 224278 599040
rect 230018 598984 230074 599040
rect 230662 598984 230718 599040
rect 233238 598984 233294 599040
rect 234710 598984 234766 599040
rect 236826 598984 236882 599040
rect 240690 598984 240746 599040
rect 242622 598984 242678 599040
rect 247774 598984 247830 599040
rect 250258 598984 250314 599040
rect 252834 598984 252890 599040
rect 193494 598440 193550 598496
rect 253938 592252 253994 592308
rect 253386 556144 253442 556200
rect 193586 536152 193642 536208
rect 194138 536016 194194 536072
rect 191930 448432 191986 448488
rect 191838 443536 191894 443592
rect 191746 430888 191802 430944
rect 191010 429528 191066 429584
rect 190826 428168 190882 428224
rect 190826 426808 190882 426864
rect 191746 425448 191802 425504
rect 191746 423816 191802 423872
rect 191010 422456 191066 422512
rect 191746 421096 191802 421152
rect 192574 475496 192630 475552
rect 193034 443672 193090 443728
rect 192482 419736 192538 419792
rect 191746 418376 191802 418432
rect 191746 417016 191802 417072
rect 190642 415384 190698 415440
rect 191470 414024 191526 414080
rect 191746 412684 191802 412720
rect 191746 412664 191748 412684
rect 191748 412664 191800 412684
rect 191800 412664 191802 412684
rect 197266 535472 197322 535528
rect 194598 515344 194654 515400
rect 195058 458904 195114 458960
rect 198002 530576 198058 530632
rect 197358 512624 197414 512680
rect 195334 511400 195390 511456
rect 198002 502968 198058 503024
rect 195334 461488 195390 461544
rect 199842 533976 199898 534032
rect 196714 482160 196770 482216
rect 196622 459040 196678 459096
rect 197358 465704 197414 465760
rect 196714 456320 196770 456376
rect 195610 452648 195666 452704
rect 197910 454008 197966 454064
rect 202970 538056 203026 538112
rect 203338 530576 203394 530632
rect 203522 522280 203578 522336
rect 204902 532072 204958 532128
rect 202234 480800 202290 480856
rect 204166 464480 204222 464536
rect 201590 462168 201646 462224
rect 202234 462168 202290 462224
rect 202326 461488 202382 461544
rect 201590 460944 201646 461000
rect 201406 459040 201462 459096
rect 200854 452920 200910 452976
rect 201406 452920 201462 452976
rect 199382 450336 199438 450392
rect 195242 449928 195298 449984
rect 203154 452648 203210 452704
rect 204074 451288 204130 451344
rect 204994 522416 205050 522472
rect 205086 464344 205142 464400
rect 204994 458768 205050 458824
rect 204902 454688 204958 454744
rect 206282 535472 206338 535528
rect 207386 538192 207442 538248
rect 208122 535472 208178 535528
rect 207662 485016 207718 485072
rect 206282 468424 206338 468480
rect 208398 461624 208454 461680
rect 210514 481616 210570 481672
rect 211802 531936 211858 531992
rect 211802 471280 211858 471336
rect 212630 532072 212686 532128
rect 213090 533432 213146 533488
rect 214654 509768 214710 509824
rect 212630 467880 212686 467936
rect 213274 467880 213330 467936
rect 214654 486512 214710 486568
rect 215482 464344 215538 464400
rect 217414 535472 217470 535528
rect 219530 535472 219586 535528
rect 218794 530712 218850 530768
rect 217322 476720 217378 476776
rect 220082 527720 220138 527776
rect 218794 475360 218850 475416
rect 216678 469784 216734 469840
rect 218702 465840 218758 465896
rect 216770 463664 216826 463720
rect 215942 459720 215998 459776
rect 218058 459856 218114 459912
rect 218702 459856 218758 459912
rect 222106 537376 222162 537432
rect 222934 535472 222990 535528
rect 224682 535336 224738 535392
rect 223670 534112 223726 534168
rect 224682 534112 224738 534168
rect 222934 497392 222990 497448
rect 222842 461488 222898 461544
rect 222106 454144 222162 454200
rect 226522 535472 226578 535528
rect 224958 523640 225014 523696
rect 224958 463664 225014 463720
rect 223670 456864 223726 456920
rect 223670 454008 223726 454064
rect 229742 530576 229798 530632
rect 227718 509768 227774 509824
rect 226246 463664 226302 463720
rect 227718 468016 227774 468072
rect 231122 526360 231178 526416
rect 230478 475360 230534 475416
rect 232502 511264 232558 511320
rect 231858 478080 231914 478136
rect 232502 465568 232558 465624
rect 228730 451560 228786 451616
rect 232134 458768 232190 458824
rect 231214 456864 231270 456920
rect 233238 465568 233294 465624
rect 233238 465160 233294 465216
rect 233146 458768 233202 458824
rect 232594 455504 232650 455560
rect 233238 452784 233294 452840
rect 238206 533296 238262 533352
rect 235906 483792 235962 483848
rect 239402 518880 239458 518936
rect 237378 471824 237434 471880
rect 238022 471824 238078 471880
rect 237378 470600 237434 470656
rect 235998 463528 236054 463584
rect 234618 462168 234674 462224
rect 235906 462168 235962 462224
rect 235906 460944 235962 461000
rect 233882 450608 233938 450664
rect 237470 458224 237526 458280
rect 239494 476176 239550 476232
rect 239402 471144 239458 471200
rect 238114 458224 238170 458280
rect 240782 481480 240838 481536
rect 239494 462848 239550 462904
rect 240782 457408 240838 457464
rect 238850 452784 238906 452840
rect 244922 535472 244978 535528
rect 245106 537376 245162 537432
rect 243174 528536 243230 528592
rect 241702 498752 241758 498808
rect 244278 505688 244334 505744
rect 241610 463528 241666 463584
rect 242162 463528 242218 463584
rect 241610 462304 241666 462360
rect 238850 451152 238906 451208
rect 246762 536696 246818 536752
rect 246302 535472 246358 535528
rect 244370 496576 244426 496632
rect 244922 452784 244978 452840
rect 244278 450472 244334 450528
rect 245750 449928 245806 449984
rect 249890 526360 249946 526416
rect 248602 474000 248658 474056
rect 249062 474000 249118 474056
rect 249614 449928 249670 449984
rect 251086 452512 251142 452568
rect 250626 451424 250682 451480
rect 251454 539008 251510 539064
rect 252466 529080 252522 529136
rect 251546 452920 251602 452976
rect 252558 484372 252560 484392
rect 252560 484372 252612 484392
rect 252612 484372 252614 484392
rect 252558 484336 252614 484372
rect 252466 481616 252522 481672
rect 252466 480800 252522 480856
rect 253386 541048 253442 541104
rect 254030 586880 254086 586936
rect 254582 599528 254638 599584
rect 254766 600616 254822 600672
rect 255962 598848 256018 598904
rect 255410 593816 255466 593872
rect 255410 593000 255466 593056
rect 254766 592592 254822 592648
rect 256606 597624 256662 597680
rect 256606 595176 256662 595232
rect 255410 589872 255466 589928
rect 255962 589872 256018 589928
rect 255502 589328 255558 589384
rect 255962 587968 256018 588024
rect 255502 587152 255558 587208
rect 255318 585112 255374 585168
rect 254122 582256 254178 582312
rect 255502 584296 255558 584352
rect 255410 584160 255466 584216
rect 255410 582528 255466 582584
rect 255502 580216 255558 580272
rect 255410 579808 255466 579864
rect 255318 578584 255374 578640
rect 254122 554920 254178 554976
rect 254214 545128 254270 545184
rect 253294 476176 253350 476232
rect 252098 455368 252154 455424
rect 247038 449656 247094 449712
rect 254214 462848 254270 462904
rect 253938 448704 253994 448760
rect 254030 448568 254086 448624
rect 253570 429800 253626 429856
rect 192850 411324 192906 411360
rect 192850 411304 192852 411324
rect 192852 411304 192904 411324
rect 192904 411304 192906 411324
rect 193126 411304 193182 411360
rect 189722 396072 189778 396128
rect 189722 380840 189778 380896
rect 189170 380160 189226 380216
rect 189170 346432 189226 346488
rect 189078 330384 189134 330440
rect 190274 311072 190330 311128
rect 189814 301008 189870 301064
rect 190182 295432 190238 295488
rect 188434 272448 188490 272504
rect 188342 251776 188398 251832
rect 187698 244840 187754 244896
rect 188342 244432 188398 244488
rect 187698 241032 187754 241088
rect 189722 285640 189778 285696
rect 189722 281424 189778 281480
rect 188526 240896 188582 240952
rect 188434 239808 188490 239864
rect 190458 409944 190514 410000
rect 191746 408584 191802 408640
rect 191746 406952 191802 407008
rect 191654 405592 191710 405648
rect 191746 404232 191802 404288
rect 193126 402872 193182 402928
rect 191562 401512 191618 401568
rect 191746 400152 191802 400208
rect 191746 398520 191802 398576
rect 191010 394440 191066 394496
rect 191746 391720 191802 391776
rect 191930 393080 191986 393136
rect 191838 387640 191894 387696
rect 191838 387368 191894 387424
rect 190458 375400 190514 375456
rect 192482 391040 192538 391096
rect 192022 390632 192078 390688
rect 192022 387640 192078 387696
rect 190550 372680 190606 372736
rect 191102 342896 191158 342952
rect 190550 335960 190606 336016
rect 190458 326304 190514 326360
rect 193034 329024 193090 329080
rect 191102 323584 191158 323640
rect 190918 299784 190974 299840
rect 191102 299784 191158 299840
rect 191746 298696 191802 298752
rect 191746 297608 191802 297664
rect 192022 295976 192078 296032
rect 192022 295296 192078 295352
rect 191746 294344 191802 294400
rect 191562 293256 191618 293312
rect 193310 397976 193366 398032
rect 254214 447480 254270 447536
rect 254214 427896 254270 427952
rect 254122 405320 254178 405376
rect 254030 396888 254086 396944
rect 254030 395528 254086 395584
rect 193402 391040 193458 391096
rect 212446 390904 212502 390960
rect 249706 390904 249762 390960
rect 195242 387640 195298 387696
rect 195242 351872 195298 351928
rect 193310 315288 193366 315344
rect 193402 314880 193458 314936
rect 193034 292168 193090 292224
rect 190366 291352 190422 291408
rect 193034 291352 193090 291408
rect 189998 274624 190054 274680
rect 190274 274624 190330 274680
rect 189814 238040 189870 238096
rect 191654 291080 191710 291136
rect 191194 290028 191196 290048
rect 191196 290028 191248 290048
rect 191248 290028 191250 290048
rect 191194 289992 191250 290028
rect 191746 288904 191802 288960
rect 191746 286728 191802 286784
rect 191746 284552 191802 284608
rect 191746 283464 191802 283520
rect 191746 282376 191802 282432
rect 191746 281288 191802 281344
rect 192022 280200 192078 280256
rect 191746 279112 191802 279168
rect 191562 278024 191618 278080
rect 191746 276936 191802 276992
rect 191746 275848 191802 275904
rect 191746 274624 191802 274680
rect 191746 273672 191802 273728
rect 191286 272584 191342 272640
rect 191746 271496 191802 271552
rect 191194 270444 191196 270464
rect 191196 270444 191248 270464
rect 191248 270444 191250 270464
rect 191194 270408 191250 270444
rect 194414 305632 194470 305688
rect 195242 349696 195298 349752
rect 197358 387640 197414 387696
rect 198186 387640 198242 387696
rect 197358 387368 197414 387424
rect 201130 386008 201186 386064
rect 199106 384376 199162 384432
rect 204350 389816 204406 389872
rect 203522 386008 203578 386064
rect 199382 366288 199438 366344
rect 196622 340040 196678 340096
rect 196714 319368 196770 319424
rect 196622 310664 196678 310720
rect 195058 309032 195114 309088
rect 195058 307808 195114 307864
rect 194598 303728 194654 303784
rect 195610 303728 195666 303784
rect 197450 331200 197506 331256
rect 197450 326984 197506 327040
rect 198002 312432 198058 312488
rect 199198 306312 199254 306368
rect 199014 300872 199070 300928
rect 202142 363568 202198 363624
rect 200762 359352 200818 359408
rect 201682 349832 201738 349888
rect 201498 338680 201554 338736
rect 200118 334056 200174 334112
rect 200762 334056 200818 334112
rect 199382 306312 199438 306368
rect 201590 331744 201646 331800
rect 202142 343032 202198 343088
rect 204810 389136 204866 389192
rect 204810 386280 204866 386336
rect 206466 378800 206522 378856
rect 204902 346976 204958 347032
rect 202878 334736 202934 334792
rect 201682 303592 201738 303648
rect 202786 303592 202842 303648
rect 204166 334600 204222 334656
rect 203062 322224 203118 322280
rect 204350 317600 204406 317656
rect 205638 338000 205694 338056
rect 205638 336776 205694 336832
rect 204902 314064 204958 314120
rect 205822 305088 205878 305144
rect 209594 385600 209650 385656
rect 208398 375128 208454 375184
rect 209042 362208 209098 362264
rect 206558 352552 206614 352608
rect 207662 340176 207718 340232
rect 207202 338816 207258 338872
rect 206558 338000 206614 338056
rect 207110 331880 207166 331936
rect 206282 305088 206338 305144
rect 208398 313248 208454 313304
rect 213458 387504 213514 387560
rect 209778 349696 209834 349752
rect 209318 313928 209374 313984
rect 209318 313248 209374 313304
rect 209134 311072 209190 311128
rect 209042 306584 209098 306640
rect 211342 328616 211398 328672
rect 210238 309304 210294 309360
rect 210422 309304 210478 309360
rect 211066 303592 211122 303648
rect 211434 326304 211490 326360
rect 214654 369008 214710 369064
rect 211894 348336 211950 348392
rect 211894 328616 211950 328672
rect 212446 309712 212502 309768
rect 212446 302504 212502 302560
rect 213918 324944 213974 325000
rect 216678 383424 216734 383480
rect 215390 381928 215446 381984
rect 215390 380976 215446 381032
rect 215942 380976 215998 381032
rect 216678 360032 216734 360088
rect 217414 360032 217470 360088
rect 215482 335960 215538 336016
rect 214838 304136 214894 304192
rect 217414 335960 217470 336016
rect 216862 301552 216918 301608
rect 220082 384240 220138 384296
rect 220174 382064 220230 382120
rect 220910 380296 220966 380352
rect 220266 373360 220322 373416
rect 220174 349832 220230 349888
rect 224866 384784 224922 384840
rect 221462 370504 221518 370560
rect 220266 345616 220322 345672
rect 219438 338136 219494 338192
rect 218702 311752 218758 311808
rect 218058 306992 218114 307048
rect 218702 305632 218758 305688
rect 218150 301144 218206 301200
rect 220818 336640 220874 336696
rect 220818 335416 220874 335472
rect 220174 307944 220230 308000
rect 220910 327664 220966 327720
rect 221554 348472 221610 348528
rect 221554 336640 221610 336696
rect 222290 330384 222346 330440
rect 221002 324400 221058 324456
rect 224222 360848 224278 360904
rect 224314 351056 224370 351112
rect 224222 338680 224278 338736
rect 223578 338000 223634 338056
rect 223578 337320 223634 337376
rect 223486 312432 223542 312488
rect 222842 311072 222898 311128
rect 223394 306720 223450 306776
rect 224314 338000 224370 338056
rect 223670 320048 223726 320104
rect 224222 320048 224278 320104
rect 223670 318824 223726 318880
rect 223486 302232 223542 302288
rect 229742 375944 229798 376000
rect 227626 371864 227682 371920
rect 226246 346432 226302 346488
rect 225142 327800 225198 327856
rect 226338 334600 226394 334656
rect 226982 320728 227038 320784
rect 229282 328480 229338 328536
rect 229742 328480 229798 328536
rect 230570 389272 230626 389328
rect 231122 381520 231178 381576
rect 232594 382880 232650 382936
rect 232502 374584 232558 374640
rect 232502 351872 232558 351928
rect 231122 341400 231178 341456
rect 230662 332560 230718 332616
rect 231858 331200 231914 331256
rect 231122 309168 231178 309224
rect 232226 303592 232282 303648
rect 234342 377304 234398 377360
rect 233882 357992 233938 358048
rect 232594 346976 232650 347032
rect 236642 388592 236698 388648
rect 237194 388592 237250 388648
rect 238022 386960 238078 387016
rect 235262 373224 235318 373280
rect 233882 329840 233938 329896
rect 236642 356632 236698 356688
rect 239402 375264 239458 375320
rect 238114 370640 238170 370696
rect 238022 342896 238078 342952
rect 234710 314744 234766 314800
rect 234526 301688 234582 301744
rect 235262 327664 235318 327720
rect 235262 314744 235318 314800
rect 237470 318008 237526 318064
rect 240782 381656 240838 381712
rect 237470 310528 237526 310584
rect 240046 339768 240102 339824
rect 240138 307672 240194 307728
rect 244738 389000 244794 389056
rect 245566 388320 245622 388376
rect 244922 386144 244978 386200
rect 243082 382200 243138 382256
rect 243082 380976 243138 381032
rect 244186 380976 244242 381032
rect 241242 307672 241298 307728
rect 241242 306448 241298 306504
rect 240046 303864 240102 303920
rect 238850 302232 238906 302288
rect 239402 302096 239458 302152
rect 241794 304952 241850 305008
rect 241426 302368 241482 302424
rect 243082 301552 243138 301608
rect 244370 310392 244426 310448
rect 244370 309168 244426 309224
rect 236734 301416 236790 301472
rect 244922 334600 244978 334656
rect 245014 310392 245070 310448
rect 245566 306448 245622 306504
rect 244462 305768 244518 305824
rect 244462 304952 244518 305008
rect 246210 306992 246266 307048
rect 246394 306992 246450 307048
rect 248602 389000 248658 389056
rect 249522 389000 249578 389056
rect 247222 388456 247278 388512
rect 247130 378664 247186 378720
rect 247038 372544 247094 372600
rect 249062 374584 249118 374640
rect 247222 366288 247278 366344
rect 248326 330384 248382 330440
rect 247682 307808 247738 307864
rect 246946 304272 247002 304328
rect 247222 304136 247278 304192
rect 246302 302096 246358 302152
rect 248694 311752 248750 311808
rect 248602 310936 248658 310992
rect 217874 300872 217930 300928
rect 250442 389408 250498 389464
rect 249706 373904 249762 373960
rect 249614 361564 249616 361584
rect 249616 361564 249668 361584
rect 249668 361564 249670 361584
rect 249614 361528 249670 361564
rect 249062 329160 249118 329216
rect 249614 311752 249670 311808
rect 250442 368328 250498 368384
rect 249890 331200 249946 331256
rect 253938 391992 253994 392048
rect 252466 384920 252522 384976
rect 254030 389408 254086 389464
rect 254490 447500 254546 447536
rect 254490 447480 254492 447500
rect 254492 447480 254544 447500
rect 254544 447480 254546 447500
rect 255410 577632 255466 577688
rect 255410 576952 255466 577008
rect 255410 575864 255466 575920
rect 255410 574640 255466 574696
rect 255594 574096 255650 574152
rect 255502 571920 255558 571976
rect 255410 571512 255466 571568
rect 255410 570560 255466 570616
rect 255502 569200 255558 569256
rect 255410 568656 255466 568712
rect 255686 572872 255742 572928
rect 255594 566208 255650 566264
rect 255502 565956 255558 565992
rect 255502 565936 255504 565956
rect 255504 565936 255556 565956
rect 255556 565936 255558 565956
rect 255502 564712 255558 564768
rect 255686 561720 255742 561776
rect 255502 560768 255558 560824
rect 255594 559544 255650 559600
rect 255502 559136 255558 559192
rect 255594 557912 255650 557968
rect 255594 556824 255650 556880
rect 255686 554104 255742 554160
rect 255594 553560 255650 553616
rect 255594 552744 255650 552800
rect 255594 550840 255650 550896
rect 255594 549908 255650 549944
rect 255594 549888 255596 549908
rect 255596 549888 255648 549908
rect 255648 549888 255650 549908
rect 255594 548392 255650 548448
rect 255870 547848 255926 547904
rect 255502 546760 255558 546816
rect 255502 545808 255558 545864
rect 255594 542816 255650 542872
rect 255502 542428 255558 542464
rect 255502 542408 255504 542428
rect 255504 542408 255556 542428
rect 255556 542408 255558 542428
rect 255502 540096 255558 540152
rect 255502 539416 255558 539472
rect 256606 543768 256662 543824
rect 255594 457408 255650 457464
rect 255594 448840 255650 448896
rect 255502 446120 255558 446176
rect 255594 444760 255650 444816
rect 255502 443400 255558 443456
rect 255686 442040 255742 442096
rect 255502 439048 255558 439104
rect 255502 437688 255558 437744
rect 255502 437552 255558 437608
rect 255502 436328 255558 436384
rect 255502 434968 255558 435024
rect 255502 433608 255558 433664
rect 255962 431976 256018 432032
rect 255410 430616 255466 430672
rect 255410 426536 255466 426592
rect 255502 425176 255558 425232
rect 255502 423544 255558 423600
rect 255502 422184 255558 422240
rect 255502 420824 255558 420880
rect 255410 419484 255466 419520
rect 255410 419464 255412 419484
rect 255412 419464 255464 419484
rect 255464 419464 255466 419484
rect 255410 418104 255466 418160
rect 255410 416780 255412 416800
rect 255412 416780 255464 416800
rect 255464 416780 255466 416800
rect 255410 416744 255466 416780
rect 255318 415112 255374 415168
rect 255410 413788 255412 413808
rect 255412 413788 255464 413808
rect 255464 413788 255466 413808
rect 255410 413752 255466 413788
rect 255410 412428 255412 412448
rect 255412 412428 255464 412448
rect 255464 412428 255466 412448
rect 255410 412392 255466 412428
rect 255502 411032 255558 411088
rect 255410 409672 255466 409728
rect 255410 408312 255466 408368
rect 255502 406952 255558 407008
rect 255318 402600 255374 402656
rect 255410 401240 255466 401296
rect 255410 399880 255466 399936
rect 255410 398520 255466 398576
rect 255502 394168 255558 394224
rect 254306 392808 254362 392864
rect 254214 389272 254270 389328
rect 253938 365608 253994 365664
rect 256882 567432 256938 567488
rect 256790 530576 256846 530632
rect 256698 363568 256754 363624
rect 250994 320184 251050 320240
rect 249706 310936 249762 310992
rect 249706 310528 249762 310584
rect 250166 302368 250222 302424
rect 252466 321544 252522 321600
rect 252006 302368 252062 302424
rect 251822 301688 251878 301744
rect 251730 301144 251786 301200
rect 252558 304272 252614 304328
rect 252558 303728 252614 303784
rect 250994 301008 251050 301064
rect 251638 300872 251694 300928
rect 253386 325760 253442 325816
rect 253386 321408 253442 321464
rect 253202 311208 253258 311264
rect 253386 311072 253442 311128
rect 193678 299376 193734 299432
rect 252834 298016 252890 298072
rect 193402 269320 193458 269376
rect 191194 268232 191250 268288
rect 190642 256264 190698 256320
rect 190642 254088 190698 254144
rect 189998 237904 190054 237960
rect 188342 155216 188398 155272
rect 187698 153720 187754 153776
rect 187698 145832 187754 145888
rect 189078 149640 189134 149696
rect 189630 149640 189686 149696
rect 188986 147736 189042 147792
rect 188894 131416 188950 131472
rect 189170 134564 189226 134600
rect 189170 134544 189172 134564
rect 189172 134544 189224 134564
rect 189224 134544 189226 134564
rect 186318 89664 186374 89720
rect 187698 93064 187754 93120
rect 187698 87896 187754 87952
rect 191562 266056 191618 266112
rect 191746 264988 191802 265024
rect 191746 264968 191748 264988
rect 191748 264968 191800 264988
rect 191800 264968 191802 264988
rect 191746 263880 191802 263936
rect 191746 262792 191802 262848
rect 191562 261704 191618 261760
rect 191746 259528 191802 259584
rect 191654 252592 191710 252648
rect 191562 250824 191618 250880
rect 191746 251912 191802 251968
rect 191654 249736 191710 249792
rect 191194 238584 191250 238640
rect 191746 247560 191802 247616
rect 191746 243208 191802 243264
rect 192022 240080 192078 240136
rect 192022 237904 192078 237960
rect 192482 179968 192538 180024
rect 192482 165688 192538 165744
rect 190458 162152 190514 162208
rect 191838 159296 191894 159352
rect 193126 162016 193182 162072
rect 192574 159296 192630 159352
rect 191746 149096 191802 149152
rect 189814 136720 189870 136776
rect 191654 145832 191710 145888
rect 191654 145560 191710 145616
rect 191102 144200 191158 144256
rect 191102 137808 191158 137864
rect 190458 134680 190514 134736
rect 190366 129784 190422 129840
rect 190274 125704 190330 125760
rect 191010 120264 191066 120320
rect 191562 136312 191618 136368
rect 191562 135496 191618 135552
rect 191194 133864 191250 133920
rect 191746 129240 191802 129296
rect 191654 128424 191710 128480
rect 191746 127608 191802 127664
rect 191562 126520 191618 126576
rect 193034 147872 193090 147928
rect 192942 146920 192998 146976
rect 192850 139848 192906 139904
rect 192482 124888 192538 124944
rect 193034 138216 193090 138272
rect 192942 123800 192998 123856
rect 191746 122984 191802 123040
rect 191746 122168 191802 122224
rect 191194 121372 191250 121408
rect 191194 121352 191196 121372
rect 191196 121352 191248 121372
rect 191248 121352 191250 121372
rect 191746 119448 191802 119504
rect 191746 118632 191802 118688
rect 191102 117544 191158 117600
rect 191562 116728 191618 116784
rect 189814 116456 189870 116512
rect 189722 115912 189778 115968
rect 189078 110744 189134 110800
rect 188434 107752 188490 107808
rect 189078 93200 189134 93256
rect 188802 93064 188858 93120
rect 189078 92520 189134 92576
rect 189814 99592 189870 99648
rect 190182 99456 190238 99512
rect 189722 89392 189778 89448
rect 188434 78512 188490 78568
rect 188342 73072 188398 73128
rect 186962 70216 187018 70272
rect 190274 92520 190330 92576
rect 190642 109656 190698 109712
rect 190826 106936 190882 106992
rect 191194 106120 191250 106176
rect 191010 103400 191066 103456
rect 191102 93608 191158 93664
rect 191102 92520 191158 92576
rect 191746 115096 191802 115152
rect 191838 114008 191894 114064
rect 191746 113192 191802 113248
rect 191746 112412 191748 112432
rect 191748 112412 191800 112432
rect 191800 112412 191802 112432
rect 191746 112376 191802 112412
rect 191746 110472 191802 110528
rect 191746 108876 191748 108896
rect 191748 108876 191800 108896
rect 191800 108876 191802 108896
rect 191746 108840 191802 108876
rect 191746 105032 191802 105088
rect 191746 101496 191802 101552
rect 191654 100680 191710 100736
rect 191654 99456 191710 99512
rect 191746 97960 191802 98016
rect 191654 97144 191710 97200
rect 191654 95784 191710 95840
rect 191746 94424 191802 94480
rect 193678 242800 193734 242856
rect 193310 240080 193366 240136
rect 198094 242020 198096 242040
rect 198096 242020 198148 242040
rect 198148 242020 198150 242040
rect 193862 174528 193918 174584
rect 193862 153720 193918 153776
rect 194598 142432 194654 142488
rect 193218 140800 193274 140856
rect 196070 238040 196126 238096
rect 195978 225528 196034 225584
rect 197358 234368 197414 234424
rect 196622 215872 196678 215928
rect 197358 193840 197414 193896
rect 195242 141072 195298 141128
rect 196530 146376 196586 146432
rect 196806 168952 196862 169008
rect 196714 142296 196770 142352
rect 198094 241984 198150 242020
rect 242990 242020 242992 242040
rect 242992 242020 243044 242040
rect 243044 242020 243046 242040
rect 242990 241984 243046 242020
rect 200118 166912 200174 166968
rect 200670 166912 200726 166968
rect 198830 149640 198886 149696
rect 197910 144744 197966 144800
rect 200210 157936 200266 157992
rect 207662 241032 207718 241088
rect 204902 226888 204958 226944
rect 201314 144064 201370 144120
rect 204350 151952 204406 152008
rect 202878 142160 202934 142216
rect 203890 142160 203946 142216
rect 207018 232464 207074 232520
rect 207018 229064 207074 229120
rect 204994 153720 205050 153776
rect 212446 240896 212502 240952
rect 210422 236544 210478 236600
rect 210514 229064 210570 229120
rect 210422 227568 210478 227624
rect 207662 156168 207718 156224
rect 204902 145696 204958 145752
rect 207018 148008 207074 148064
rect 208398 162696 208454 162752
rect 207754 149640 207810 149696
rect 207662 141480 207718 141536
rect 208490 152360 208546 152416
rect 207846 141344 207902 141400
rect 208122 141344 208178 141400
rect 194966 140392 195022 140448
rect 206558 140800 206614 140856
rect 210422 226344 210478 226400
rect 211066 226344 211122 226400
rect 210422 175344 210478 175400
rect 209134 171672 209190 171728
rect 210422 155896 210478 155952
rect 210514 155352 210570 155408
rect 209042 140528 209098 140584
rect 210514 144064 210570 144120
rect 211802 192480 211858 192536
rect 211158 153720 211214 153776
rect 211066 148416 211122 148472
rect 213182 216688 213238 216744
rect 214654 200640 214710 200696
rect 211894 158752 211950 158808
rect 212446 158752 212502 158808
rect 211802 151952 211858 152008
rect 211894 151000 211950 151056
rect 212354 142432 212410 142488
rect 210146 140564 210148 140584
rect 210148 140564 210200 140584
rect 210200 140564 210202 140584
rect 210146 140528 210202 140564
rect 217322 231104 217378 231160
rect 217322 217912 217378 217968
rect 217322 172488 217378 172544
rect 216678 168952 216734 169008
rect 215298 148280 215354 148336
rect 215850 143656 215906 143712
rect 218242 142160 218298 142216
rect 220082 208256 220138 208312
rect 219438 167048 219494 167104
rect 220174 167048 220230 167104
rect 220174 150456 220230 150512
rect 222198 141072 222254 141128
rect 223578 157392 223634 157448
rect 222842 144744 222898 144800
rect 222842 141480 222898 141536
rect 223210 141072 223266 141128
rect 224774 157392 224830 157448
rect 224498 144220 224554 144256
rect 224498 144200 224500 144220
rect 224500 144200 224552 144220
rect 224552 144200 224554 144220
rect 224222 142296 224278 142352
rect 223394 140800 223450 140856
rect 222842 140664 222898 140720
rect 215390 140528 215446 140584
rect 193402 140140 193458 140176
rect 193402 140120 193404 140140
rect 193404 140120 193456 140140
rect 193456 140120 193458 140140
rect 193218 131824 193274 131880
rect 193218 131416 193274 131472
rect 225050 129648 225106 129704
rect 225142 114824 225198 114880
rect 225050 113736 225106 113792
rect 193218 104216 193274 104272
rect 193126 102584 193182 102640
rect 193126 92520 193182 92576
rect 199198 93336 199254 93392
rect 208950 93336 209006 93392
rect 213274 93064 213330 93120
rect 193218 73752 193274 73808
rect 196530 92384 196586 92440
rect 198002 92384 198058 92440
rect 197082 86808 197138 86864
rect 200762 92112 200818 92168
rect 200210 91024 200266 91080
rect 200946 91024 201002 91080
rect 203706 90480 203762 90536
rect 204442 90344 204498 90400
rect 203706 88032 203762 88088
rect 206098 92384 206154 92440
rect 205546 92112 205602 92168
rect 205638 90208 205694 90264
rect 206834 90208 206890 90264
rect 202878 77832 202934 77888
rect 203522 77832 203578 77888
rect 203522 77152 203578 77208
rect 209226 88168 209282 88224
rect 210330 89664 210386 89720
rect 211618 89664 211674 89720
rect 209870 81368 209926 81424
rect 211066 81368 211122 81424
rect 211066 80688 211122 80744
rect 215298 90208 215354 90264
rect 215206 89528 215262 89584
rect 212538 71712 212594 71768
rect 212538 70352 212594 70408
rect 213182 70352 213238 70408
rect 216402 90208 216458 90264
rect 219162 91024 219218 91080
rect 219438 90344 219494 90400
rect 219162 85312 219218 85368
rect 220082 91024 220138 91080
rect 219806 89528 219862 89584
rect 220082 82728 220138 82784
rect 224314 91024 224370 91080
rect 222290 67496 222346 67552
rect 225050 109112 225106 109168
rect 225142 94696 225198 94752
rect 230478 238584 230534 238640
rect 226154 114824 226210 114880
rect 226430 171672 226486 171728
rect 226430 134680 226486 134736
rect 226614 146512 226670 146568
rect 226706 139032 226762 139088
rect 226706 137128 226762 137184
rect 226614 136584 226670 136640
rect 226706 135496 226762 135552
rect 226614 134680 226670 134736
rect 226706 133628 226708 133648
rect 226708 133628 226760 133648
rect 226760 133628 226762 133648
rect 226706 133592 226762 133628
rect 226614 132776 226670 132832
rect 226706 131960 226762 132016
rect 226706 130872 226762 130928
rect 226798 130056 226854 130112
rect 226614 128968 226670 129024
rect 226430 128424 226486 128480
rect 226706 127336 226762 127392
rect 226706 126520 226762 126576
rect 226614 124616 226670 124672
rect 227626 123800 227682 123856
rect 226706 122984 226762 123040
rect 226522 122168 226578 122224
rect 226706 120264 226762 120320
rect 226522 118360 226578 118416
rect 226614 117544 226670 117600
rect 227626 116728 227682 116784
rect 226706 115948 226708 115968
rect 226708 115948 226760 115968
rect 226760 115948 226762 115968
rect 226706 115912 226762 115948
rect 226430 114008 226486 114064
rect 226338 112104 226394 112160
rect 226338 110472 226394 110528
rect 226338 105848 226394 105904
rect 226338 101496 226394 101552
rect 226338 99456 226394 99512
rect 226706 111288 226762 111344
rect 226522 108568 226578 108624
rect 226706 106936 226762 106992
rect 226706 105052 226762 105088
rect 226706 105032 226708 105052
rect 226708 105032 226760 105052
rect 226760 105032 226762 105052
rect 226706 104216 226762 104272
rect 226706 103400 226762 103456
rect 226706 102312 226762 102368
rect 226706 98776 226762 98832
rect 226614 97960 226670 98016
rect 226430 95104 226486 95160
rect 226706 96056 226762 96112
rect 226982 97144 227038 97200
rect 227074 95104 227130 95160
rect 225050 89392 225106 89448
rect 226706 84088 226762 84144
rect 224866 4800 224922 4856
rect 227166 93608 227222 93664
rect 229098 162832 229154 162888
rect 231858 228792 231914 228848
rect 236642 232464 236698 232520
rect 231858 227704 231914 227760
rect 233146 227704 233202 227760
rect 230478 162016 230534 162072
rect 227994 144880 228050 144936
rect 227902 129240 227958 129296
rect 227902 126928 227958 126984
rect 228362 139848 228418 139904
rect 227902 125704 227958 125760
rect 230478 158752 230534 158808
rect 227902 100680 227958 100736
rect 227994 95240 228050 95296
rect 227994 75792 228050 75848
rect 236642 220768 236698 220824
rect 235998 210296 236054 210352
rect 231950 153040 232006 153096
rect 232502 153040 232558 153096
rect 231950 151816 232006 151872
rect 233238 150592 233294 150648
rect 232502 142296 232558 142352
rect 231858 77832 231914 77888
rect 231122 73072 231178 73128
rect 232594 77832 232650 77888
rect 235998 169768 236054 169824
rect 235998 138896 236054 138952
rect 237378 164328 237434 164384
rect 238022 140800 238078 140856
rect 240230 154400 240286 154456
rect 240230 153176 240286 153232
rect 244922 241032 244978 241088
rect 242254 239944 242310 240000
rect 242714 239944 242770 240000
rect 241426 224168 241482 224224
rect 240782 154400 240838 154456
rect 240322 149096 240378 149152
rect 240782 149096 240838 149152
rect 239402 90344 239458 90400
rect 226982 3304 227038 3360
rect 244922 217912 244978 217968
rect 247498 239400 247554 239456
rect 247774 238040 247830 238096
rect 246394 236816 246450 236872
rect 245106 146920 245162 146976
rect 246394 199280 246450 199336
rect 249154 239400 249210 239456
rect 250166 241984 250222 242040
rect 249890 236544 249946 236600
rect 249890 160112 249946 160168
rect 251822 239808 251878 239864
rect 251822 238584 251878 238640
rect 252098 232464 252154 232520
rect 252834 297608 252890 297664
rect 252834 293392 252890 293448
rect 252558 220904 252614 220960
rect 252190 145560 252246 145616
rect 253938 300600 253994 300656
rect 253018 298832 253074 298888
rect 253018 297608 253074 297664
rect 253938 296520 253994 296576
rect 254030 295568 254086 295624
rect 254582 301688 254638 301744
rect 254214 299784 254270 299840
rect 254122 293120 254178 293176
rect 252834 265512 252890 265568
rect 253846 265240 253902 265296
rect 252834 258712 252890 258768
rect 258170 475360 258226 475416
rect 256882 403960 256938 404016
rect 255318 300328 255374 300384
rect 255318 297744 255374 297800
rect 255318 287544 255374 287600
rect 256606 298172 256662 298208
rect 256606 298152 256608 298172
rect 256608 298152 256660 298172
rect 256660 298152 256662 298172
rect 255594 296112 255650 296168
rect 256606 296112 256662 296168
rect 256330 294752 256386 294808
rect 256606 294344 256662 294400
rect 256146 293140 256202 293176
rect 256146 293120 256148 293140
rect 256148 293120 256200 293140
rect 256200 293120 256202 293140
rect 255962 292576 256018 292632
rect 255962 291760 256018 291816
rect 255686 291624 255742 291680
rect 256606 291080 256662 291136
rect 255502 289992 255558 290048
rect 255502 289176 255558 289232
rect 255502 287952 255558 288008
rect 258354 521600 258410 521656
rect 258906 395256 258962 395312
rect 259550 526360 259606 526416
rect 261022 529080 261078 529136
rect 261022 452920 261078 452976
rect 261114 446392 261170 446448
rect 261114 384784 261170 384840
rect 263598 389000 263654 389056
rect 262402 388320 262458 388376
rect 262310 370640 262366 370696
rect 262218 357992 262274 358048
rect 258722 324944 258778 325000
rect 258170 290808 258226 290864
rect 257434 287000 257490 287056
rect 255410 286628 255412 286648
rect 255412 286628 255464 286648
rect 255464 286628 255466 286648
rect 255410 286592 255466 286628
rect 257434 286456 257490 286512
rect 255502 286184 255558 286240
rect 256698 286048 256754 286104
rect 255410 285368 255466 285424
rect 255410 284008 255466 284064
rect 255502 283192 255558 283248
rect 255410 282376 255466 282432
rect 255502 281968 255558 282024
rect 255410 281444 255466 281480
rect 255410 281424 255412 281444
rect 255412 281424 255464 281444
rect 255464 281424 255466 281444
rect 255502 280200 255558 280256
rect 255502 278976 255558 279032
rect 255502 278432 255558 278488
rect 255410 277616 255466 277672
rect 255502 277344 255558 277400
rect 255502 276800 255558 276856
rect 255594 276392 255650 276448
rect 255410 275984 255466 276040
rect 255502 275032 255558 275088
rect 255410 274660 255412 274680
rect 255412 274660 255464 274680
rect 255464 274660 255466 274680
rect 255410 274624 255466 274660
rect 255410 274252 255412 274272
rect 255412 274252 255464 274272
rect 255464 274252 255466 274272
rect 255410 274216 255466 274252
rect 255502 273808 255558 273864
rect 255410 272448 255466 272504
rect 255410 272040 255466 272096
rect 255502 271224 255558 271280
rect 255410 269864 255466 269920
rect 255410 269456 255466 269512
rect 255410 268232 255466 268288
rect 255410 267824 255466 267880
rect 255410 266872 255466 266928
rect 255318 266056 255374 266112
rect 255502 264288 255558 264344
rect 255410 263880 255466 263936
rect 255502 263472 255558 263528
rect 255686 263472 255742 263528
rect 255686 262656 255742 262712
rect 255410 262248 255466 262304
rect 255502 261296 255558 261352
rect 255410 260480 255466 260536
rect 256422 260072 256478 260128
rect 255410 259664 255466 259720
rect 255502 259256 255558 259312
rect 255594 258304 255650 258360
rect 255410 257896 255466 257952
rect 255410 256264 255466 256320
rect 255318 255312 255374 255368
rect 254030 253680 254086 253736
rect 253938 252456 253994 252512
rect 252834 242800 252890 242856
rect 252926 242392 252982 242448
rect 254582 241440 254638 241496
rect 254582 240760 254638 240816
rect 253938 237904 253994 237960
rect 252834 236816 252890 236872
rect 253938 235728 253994 235784
rect 253938 233008 253994 233064
rect 254674 228928 254730 228984
rect 255502 254904 255558 254960
rect 255410 254532 255412 254552
rect 255412 254532 255464 254552
rect 255464 254532 255466 254552
rect 255410 254496 255466 254532
rect 255410 253272 255466 253328
rect 255410 251912 255466 251968
rect 255502 251504 255558 251560
rect 255502 251096 255558 251152
rect 255410 250688 255466 250744
rect 255410 249872 255466 249928
rect 256422 253136 256478 253192
rect 255594 249736 255650 249792
rect 255502 249328 255558 249384
rect 255410 248920 255466 248976
rect 255410 248376 255466 248432
rect 255502 248104 255558 248160
rect 255502 247152 255558 247208
rect 255686 246744 255742 246800
rect 255502 246200 255558 246256
rect 255594 245928 255650 245984
rect 255502 245556 255504 245576
rect 255504 245556 255556 245576
rect 255556 245556 255558 245576
rect 255502 245520 255558 245556
rect 255686 245112 255742 245168
rect 255594 244704 255650 244760
rect 255502 244160 255558 244216
rect 255594 243480 255650 243536
rect 255778 243616 255834 243672
rect 255594 242120 255650 242176
rect 255502 241712 255558 241768
rect 255778 241440 255834 241496
rect 255410 235728 255466 235784
rect 255318 225528 255374 225584
rect 255318 174528 255374 174584
rect 254582 89528 254638 89584
rect 256790 269048 256846 269104
rect 256882 257488 256938 257544
rect 257526 246336 257582 246392
rect 258538 299920 258594 299976
rect 258814 293800 258870 293856
rect 258446 278160 258502 278216
rect 258262 275440 258318 275496
rect 257526 238040 257582 238096
rect 257342 237360 257398 237416
rect 256882 233144 256938 233200
rect 258262 236000 258318 236056
rect 258446 237360 258502 237416
rect 258262 222128 258318 222184
rect 259366 281560 259422 281616
rect 259274 281016 259330 281072
rect 259458 279384 259514 279440
rect 259458 278024 259514 278080
rect 259642 292168 259698 292224
rect 259366 268640 259422 268696
rect 258170 204312 258226 204368
rect 258722 204312 258778 204368
rect 258078 94696 258134 94752
rect 260838 295160 260894 295216
rect 260746 291760 260802 291816
rect 260746 289756 260748 289776
rect 260748 289756 260800 289776
rect 260800 289756 260802 289776
rect 260746 289720 260802 289756
rect 259826 279792 259882 279848
rect 260930 266464 260986 266520
rect 262218 291624 262274 291680
rect 260930 235864 260986 235920
rect 260930 205692 260986 205728
rect 260930 205672 260932 205692
rect 260932 205672 260984 205692
rect 260984 205672 260986 205692
rect 259550 156032 259606 156088
rect 259458 128968 259514 129024
rect 258170 91024 258226 91080
rect 254674 4800 254730 4856
rect 262402 284960 262458 285016
rect 262402 284280 262458 284336
rect 263966 284280 264022 284336
rect 262402 271496 262458 271552
rect 262402 271088 262458 271144
rect 263690 262928 263746 262984
rect 263598 260072 263654 260128
rect 262770 257080 262826 257136
rect 262494 253272 262550 253328
rect 263506 254224 263562 254280
rect 263598 253952 263654 254008
rect 263598 246336 263654 246392
rect 260930 89664 260986 89720
rect 262218 79328 262274 79384
rect 263874 246200 263930 246256
rect 263874 224168 263930 224224
rect 265622 454144 265678 454200
rect 265162 383560 265218 383616
rect 265162 382336 265218 382392
rect 264978 318008 265034 318064
rect 264978 283464 265034 283520
rect 266358 335960 266414 336016
rect 265254 322088 265310 322144
rect 265070 280744 265126 280800
rect 264978 279384 265034 279440
rect 264334 278840 264390 278896
rect 266450 319368 266506 319424
rect 266450 316104 266506 316160
rect 265254 267144 265310 267200
rect 265254 265648 265310 265704
rect 265622 265648 265678 265704
rect 266634 361664 266690 361720
rect 267922 449928 267978 449984
rect 266634 301008 266690 301064
rect 266542 284824 266598 284880
rect 266450 282648 266506 282704
rect 266542 263064 266598 263120
rect 266450 259664 266506 259720
rect 266450 258032 266506 258088
rect 266450 251932 266506 251968
rect 266450 251912 266452 251932
rect 266452 251912 266504 251932
rect 266504 251912 266506 251932
rect 267830 320048 267886 320104
rect 268382 376624 268438 376680
rect 269394 460944 269450 461000
rect 269210 322904 269266 322960
rect 267922 319404 267924 319424
rect 267924 319404 267976 319424
rect 267976 319404 267978 319424
rect 267922 319368 267978 319404
rect 267830 309712 267886 309768
rect 267738 286456 267794 286512
rect 266726 214512 266782 214568
rect 264242 95784 264298 95840
rect 265346 3304 265402 3360
rect 269118 303864 269174 303920
rect 268014 295160 268070 295216
rect 268106 288360 268162 288416
rect 268106 240488 268162 240544
rect 269210 288360 269266 288416
rect 269762 441632 269818 441688
rect 269486 312432 269542 312488
rect 269302 269184 269358 269240
rect 270682 451560 270738 451616
rect 270774 360168 270830 360224
rect 270774 311888 270830 311944
rect 270498 307672 270554 307728
rect 270590 299784 270646 299840
rect 270498 273536 270554 273592
rect 269394 265512 269450 265568
rect 270958 273536 271014 273592
rect 271142 269048 271198 269104
rect 273258 452376 273314 452432
rect 273074 451288 273130 451344
rect 271970 243480 272026 243536
rect 271878 226888 271934 226944
rect 273442 533296 273498 533352
rect 273534 459584 273590 459640
rect 273442 452648 273498 452704
rect 274730 382200 274786 382256
rect 273442 298016 273498 298072
rect 273442 296792 273498 296848
rect 273442 281560 273498 281616
rect 273350 271088 273406 271144
rect 272522 247424 272578 247480
rect 272522 247016 272578 247072
rect 272154 246200 272210 246256
rect 270498 162696 270554 162752
rect 269118 73752 269174 73808
rect 273534 276664 273590 276720
rect 273442 213152 273498 213208
rect 273534 153720 273590 153776
rect 274730 261024 274786 261080
rect 275006 293800 275062 293856
rect 275006 292576 275062 292632
rect 275282 267144 275338 267200
rect 275282 256944 275338 257000
rect 277490 458768 277546 458824
rect 277398 348336 277454 348392
rect 277398 317464 277454 317520
rect 276202 292576 276258 292632
rect 276018 238584 276074 238640
rect 273258 86128 273314 86184
rect 277398 276664 277454 276720
rect 277766 458768 277822 458824
rect 277582 306448 277638 306504
rect 276294 264288 276350 264344
rect 276294 263608 276350 263664
rect 277490 243616 277546 243672
rect 278778 452784 278834 452840
rect 277766 317464 277822 317520
rect 278318 262112 278374 262168
rect 278318 261296 278374 261352
rect 280158 463664 280214 463720
rect 278870 340040 278926 340096
rect 278870 296792 278926 296848
rect 280434 416744 280490 416800
rect 280250 387640 280306 387696
rect 280250 369688 280306 369744
rect 281446 387640 281502 387696
rect 281538 380840 281594 380896
rect 280526 325760 280582 325816
rect 281630 286320 281686 286376
rect 281538 283464 281594 283520
rect 280342 256672 280398 256728
rect 280158 235728 280214 235784
rect 282918 313928 282974 313984
rect 281814 304136 281870 304192
rect 281722 152360 281778 152416
rect 281630 126928 281686 126984
rect 283102 386008 283158 386064
rect 283194 279384 283250 279440
rect 288622 604424 288678 604480
rect 289726 604460 289728 604480
rect 289728 604460 289780 604480
rect 289780 604460 289782 604480
rect 289726 604424 289782 604460
rect 285586 536696 285642 536752
rect 285586 536016 285642 536072
rect 284390 390496 284446 390552
rect 284390 389136 284446 389192
rect 284390 385600 284446 385656
rect 285770 302368 285826 302424
rect 284942 298696 284998 298752
rect 285678 291760 285734 291816
rect 284942 133456 284998 133512
rect 284390 88032 284446 88088
rect 287058 452512 287114 452568
rect 287058 450472 287114 450528
rect 285954 264288 286010 264344
rect 287242 467880 287298 467936
rect 287150 268368 287206 268424
rect 287058 242800 287114 242856
rect 285954 144064 286010 144120
rect 288438 459720 288494 459776
rect 287334 455504 287390 455560
rect 288346 455504 288402 455560
rect 287426 418240 287482 418296
rect 288530 452512 288586 452568
rect 288530 267008 288586 267064
rect 288438 264152 288494 264208
rect 289818 456864 289874 456920
rect 288622 261432 288678 261488
rect 288530 250416 288586 250472
rect 288530 224848 288586 224904
rect 288438 157936 288494 157992
rect 291198 375264 291254 375320
rect 291198 301552 291254 301608
rect 289818 147736 289874 147792
rect 292578 366968 292634 367024
rect 294050 470600 294106 470656
rect 291290 272448 291346 272504
rect 582470 697176 582526 697232
rect 582378 617480 582434 617536
rect 295430 536016 295486 536072
rect 294050 320184 294106 320240
rect 292670 278024 292726 278080
rect 582378 590960 582434 591016
rect 295430 310528 295486 310584
rect 295338 309168 295394 309224
rect 294050 155896 294106 155952
rect 294694 155896 294750 155952
rect 291842 82048 291898 82104
rect 299478 465160 299534 465216
rect 298190 458224 298246 458280
rect 298282 331744 298338 331800
rect 296810 253136 296866 253192
rect 299570 462304 299626 462360
rect 299662 307808 299718 307864
rect 299570 305632 299626 305688
rect 299478 298696 299534 298752
rect 291842 3304 291898 3360
rect 582378 577632 582434 577688
rect 582562 683848 582618 683904
rect 582654 644000 582710 644056
rect 582746 630808 582802 630864
rect 582930 670656 582986 670712
rect 582746 607824 582802 607880
rect 582654 603608 582710 603664
rect 582378 537784 582434 537840
rect 580170 484608 580226 484664
rect 580170 458088 580226 458144
rect 582838 564304 582894 564360
rect 582746 524456 582802 524512
rect 582654 511264 582710 511320
rect 582470 471416 582526 471472
rect 580262 418240 580318 418296
rect 582378 378392 582434 378448
rect 582470 365064 582526 365120
rect 580906 325216 580962 325272
rect 582378 302232 582434 302288
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580722 258848 580778 258904
rect 304262 250416 304318 250472
rect 580170 232328 580226 232384
rect 580262 219000 580318 219056
rect 580354 205672 580410 205728
rect 302238 205536 302294 205592
rect 579986 192480 580042 192536
rect 580170 179152 580226 179208
rect 301962 3304 302018 3360
rect 306378 40568 306434 40624
rect 317418 133048 317474 133104
rect 310518 84768 310574 84824
rect 323582 142160 323638 142216
rect 334622 91704 334678 91760
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 46280 580226 46336
rect 582746 431568 582802 431624
rect 582654 404912 582710 404968
rect 582746 390496 582802 390552
rect 582562 351872 582618 351928
rect 582654 312024 582710 312080
rect 582562 289856 582618 289912
rect 582470 252456 582526 252512
rect 582470 245520 582526 245576
rect 582654 236000 582710 236056
rect 582838 165824 582894 165880
rect 582654 152632 582710 152688
rect 582930 150456 582986 150512
rect 583022 139304 583078 139360
rect 583114 125976 583170 126032
rect 582930 112784 582986 112840
rect 582838 87488 582894 87544
rect 582746 59608 582802 59664
rect 582654 19760 582710 19816
rect 582930 80688 582986 80744
rect 583022 72936 583078 72992
rect 582930 33088 582986 33144
rect 582838 6568 582894 6624
<< metal3 >>
rect 72969 699820 73035 699821
rect 72918 699818 72924 699820
rect 72878 699758 72924 699818
rect 72988 699816 73035 699820
rect 73030 699760 73035 699816
rect 72918 699756 72924 699758
rect 72988 699756 73035 699760
rect 72969 699755 73035 699756
rect -960 697220 480 697460
rect 582465 697234 582531 697237
rect 583520 697234 584960 697324
rect 582465 697232 584960 697234
rect 582465 697176 582470 697232
rect 582526 697176 584960 697232
rect 582465 697174 584960 697176
rect 582465 697171 582531 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582557 683906 582623 683909
rect 583520 683906 584960 683996
rect 582557 683904 584960 683906
rect 582557 683848 582562 683904
rect 582618 683848 584960 683904
rect 582557 683846 584960 683848
rect 582557 683843 582623 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582925 670714 582991 670717
rect 583520 670714 584960 670804
rect 582925 670712 584960 670714
rect 582925 670656 582930 670712
rect 582986 670656 584960 670712
rect 582925 670654 584960 670656
rect 582925 670651 582991 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582649 644058 582715 644061
rect 583520 644058 584960 644148
rect 582649 644056 584960 644058
rect 582649 644000 582654 644056
rect 582710 644000 584960 644056
rect 582649 643998 584960 644000
rect 582649 643995 582715 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582741 630866 582807 630869
rect 583520 630866 584960 630956
rect 582741 630864 584960 630866
rect 582741 630808 582746 630864
rect 582802 630808 584960 630864
rect 582741 630806 584960 630808
rect 582741 630803 582807 630806
rect 583520 630716 584960 630806
rect 162710 619652 162716 619716
rect 162780 619714 162786 619716
rect 227713 619714 227779 619717
rect 162780 619712 227779 619714
rect 162780 619656 227718 619712
rect 227774 619656 227779 619712
rect 162780 619654 227779 619656
rect 162780 619652 162786 619654
rect 227713 619651 227779 619654
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582373 617538 582439 617541
rect 583520 617538 584960 617628
rect 582373 617536 584960 617538
rect 582373 617480 582378 617536
rect 582434 617480 584960 617536
rect 582373 617478 584960 617480
rect 582373 617475 582439 617478
rect 583520 617388 584960 617478
rect 180006 609996 180012 610060
rect 180076 610058 180082 610060
rect 207657 610058 207723 610061
rect 180076 610056 207723 610058
rect 180076 610000 207662 610056
rect 207718 610000 207723 610056
rect 180076 609998 207723 610000
rect 180076 609996 180082 609998
rect 207657 609995 207723 609998
rect 184054 608772 184060 608836
rect 184124 608834 184130 608836
rect 208393 608834 208459 608837
rect 184124 608832 208459 608834
rect 184124 608776 208398 608832
rect 208454 608776 208459 608832
rect 184124 608774 208459 608776
rect 184124 608772 184130 608774
rect 208393 608771 208459 608774
rect 175181 608698 175247 608701
rect 226425 608698 226491 608701
rect 175181 608696 226491 608698
rect 175181 608640 175186 608696
rect 175242 608640 226430 608696
rect 226486 608640 226491 608696
rect 175181 608638 226491 608640
rect 175181 608635 175247 608638
rect 226425 608635 226491 608638
rect 191649 607882 191715 607885
rect 582741 607882 582807 607885
rect 191649 607880 582807 607882
rect 191649 607824 191654 607880
rect 191710 607824 582746 607880
rect 582802 607824 582807 607880
rect 191649 607822 582807 607824
rect 191649 607819 191715 607822
rect 582741 607819 582807 607822
rect 192334 607276 192340 607340
rect 192404 607338 192410 607340
rect 209405 607338 209471 607341
rect 192404 607336 209471 607338
rect 192404 607280 209410 607336
rect 209466 607280 209471 607336
rect 192404 607278 209471 607280
rect 192404 607276 192410 607278
rect 209405 607275 209471 607278
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 189717 605978 189783 605981
rect 222101 605978 222167 605981
rect 189717 605976 222167 605978
rect 189717 605920 189722 605976
rect 189778 605920 222106 605976
rect 222162 605920 222167 605976
rect 189717 605918 222167 605920
rect 189717 605915 189783 605918
rect 222101 605915 222167 605918
rect 180701 604618 180767 604621
rect 234061 604618 234127 604621
rect 180701 604616 234127 604618
rect 180701 604560 180706 604616
rect 180762 604560 234066 604616
rect 234122 604560 234127 604616
rect 180701 604558 234127 604560
rect 180701 604555 180767 604558
rect 234061 604555 234127 604558
rect 188429 604482 188495 604485
rect 196709 604482 196775 604485
rect 288617 604482 288683 604485
rect 289721 604482 289787 604485
rect 188429 604480 289787 604482
rect 188429 604424 188434 604480
rect 188490 604424 196714 604480
rect 196770 604424 288622 604480
rect 288678 604424 289726 604480
rect 289782 604424 289787 604480
rect 188429 604422 289787 604424
rect 188429 604419 188495 604422
rect 196709 604419 196775 604422
rect 288617 604419 288683 604422
rect 289721 604419 289787 604422
rect 583520 604060 584960 604300
rect 191741 603666 191807 603669
rect 582649 603666 582715 603669
rect 191741 603664 582715 603666
rect 191741 603608 191746 603664
rect 191802 603608 582654 603664
rect 582710 603608 582715 603664
rect 191741 603606 582715 603608
rect 191741 603603 191807 603606
rect 582649 603603 582715 603606
rect 88977 603258 89043 603261
rect 230105 603258 230171 603261
rect 88977 603256 230171 603258
rect 88977 603200 88982 603256
rect 89038 603200 230110 603256
rect 230166 603200 230171 603256
rect 88977 603198 230171 603200
rect 88977 603195 89043 603198
rect 230105 603195 230171 603198
rect 226333 603122 226399 603125
rect 258390 603122 258396 603124
rect 226333 603120 258396 603122
rect 226333 603064 226338 603120
rect 226394 603064 258396 603120
rect 226333 603062 258396 603064
rect 226333 603059 226399 603062
rect 258390 603060 258396 603062
rect 258460 603060 258466 603124
rect 171041 602034 171107 602037
rect 201125 602034 201191 602037
rect 171041 602032 201191 602034
rect 171041 601976 171046 602032
rect 171102 601976 201130 602032
rect 201186 601976 201191 602032
rect 171041 601974 201191 601976
rect 171041 601971 171107 601974
rect 201125 601971 201191 601974
rect 194133 601898 194199 601901
rect 204805 601898 204871 601901
rect 194133 601896 204871 601898
rect 194133 601840 194138 601896
rect 194194 601840 204810 601896
rect 204866 601840 204871 601896
rect 194133 601838 204871 601840
rect 194133 601835 194199 601838
rect 204805 601835 204871 601838
rect 230105 601898 230171 601901
rect 244590 601898 244596 601900
rect 230105 601896 244596 601898
rect 230105 601840 230110 601896
rect 230166 601840 244596 601896
rect 230105 601838 244596 601840
rect 230105 601835 230171 601838
rect 244590 601836 244596 601838
rect 244660 601836 244666 601900
rect 239213 601762 239279 601765
rect 259494 601762 259500 601764
rect 239213 601760 259500 601762
rect 239213 601704 239218 601760
rect 239274 601704 259500 601760
rect 239213 601702 259500 601704
rect 239213 601699 239279 601702
rect 259494 601700 259500 601702
rect 259564 601700 259570 601764
rect 154430 600884 154436 600948
rect 154500 600946 154506 600948
rect 194133 600946 194199 600949
rect 154500 600944 194199 600946
rect 154500 600888 194138 600944
rect 194194 600888 194199 600944
rect 154500 600886 194199 600888
rect 154500 600884 154506 600886
rect 194133 600883 194199 600886
rect 192569 600810 192635 600813
rect 204253 600810 204319 600813
rect 192569 600808 204319 600810
rect 192569 600752 192574 600808
rect 192630 600752 204258 600808
rect 204314 600752 204319 600808
rect 192569 600750 204319 600752
rect 192569 600747 192635 600750
rect 204253 600747 204319 600750
rect 209957 600810 210023 600813
rect 219934 600810 219940 600812
rect 209957 600808 219940 600810
rect 209957 600752 209962 600808
rect 210018 600752 219940 600808
rect 209957 600750 219940 600752
rect 209957 600747 210023 600750
rect 219934 600748 219940 600750
rect 220004 600748 220010 600812
rect 186957 600674 187023 600677
rect 199837 600674 199903 600677
rect 186957 600672 199903 600674
rect 186957 600616 186962 600672
rect 187018 600616 199842 600672
rect 199898 600616 199903 600672
rect 186957 600614 199903 600616
rect 186957 600611 187023 600614
rect 199837 600611 199903 600614
rect 202413 600674 202479 600677
rect 232446 600674 232452 600676
rect 202413 600672 232452 600674
rect 202413 600616 202418 600672
rect 202474 600616 232452 600672
rect 202413 600614 232452 600616
rect 202413 600611 202479 600614
rect 232446 600612 232452 600614
rect 232516 600612 232522 600676
rect 244181 600674 244247 600677
rect 254761 600674 254827 600677
rect 244181 600672 254827 600674
rect 244181 600616 244186 600672
rect 244242 600616 254766 600672
rect 254822 600616 254827 600672
rect 244181 600614 254827 600616
rect 244181 600611 244247 600614
rect 254761 600611 254827 600614
rect 193438 600476 193444 600540
rect 193508 600538 193514 600540
rect 222929 600538 222995 600541
rect 193508 600536 222995 600538
rect 193508 600480 222934 600536
rect 222990 600480 222995 600536
rect 193508 600478 222995 600480
rect 193508 600476 193514 600478
rect 222929 600475 222995 600478
rect 231761 600538 231827 600541
rect 246205 600538 246271 600541
rect 231761 600536 246271 600538
rect 231761 600480 231766 600536
rect 231822 600480 246210 600536
rect 246266 600480 246271 600536
rect 231761 600478 246271 600480
rect 231761 600475 231827 600478
rect 246205 600475 246271 600478
rect 246757 600538 246823 600541
rect 263542 600538 263548 600540
rect 246757 600536 263548 600538
rect 246757 600480 246762 600536
rect 246818 600480 263548 600536
rect 246757 600478 263548 600480
rect 246757 600475 246823 600478
rect 263542 600476 263548 600478
rect 263612 600476 263618 600540
rect 215293 600404 215359 600405
rect 215293 600402 215340 600404
rect 215212 600400 215340 600402
rect 215404 600402 215410 600404
rect 216397 600402 216463 600405
rect 215404 600400 216463 600402
rect 215212 600344 215298 600400
rect 215404 600344 216402 600400
rect 216458 600344 216463 600400
rect 215212 600342 215340 600344
rect 215293 600340 215340 600342
rect 215404 600342 216463 600344
rect 215404 600340 215410 600342
rect 215293 600339 215359 600340
rect 216397 600339 216463 600342
rect 218237 600402 218303 600405
rect 218646 600402 218652 600404
rect 218237 600400 218652 600402
rect 218237 600344 218242 600400
rect 218298 600344 218652 600400
rect 218237 600342 218652 600344
rect 218237 600339 218303 600342
rect 218646 600340 218652 600342
rect 218716 600402 218722 600404
rect 219341 600402 219407 600405
rect 218716 600400 219407 600402
rect 218716 600344 219346 600400
rect 219402 600344 219407 600400
rect 218716 600342 219407 600344
rect 218716 600340 218722 600342
rect 219341 600339 219407 600342
rect 225781 600402 225847 600405
rect 230974 600402 230980 600404
rect 225781 600400 230980 600402
rect 225781 600344 225786 600400
rect 225842 600344 230980 600400
rect 225781 600342 230980 600344
rect 225781 600339 225847 600342
rect 230974 600340 230980 600342
rect 231044 600340 231050 600404
rect 250069 600402 250135 600405
rect 276238 600402 276244 600404
rect 250069 600400 276244 600402
rect 250069 600344 250074 600400
rect 250130 600344 276244 600400
rect 250069 600342 276244 600344
rect 250069 600339 250135 600342
rect 276238 600340 276244 600342
rect 276308 600340 276314 600404
rect 178769 599586 178835 599589
rect 205633 599586 205699 599589
rect 206829 599586 206895 599589
rect 178769 599584 206895 599586
rect 178769 599528 178774 599584
rect 178830 599528 205638 599584
rect 205694 599528 206834 599584
rect 206890 599528 206895 599584
rect 178769 599526 206895 599528
rect 178769 599523 178835 599526
rect 205633 599523 205699 599526
rect 206829 599523 206895 599526
rect 248321 599586 248387 599589
rect 254577 599586 254643 599589
rect 248321 599584 254643 599586
rect 248321 599528 248326 599584
rect 248382 599528 254582 599584
rect 254638 599528 254643 599584
rect 248321 599526 254643 599528
rect 248321 599523 248387 599526
rect 254577 599523 254643 599526
rect 192661 599450 192727 599453
rect 198549 599450 198615 599453
rect 212441 599452 212507 599453
rect 212390 599450 212396 599452
rect 192661 599448 198615 599450
rect 192661 599392 192666 599448
rect 192722 599392 198554 599448
rect 198610 599392 198615 599448
rect 192661 599390 198615 599392
rect 212350 599390 212396 599450
rect 212460 599448 212507 599452
rect 212502 599392 212507 599448
rect 192661 599387 192727 599390
rect 198549 599387 198615 599390
rect 212390 599388 212396 599390
rect 212460 599388 212507 599392
rect 212441 599387 212507 599388
rect 226333 599452 226399 599453
rect 226333 599448 226380 599452
rect 226444 599450 226450 599452
rect 236361 599450 236427 599453
rect 238518 599450 238524 599452
rect 226333 599392 226338 599448
rect 226333 599388 226380 599392
rect 226444 599390 226490 599450
rect 236361 599448 238524 599450
rect 236361 599392 236366 599448
rect 236422 599392 238524 599448
rect 236361 599390 238524 599392
rect 226444 599388 226450 599390
rect 226333 599387 226399 599388
rect 236361 599387 236427 599390
rect 238518 599388 238524 599390
rect 238588 599388 238594 599452
rect 75913 599314 75979 599317
rect 249333 599314 249399 599317
rect 75913 599312 249399 599314
rect 75913 599256 75918 599312
rect 75974 599256 249338 599312
rect 249394 599256 249399 599312
rect 75913 599254 249399 599256
rect 75913 599251 75979 599254
rect 249333 599251 249399 599254
rect 204437 599178 204503 599181
rect 204846 599178 204852 599180
rect 204437 599176 204852 599178
rect 204437 599120 204442 599176
rect 204498 599120 204852 599176
rect 204437 599118 204852 599120
rect 204437 599115 204503 599118
rect 204846 599116 204852 599118
rect 204916 599116 204922 599180
rect 213269 599178 213335 599181
rect 222694 599178 222700 599180
rect 213269 599176 222700 599178
rect 213269 599120 213274 599176
rect 213330 599120 222700 599176
rect 213269 599118 222700 599120
rect 213269 599115 213335 599118
rect 222694 599116 222700 599118
rect 222764 599116 222770 599180
rect 229686 599116 229692 599180
rect 229756 599178 229762 599180
rect 231209 599178 231275 599181
rect 229756 599176 231275 599178
rect 229756 599120 231214 599176
rect 231270 599120 231275 599176
rect 229756 599118 231275 599120
rect 229756 599116 229762 599118
rect 231209 599115 231275 599118
rect 236821 599178 236887 599181
rect 237414 599178 237420 599180
rect 236821 599176 237420 599178
rect 236821 599120 236826 599176
rect 236882 599120 237420 599176
rect 236821 599118 237420 599120
rect 236821 599115 236887 599118
rect 237414 599116 237420 599118
rect 237484 599116 237490 599180
rect 240041 599178 240107 599181
rect 241646 599178 241652 599180
rect 240041 599176 241652 599178
rect 240041 599120 240046 599176
rect 240102 599120 241652 599176
rect 240041 599118 241652 599120
rect 240041 599115 240107 599118
rect 241646 599116 241652 599118
rect 241716 599116 241722 599180
rect 243905 599178 243971 599181
rect 262254 599178 262260 599180
rect 243905 599176 262260 599178
rect 243905 599120 243910 599176
rect 243966 599120 262260 599176
rect 243905 599118 262260 599120
rect 243905 599115 243971 599118
rect 262254 599116 262260 599118
rect 262324 599116 262330 599180
rect 193121 599110 193187 599113
rect 193121 599108 193660 599110
rect 193121 599052 193126 599108
rect 193182 599052 193660 599108
rect 193121 599050 193660 599052
rect 193121 599047 193187 599050
rect 194593 599044 194659 599045
rect 197169 599044 197235 599045
rect 201585 599044 201651 599045
rect 203057 599044 203123 599045
rect 207105 599044 207171 599045
rect 210785 599044 210851 599045
rect 194542 598980 194548 599044
rect 194612 599042 194659 599044
rect 197118 599042 197124 599044
rect 194612 599040 194704 599042
rect 194654 598984 194704 599040
rect 194612 598982 194704 598984
rect 197078 598982 197124 599042
rect 197188 599040 197235 599044
rect 201534 599042 201540 599044
rect 197230 598984 197235 599040
rect 194612 598980 194659 598982
rect 197118 598980 197124 598982
rect 197188 598980 197235 598984
rect 201494 598982 201540 599042
rect 201604 599040 201651 599044
rect 203006 599042 203012 599044
rect 201646 598984 201651 599040
rect 201534 598980 201540 598982
rect 201604 598980 201651 598984
rect 202966 598982 203012 599042
rect 203076 599040 203123 599044
rect 207054 599042 207060 599044
rect 203118 598984 203123 599040
rect 203006 598980 203012 598982
rect 203076 598980 203123 598984
rect 207014 598982 207060 599042
rect 207124 599040 207171 599044
rect 210734 599042 210740 599044
rect 207166 598984 207171 599040
rect 207054 598980 207060 598982
rect 207124 598980 207171 598984
rect 210694 598982 210740 599042
rect 210804 599040 210851 599044
rect 210846 598984 210851 599040
rect 210734 598980 210740 598982
rect 210804 598980 210851 598984
rect 219566 598980 219572 599044
rect 219636 599042 219642 599044
rect 219709 599042 219775 599045
rect 220905 599044 220971 599045
rect 223849 599044 223915 599045
rect 220854 599042 220860 599044
rect 219636 599040 219775 599042
rect 219636 598984 219714 599040
rect 219770 598984 219775 599040
rect 219636 598982 219775 598984
rect 220814 598982 220860 599042
rect 220924 599040 220971 599044
rect 223798 599042 223804 599044
rect 220966 598984 220971 599040
rect 219636 598980 219642 598982
rect 194593 598979 194659 598980
rect 197169 598979 197235 598980
rect 201585 598979 201651 598980
rect 203057 598979 203123 598980
rect 207105 598979 207171 598980
rect 210785 598979 210851 598980
rect 219709 598979 219775 598982
rect 220854 598980 220860 598982
rect 220924 598980 220971 598984
rect 223758 598982 223804 599042
rect 223868 599040 223915 599044
rect 223910 598984 223915 599040
rect 223798 598980 223804 598982
rect 223868 598980 223915 598984
rect 223982 598980 223988 599044
rect 224052 599042 224058 599044
rect 224217 599042 224283 599045
rect 224052 599040 224283 599042
rect 224052 598984 224222 599040
rect 224278 598984 224283 599040
rect 224052 598982 224283 598984
rect 224052 598980 224058 598982
rect 220905 598979 220971 598980
rect 223849 598979 223915 598980
rect 224217 598979 224283 598982
rect 228214 598980 228220 599044
rect 228284 599042 228290 599044
rect 230013 599042 230079 599045
rect 230657 599044 230723 599045
rect 233233 599044 233299 599045
rect 234705 599044 234771 599045
rect 230606 599042 230612 599044
rect 228284 599040 230079 599042
rect 228284 598984 230018 599040
rect 230074 598984 230079 599040
rect 228284 598982 230079 598984
rect 230566 598982 230612 599042
rect 230676 599040 230723 599044
rect 233182 599042 233188 599044
rect 230718 598984 230723 599040
rect 228284 598980 228290 598982
rect 230013 598979 230079 598982
rect 230606 598980 230612 598982
rect 230676 598980 230723 598984
rect 233142 598982 233188 599042
rect 233252 599040 233299 599044
rect 234654 599042 234660 599044
rect 233294 598984 233299 599040
rect 233182 598980 233188 598982
rect 233252 598980 233299 598984
rect 234614 598982 234660 599042
rect 234724 599040 234771 599044
rect 234766 598984 234771 599040
rect 234654 598980 234660 598982
rect 234724 598980 234771 598984
rect 236494 598980 236500 599044
rect 236564 599042 236570 599044
rect 236821 599042 236887 599045
rect 236564 599040 236887 599042
rect 236564 598984 236826 599040
rect 236882 598984 236887 599040
rect 236564 598982 236887 598984
rect 236564 598980 236570 598982
rect 230657 598979 230723 598980
rect 233233 598979 233299 598980
rect 234705 598979 234771 598980
rect 236821 598979 236887 598982
rect 240685 599044 240751 599045
rect 240685 599040 240732 599044
rect 240796 599042 240802 599044
rect 242617 599042 242683 599045
rect 247769 599044 247835 599045
rect 242934 599042 242940 599044
rect 240685 598984 240690 599040
rect 240685 598980 240732 598984
rect 240796 598982 240842 599042
rect 242617 599040 242940 599042
rect 242617 598984 242622 599040
rect 242678 598984 242940 599040
rect 242617 598982 242940 598984
rect 240796 598980 240802 598982
rect 240685 598979 240751 598980
rect 242617 598979 242683 598982
rect 242934 598980 242940 598982
rect 243004 598980 243010 599044
rect 247718 599042 247724 599044
rect 247678 598982 247724 599042
rect 247788 599040 247835 599044
rect 247830 598984 247835 599040
rect 247718 598980 247724 598982
rect 247788 598980 247835 598984
rect 249926 598980 249932 599044
rect 249996 599042 250002 599044
rect 250253 599042 250319 599045
rect 249996 599040 250319 599042
rect 249996 598984 250258 599040
rect 250314 598984 250319 599040
rect 249996 598982 250319 598984
rect 249996 598980 250002 598982
rect 247769 598979 247835 598980
rect 250253 598979 250319 598982
rect 252502 598980 252508 599044
rect 252572 599042 252578 599044
rect 252829 599042 252895 599045
rect 252572 599040 252895 599042
rect 252572 598984 252834 599040
rect 252890 598984 252895 599040
rect 252572 598982 252895 598984
rect 252572 598980 252578 598982
rect 252829 598979 252895 598982
rect 255957 598906 256023 598909
rect 253430 598904 256023 598906
rect 253430 598848 255962 598904
rect 256018 598848 256023 598904
rect 253430 598846 256023 598848
rect 253430 598808 253490 598846
rect 255957 598843 256023 598846
rect 193254 598436 193260 598500
rect 193324 598498 193330 598500
rect 193489 598498 193555 598501
rect 193324 598496 193555 598498
rect 193324 598440 193494 598496
rect 193550 598440 193555 598496
rect 193324 598438 193555 598440
rect 193324 598436 193330 598438
rect 193489 598435 193555 598438
rect 133689 598226 133755 598229
rect 192334 598226 192340 598228
rect 133689 598224 192340 598226
rect 133689 598168 133694 598224
rect 133750 598168 192340 598224
rect 133689 598166 192340 598168
rect 133689 598163 133755 598166
rect 192334 598164 192340 598166
rect 192404 598164 192410 598228
rect 191005 597954 191071 597957
rect 193630 597954 193690 598264
rect 191005 597952 193690 597954
rect 191005 597896 191010 597952
rect 191066 597896 193690 597952
rect 191005 597894 193690 597896
rect 191005 597891 191071 597894
rect 253430 597682 253490 597720
rect 256601 597682 256667 597685
rect 253430 597680 256667 597682
rect 253430 597624 256606 597680
rect 256662 597624 256667 597680
rect 253430 597622 256667 597624
rect 256601 597619 256667 597622
rect 191649 597274 191715 597277
rect 191649 597272 193690 597274
rect 191649 597216 191654 597272
rect 191710 597216 193690 597272
rect 191649 597214 193690 597216
rect 191649 597211 191715 597214
rect 193630 597176 193690 597214
rect 188245 596866 188311 596869
rect 193438 596866 193444 596868
rect 188245 596864 193444 596866
rect 188245 596808 188250 596864
rect 188306 596808 193444 596864
rect 188245 596806 193444 596808
rect 188245 596803 188311 596806
rect 193438 596804 193444 596806
rect 193508 596804 193514 596868
rect 188245 596324 188311 596325
rect 188245 596320 188292 596324
rect 188356 596322 188362 596324
rect 191373 596322 191439 596325
rect 193630 596322 193690 596360
rect 188245 596264 188250 596320
rect 188245 596260 188292 596264
rect 188356 596262 188402 596322
rect 191373 596320 193690 596322
rect 191373 596264 191378 596320
rect 191434 596264 193690 596320
rect 191373 596262 193690 596264
rect 253430 596322 253490 596904
rect 270534 596322 270540 596324
rect 253430 596262 270540 596322
rect 188356 596260 188362 596262
rect 188245 596259 188311 596260
rect 191373 596259 191439 596262
rect 270534 596260 270540 596262
rect 270604 596260 270610 596324
rect 186221 595506 186287 595509
rect 193254 595506 193260 595508
rect 186221 595504 193260 595506
rect 186221 595448 186226 595504
rect 186282 595448 193260 595504
rect 186221 595446 193260 595448
rect 186221 595443 186287 595446
rect 193254 595444 193260 595446
rect 193324 595444 193330 595508
rect 191097 594962 191163 594965
rect 193630 594962 193690 595544
rect 253430 595234 253490 595816
rect 256601 595234 256667 595237
rect 253430 595232 256667 595234
rect 253430 595176 256606 595232
rect 256662 595176 256667 595232
rect 253430 595174 256667 595176
rect 256601 595171 256667 595174
rect 191097 594960 193690 594962
rect 191097 594904 191102 594960
rect 191158 594904 193690 594960
rect 191097 594902 193690 594904
rect 191097 594899 191163 594902
rect 253430 594826 253490 595000
rect 258390 594826 258396 594828
rect 253430 594766 258396 594826
rect 258390 594764 258396 594766
rect 258460 594764 258466 594828
rect 191281 594010 191347 594013
rect 193630 594010 193690 594456
rect 191281 594008 193690 594010
rect 191281 593952 191286 594008
rect 191342 593952 193690 594008
rect 191281 593950 193690 593952
rect 191281 593947 191347 593950
rect 253430 593874 253490 594184
rect 255405 593874 255471 593877
rect 253430 593872 255471 593874
rect 253430 593816 255410 593872
rect 255466 593816 255471 593872
rect 253430 593814 255471 593816
rect 255405 593811 255471 593814
rect 193029 593466 193095 593469
rect 193630 593466 193690 593640
rect 193029 593464 193690 593466
rect 193029 593408 193034 593464
rect 193090 593408 193690 593464
rect 193029 593406 193690 593408
rect 193029 593403 193095 593406
rect 142613 593330 142679 593333
rect 143441 593330 143507 593333
rect 191189 593330 191255 593333
rect 142613 593328 191255 593330
rect 142613 593272 142618 593328
rect 142674 593272 143446 593328
rect 143502 593272 191194 593328
rect 191250 593272 191255 593328
rect 142613 593270 191255 593272
rect 142613 593267 142679 593270
rect 143441 593267 143507 593270
rect 191189 593267 191255 593270
rect -960 592908 480 593148
rect 253430 593058 253490 593096
rect 255405 593058 255471 593061
rect 253430 593056 255471 593058
rect 253430 593000 255410 593056
rect 255466 593000 255471 593056
rect 253430 592998 255471 593000
rect 255405 592995 255471 592998
rect 254761 592650 254827 592653
rect 269062 592650 269068 592652
rect 254761 592648 269068 592650
rect 254761 592592 254766 592648
rect 254822 592592 269068 592648
rect 254761 592590 269068 592592
rect 254761 592587 254827 592590
rect 269062 592588 269068 592590
rect 269132 592588 269138 592652
rect 191373 592106 191439 592109
rect 193630 592106 193690 592552
rect 253933 592310 253999 592313
rect 253460 592308 253999 592310
rect 253460 592252 253938 592308
rect 253994 592252 253999 592308
rect 253460 592250 253999 592252
rect 253933 592247 253999 592250
rect 191373 592104 193690 592106
rect 191373 592048 191378 592104
rect 191434 592048 193690 592104
rect 191373 592046 193690 592048
rect 191373 592043 191439 592046
rect 191281 591290 191347 591293
rect 193630 591290 193690 591736
rect 191281 591288 193690 591290
rect 191281 591232 191286 591288
rect 191342 591232 193690 591288
rect 191281 591230 193690 591232
rect 191281 591227 191347 591230
rect 253430 590746 253490 591192
rect 582373 591018 582439 591021
rect 583520 591018 584960 591108
rect 582373 591016 584960 591018
rect 582373 590960 582378 591016
rect 582434 590960 584960 591016
rect 582373 590958 584960 590960
rect 582373 590955 582439 590958
rect 583520 590868 584960 590958
rect 267774 590746 267780 590748
rect 253430 590686 267780 590746
rect 267774 590684 267780 590686
rect 267844 590684 267850 590748
rect 193814 590204 193874 590648
rect 193806 590140 193812 590204
rect 193876 590140 193882 590204
rect 253430 589930 253490 590376
rect 255405 589930 255471 589933
rect 253430 589928 255471 589930
rect 253430 589872 255410 589928
rect 255466 589872 255471 589928
rect 253430 589870 255471 589872
rect 255405 589867 255471 589870
rect 255957 589930 256023 589933
rect 281574 589930 281580 589932
rect 255957 589928 281580 589930
rect 255957 589872 255962 589928
rect 256018 589872 281580 589928
rect 255957 589870 281580 589872
rect 255957 589867 256023 589870
rect 281574 589868 281580 589870
rect 281644 589868 281650 589932
rect 191373 589386 191439 589389
rect 193630 589386 193690 589832
rect 255497 589386 255563 589389
rect 191373 589384 193690 589386
rect 191373 589328 191378 589384
rect 191434 589328 193690 589384
rect 191373 589326 193690 589328
rect 253430 589384 255563 589386
rect 253430 589328 255502 589384
rect 255558 589328 255563 589384
rect 253430 589326 255563 589328
rect 191373 589323 191439 589326
rect 253430 589288 253490 589326
rect 255497 589323 255563 589326
rect 190545 588162 190611 588165
rect 193630 588162 193690 588744
rect 190545 588160 193690 588162
rect 190545 588104 190550 588160
rect 190606 588104 193690 588160
rect 190545 588102 193690 588104
rect 190545 588099 190611 588102
rect 159766 587964 159772 588028
rect 159836 588026 159842 588028
rect 253430 588026 253490 588472
rect 255957 588026 256023 588029
rect 159836 587966 193690 588026
rect 253430 588024 256023 588026
rect 253430 587968 255962 588024
rect 256018 587968 256023 588024
rect 253430 587966 256023 587968
rect 159836 587964 159842 587966
rect 193630 587928 193690 587966
rect 255957 587963 256023 587966
rect 190453 586530 190519 586533
rect 190453 586528 190562 586530
rect 190453 586472 190458 586528
rect 190514 586472 190562 586528
rect 190453 586467 190562 586472
rect 190502 586394 190562 586467
rect 193630 586394 193690 587112
rect 253430 586938 253490 587384
rect 255497 587210 255563 587213
rect 265750 587210 265756 587212
rect 255497 587208 265756 587210
rect 255497 587152 255502 587208
rect 255558 587152 265756 587208
rect 255497 587150 265756 587152
rect 255497 587147 255563 587150
rect 265750 587148 265756 587150
rect 265820 587148 265826 587212
rect 254025 586938 254091 586941
rect 253430 586936 254091 586938
rect 253430 586880 254030 586936
rect 254086 586880 254091 586936
rect 253430 586878 254091 586880
rect 254025 586875 254091 586878
rect 190502 586334 193690 586394
rect 253430 586394 253490 586568
rect 266302 586468 266308 586532
rect 266372 586468 266378 586532
rect 266310 586394 266370 586468
rect 253430 586334 266370 586394
rect 191741 586122 191807 586125
rect 191741 586120 193690 586122
rect 191741 586064 191746 586120
rect 191802 586064 193690 586120
rect 191741 586062 193690 586064
rect 191741 586059 191807 586062
rect 193630 586024 193690 586062
rect 191005 585170 191071 585173
rect 193630 585170 193690 585208
rect 191005 585168 193690 585170
rect 191005 585112 191010 585168
rect 191066 585112 193690 585168
rect 191005 585110 193690 585112
rect 253430 585170 253490 585480
rect 255313 585170 255379 585173
rect 253430 585168 255379 585170
rect 253430 585112 255318 585168
rect 255374 585112 255379 585168
rect 253430 585110 255379 585112
rect 191005 585107 191071 585110
rect 255313 585107 255379 585110
rect 253430 584354 253490 584664
rect 255497 584354 255563 584357
rect 253430 584352 255563 584354
rect 253430 584296 255502 584352
rect 255558 584296 255563 584352
rect 253430 584294 255563 584296
rect 255497 584291 255563 584294
rect 255405 584218 255471 584221
rect 253430 584216 255471 584218
rect 253430 584160 255410 584216
rect 255466 584160 255471 584216
rect 253430 584158 255471 584160
rect 191741 583946 191807 583949
rect 193630 583946 193690 584120
rect 191741 583944 193690 583946
rect 191741 583888 191746 583944
rect 191802 583888 193690 583944
rect 191741 583886 193690 583888
rect 191741 583883 191807 583886
rect 253430 583848 253490 584158
rect 255405 584155 255471 584158
rect 94865 583402 94931 583405
rect 98637 583402 98703 583405
rect 94865 583400 98703 583402
rect 94865 583344 94870 583400
rect 94926 583344 98642 583400
rect 98698 583344 98703 583400
rect 94865 583342 98703 583344
rect 94865 583339 94931 583342
rect 98637 583339 98703 583342
rect 82721 582722 82787 582725
rect 119337 582722 119403 582725
rect 82721 582720 119403 582722
rect 82721 582664 82726 582720
rect 82782 582664 119342 582720
rect 119398 582664 119403 582720
rect 82721 582662 119403 582664
rect 82721 582659 82787 582662
rect 119337 582659 119403 582662
rect 191281 582722 191347 582725
rect 193630 582722 193690 583304
rect 191281 582720 193690 582722
rect 191281 582664 191286 582720
rect 191342 582664 193690 582720
rect 191281 582662 193690 582664
rect 191281 582659 191347 582662
rect 73521 582586 73587 582589
rect 95877 582586 95943 582589
rect 73521 582584 95943 582586
rect 73521 582528 73526 582584
rect 73582 582528 95882 582584
rect 95938 582528 95943 582584
rect 73521 582526 95943 582528
rect 253430 582586 253490 582760
rect 255405 582586 255471 582589
rect 253430 582584 255471 582586
rect 253430 582528 255410 582584
rect 255466 582528 255471 582584
rect 253430 582526 255471 582528
rect 73521 582523 73587 582526
rect 95877 582523 95943 582526
rect 255405 582523 255471 582526
rect 254117 582314 254183 582317
rect 253430 582312 254183 582314
rect 253430 582256 254122 582312
rect 254178 582256 254183 582312
rect 253430 582254 254183 582256
rect 191189 581770 191255 581773
rect 193630 581770 193690 582216
rect 253430 581944 253490 582254
rect 254117 582251 254183 582254
rect 191189 581768 193690 581770
rect 191189 581712 191194 581768
rect 191250 581712 193690 581768
rect 191189 581710 193690 581712
rect 191189 581707 191255 581710
rect 93761 581226 93827 581229
rect 106917 581226 106983 581229
rect 93761 581224 106983 581226
rect 93761 581168 93766 581224
rect 93822 581168 106922 581224
rect 106978 581168 106983 581224
rect 93761 581166 106983 581168
rect 93761 581163 93827 581166
rect 106917 581163 106983 581166
rect 191741 581226 191807 581229
rect 193630 581226 193690 581400
rect 191741 581224 193690 581226
rect 191741 581168 191746 581224
rect 191802 581168 193690 581224
rect 191741 581166 193690 581168
rect 191741 581163 191807 581166
rect 67449 581090 67515 581093
rect 160829 581090 160895 581093
rect 67449 581088 160895 581090
rect 67449 581032 67454 581088
rect 67510 581032 160834 581088
rect 160890 581032 160895 581088
rect 67449 581030 160895 581032
rect 67449 581027 67515 581030
rect 160829 581027 160895 581030
rect 75361 580954 75427 580957
rect 75678 580954 75684 580956
rect 75361 580952 75684 580954
rect 75361 580896 75366 580952
rect 75422 580896 75684 580952
rect 75361 580894 75684 580896
rect 75361 580891 75427 580894
rect 75678 580892 75684 580894
rect 75748 580892 75754 580956
rect 70945 580820 71011 580821
rect 79961 580820 80027 580821
rect 70894 580818 70900 580820
rect 70854 580758 70900 580818
rect 70964 580816 71011 580820
rect 79910 580818 79916 580820
rect 71006 580760 71011 580816
rect 70894 580756 70900 580758
rect 70964 580756 71011 580760
rect 79870 580758 79916 580818
rect 79980 580816 80027 580820
rect 80022 580760 80027 580816
rect 79910 580756 79916 580758
rect 79980 580756 80027 580760
rect 70945 580755 71011 580756
rect 79961 580755 80027 580756
rect 84653 580820 84719 580821
rect 89253 580820 89319 580821
rect 84653 580816 84700 580820
rect 84764 580818 84770 580820
rect 84653 580760 84658 580816
rect 84653 580756 84700 580760
rect 84764 580758 84810 580818
rect 89253 580816 89300 580820
rect 89364 580818 89370 580820
rect 89253 580760 89258 580816
rect 84764 580756 84770 580758
rect 89253 580756 89300 580760
rect 89364 580758 89410 580818
rect 89364 580756 89370 580758
rect 84653 580755 84719 580756
rect 89253 580755 89319 580756
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 66897 580002 66963 580005
rect 68878 580002 68938 580584
rect 66897 580000 68938 580002
rect 66897 579944 66902 580000
rect 66958 579944 68938 580000
rect 66897 579942 68938 579944
rect 66897 579939 66963 579942
rect 191557 579730 191623 579733
rect 193630 579730 193690 580312
rect 253430 580274 253490 580856
rect 255497 580274 255563 580277
rect 253430 580272 255563 580274
rect 253430 580216 255502 580272
rect 255558 580216 255563 580272
rect 253430 580214 255563 580216
rect 255497 580211 255563 580214
rect 253430 579866 253490 580040
rect 255405 579866 255471 579869
rect 253430 579864 255471 579866
rect 253430 579808 255410 579864
rect 255466 579808 255471 579864
rect 253430 579806 255471 579808
rect 255405 579803 255471 579806
rect 191557 579728 193690 579730
rect 191557 579672 191562 579728
rect 191618 579672 193690 579728
rect 191557 579670 193690 579672
rect 191557 579667 191623 579670
rect 66662 578580 66668 578644
rect 66732 578642 66738 578644
rect 68878 578642 68938 579224
rect 94638 578914 94698 579496
rect 190913 579050 190979 579053
rect 193630 579050 193690 579496
rect 190913 579048 193690 579050
rect 190913 578992 190918 579048
rect 190974 578992 193690 579048
rect 190913 578990 193690 578992
rect 190913 578987 190979 578990
rect 96889 578914 96955 578917
rect 94638 578912 96955 578914
rect 94638 578856 96894 578912
rect 96950 578856 96955 578912
rect 94638 578854 96955 578856
rect 96889 578851 96955 578854
rect 156638 578852 156644 578916
rect 156708 578914 156714 578916
rect 191557 578914 191623 578917
rect 156708 578912 191623 578914
rect 156708 578856 191562 578912
rect 191618 578856 191623 578912
rect 156708 578854 191623 578856
rect 156708 578852 156714 578854
rect 191557 578851 191623 578854
rect 66732 578582 68938 578642
rect 253430 578642 253490 578952
rect 255313 578642 255379 578645
rect 253430 578640 255379 578642
rect 253430 578584 255318 578640
rect 255374 578584 255379 578640
rect 253430 578582 255379 578584
rect 66732 578580 66738 578582
rect 255313 578579 255379 578582
rect 191649 578370 191715 578373
rect 193630 578370 193690 578408
rect 191649 578368 193690 578370
rect 191649 578312 191654 578368
rect 191710 578312 193690 578368
rect 191649 578310 193690 578312
rect 191649 578307 191715 578310
rect 67541 577282 67607 577285
rect 68878 577282 68938 577864
rect 94638 577554 94698 578136
rect 191741 578098 191807 578101
rect 191741 578096 193690 578098
rect 191741 578040 191746 578096
rect 191802 578040 193690 578096
rect 191741 578038 193690 578040
rect 191741 578035 191807 578038
rect 193630 577592 193690 578038
rect 253430 577690 253490 578136
rect 255405 577690 255471 577693
rect 253430 577688 255471 577690
rect 253430 577632 255410 577688
rect 255466 577632 255471 577688
rect 253430 577630 255471 577632
rect 255405 577627 255471 577630
rect 582373 577690 582439 577693
rect 583520 577690 584960 577780
rect 582373 577688 584960 577690
rect 582373 577632 582378 577688
rect 582434 577632 584960 577688
rect 582373 577630 584960 577632
rect 582373 577627 582439 577630
rect 97901 577554 97967 577557
rect 94638 577552 97967 577554
rect 94638 577496 97906 577552
rect 97962 577496 97967 577552
rect 583520 577540 584960 577630
rect 94638 577494 97967 577496
rect 97901 577491 97967 577494
rect 67541 577280 68938 577282
rect 67541 577224 67546 577280
rect 67602 577224 68938 577280
rect 67541 577222 68938 577224
rect 67541 577219 67607 577222
rect 253430 577010 253490 577048
rect 255405 577010 255471 577013
rect 253430 577008 255471 577010
rect 253430 576952 255410 577008
rect 255466 576952 255471 577008
rect 253430 576950 255471 576952
rect 255405 576947 255471 576950
rect 94638 576738 94698 576776
rect 97901 576738 97967 576741
rect 94638 576736 97967 576738
rect 94638 576680 97906 576736
rect 97962 576680 97967 576736
rect 94638 576678 97967 576680
rect 97901 576675 97967 576678
rect 66161 575922 66227 575925
rect 67725 575922 67791 575925
rect 68878 575922 68938 576504
rect 191649 576194 191715 576197
rect 193630 576194 193690 576776
rect 191649 576192 193690 576194
rect 191649 576136 191654 576192
rect 191710 576136 193690 576192
rect 191649 576134 193690 576136
rect 191649 576131 191715 576134
rect 66161 575920 68938 575922
rect 66161 575864 66166 575920
rect 66222 575864 67730 575920
rect 67786 575864 68938 575920
rect 66161 575862 68938 575864
rect 253430 575922 253490 576232
rect 255405 575922 255471 575925
rect 253430 575920 255471 575922
rect 253430 575864 255410 575920
rect 255466 575864 255471 575920
rect 253430 575862 255471 575864
rect 66161 575859 66227 575862
rect 67725 575859 67791 575862
rect 255405 575859 255471 575862
rect 191741 575650 191807 575653
rect 193630 575650 193690 575688
rect 191741 575648 193690 575650
rect 191741 575592 191746 575648
rect 191802 575592 193690 575648
rect 191741 575590 193690 575592
rect 191741 575587 191807 575590
rect 67357 575106 67423 575109
rect 68878 575106 68938 575144
rect 67357 575104 68938 575106
rect 67357 575048 67362 575104
rect 67418 575048 68938 575104
rect 67357 575046 68938 575048
rect 94638 575106 94698 575416
rect 97901 575106 97967 575109
rect 94638 575104 97967 575106
rect 94638 575048 97906 575104
rect 97962 575048 97967 575104
rect 94638 575046 97967 575048
rect 67357 575043 67423 575046
rect 97901 575043 97967 575046
rect 190821 574562 190887 574565
rect 193630 574562 193690 574872
rect 253430 574698 253490 575144
rect 255405 574698 255471 574701
rect 253430 574696 255471 574698
rect 253430 574640 255410 574696
rect 255466 574640 255471 574696
rect 253430 574638 255471 574640
rect 255405 574635 255471 574638
rect 190821 574560 193690 574562
rect 190821 574504 190826 574560
rect 190882 574504 193690 574560
rect 190821 574502 193690 574504
rect 190821 574499 190887 574502
rect 253430 574154 253490 574328
rect 255589 574154 255655 574157
rect 253430 574152 255655 574154
rect 253430 574096 255594 574152
rect 255650 574096 255655 574152
rect 253430 574094 255655 574096
rect 255589 574091 255655 574094
rect 66805 573202 66871 573205
rect 68878 573202 68938 573784
rect 94638 573474 94698 574056
rect 97533 573474 97599 573477
rect 94638 573472 97599 573474
rect 94638 573416 97538 573472
rect 97594 573416 97599 573472
rect 94638 573414 97599 573416
rect 97533 573411 97599 573414
rect 193630 573202 193690 573784
rect 66805 573200 68938 573202
rect 66805 573144 66810 573200
rect 66866 573144 68938 573200
rect 66805 573142 68938 573144
rect 180750 573142 193690 573202
rect 66805 573139 66871 573142
rect 178534 572732 178540 572796
rect 178604 572794 178610 572796
rect 180750 572794 180810 573142
rect 178604 572734 180810 572794
rect 191741 572794 191807 572797
rect 193630 572794 193690 572968
rect 253430 572930 253490 573512
rect 255681 572930 255747 572933
rect 253430 572928 255747 572930
rect 253430 572872 255686 572928
rect 255742 572872 255747 572928
rect 253430 572870 255747 572872
rect 255681 572867 255747 572870
rect 191741 572792 193690 572794
rect 191741 572736 191746 572792
rect 191802 572736 193690 572792
rect 191741 572734 193690 572736
rect 178604 572732 178610 572734
rect 191741 572731 191807 572734
rect 67449 572658 67515 572661
rect 94638 572658 94698 572696
rect 97257 572658 97323 572661
rect 67449 572656 68938 572658
rect 67449 572600 67454 572656
rect 67510 572600 68938 572656
rect 67449 572598 68938 572600
rect 94638 572656 97323 572658
rect 94638 572600 97262 572656
rect 97318 572600 97323 572656
rect 94638 572598 97323 572600
rect 67449 572595 67515 572598
rect 68878 572424 68938 572598
rect 97257 572595 97323 572598
rect 190821 572250 190887 572253
rect 190821 572248 193690 572250
rect 190821 572192 190826 572248
rect 190882 572192 193690 572248
rect 190821 572190 193690 572192
rect 190821 572187 190887 572190
rect 193630 571880 193690 572190
rect 253430 571978 253490 572424
rect 255497 571978 255563 571981
rect 253430 571976 255563 571978
rect 253430 571920 255502 571976
rect 255558 571920 255563 571976
rect 253430 571918 255563 571920
rect 255497 571915 255563 571918
rect 253430 571570 253490 571608
rect 255405 571570 255471 571573
rect 253430 571568 255471 571570
rect 253430 571512 255410 571568
rect 255466 571512 255471 571568
rect 253430 571510 255471 571512
rect 255405 571507 255471 571510
rect 97717 571434 97783 571437
rect 94638 571432 97783 571434
rect 94638 571376 97722 571432
rect 97778 571376 97783 571432
rect 94638 571374 97783 571376
rect 94638 571336 94698 571374
rect 97717 571371 97783 571374
rect 191741 570890 191807 570893
rect 193630 570890 193690 571064
rect 191741 570888 193690 570890
rect 191741 570832 191746 570888
rect 191802 570832 193690 570888
rect 191741 570830 193690 570832
rect 191741 570827 191807 570830
rect 67449 570210 67515 570213
rect 68878 570210 68938 570792
rect 255262 570618 255268 570620
rect 253430 570558 255268 570618
rect 253430 570520 253490 570558
rect 255262 570556 255268 570558
rect 255332 570618 255338 570620
rect 255405 570618 255471 570621
rect 255332 570616 255471 570618
rect 255332 570560 255410 570616
rect 255466 570560 255471 570616
rect 255332 570558 255471 570560
rect 255332 570556 255338 570558
rect 255405 570555 255471 570558
rect 67449 570208 68938 570210
rect 67449 570152 67454 570208
rect 67510 570152 68938 570208
rect 67449 570150 68938 570152
rect 67449 570147 67515 570150
rect 97901 570074 97967 570077
rect 94638 570072 97967 570074
rect 94638 570016 97906 570072
rect 97962 570016 97967 570072
rect 94638 570014 97967 570016
rect 94638 569976 94698 570014
rect 97901 570011 97967 570014
rect 191741 570074 191807 570077
rect 191741 570072 193690 570074
rect 191741 570016 191746 570072
rect 191802 570016 193690 570072
rect 191741 570014 193690 570016
rect 191741 570011 191807 570014
rect 193630 569976 193690 570014
rect 65977 569938 66043 569941
rect 65977 569936 68938 569938
rect 65977 569880 65982 569936
rect 66038 569880 68938 569936
rect 65977 569878 68938 569880
rect 65977 569875 66043 569878
rect 68878 569432 68938 569878
rect 253430 569258 253490 569704
rect 255497 569258 255563 569261
rect 253430 569256 255563 569258
rect 253430 569200 255502 569256
rect 255558 569200 255563 569256
rect 253430 569198 255563 569200
rect 255497 569195 255563 569198
rect 96705 569122 96771 569125
rect 97901 569122 97967 569125
rect 94638 569120 97967 569122
rect 94638 569064 96710 569120
rect 96766 569064 97906 569120
rect 97962 569064 97967 569120
rect 94638 569062 97967 569064
rect 94638 568616 94698 569062
rect 96705 569059 96771 569062
rect 97901 569059 97967 569062
rect 172094 568652 172100 568716
rect 172164 568714 172170 568716
rect 193630 568714 193690 569160
rect 255405 568714 255471 568717
rect 172164 568654 193690 568714
rect 253430 568712 255471 568714
rect 253430 568656 255410 568712
rect 255466 568656 255471 568712
rect 253430 568654 255471 568656
rect 172164 568652 172170 568654
rect 253430 568616 253490 568654
rect 255405 568651 255471 568654
rect 66897 567490 66963 567493
rect 68878 567490 68938 568072
rect 164969 567898 165035 567901
rect 191097 567898 191163 567901
rect 164969 567896 191163 567898
rect 164969 567840 164974 567896
rect 165030 567840 191102 567896
rect 191158 567840 191163 567896
rect 164969 567838 191163 567840
rect 164969 567835 165035 567838
rect 191097 567835 191163 567838
rect 66897 567488 68938 567490
rect 66897 567432 66902 567488
rect 66958 567432 68938 567488
rect 66897 567430 68938 567432
rect 189717 567490 189783 567493
rect 193630 567490 193690 568072
rect 189717 567488 193690 567490
rect 189717 567432 189722 567488
rect 189778 567432 193690 567488
rect 189717 567430 193690 567432
rect 253430 567490 253490 567800
rect 256877 567490 256943 567493
rect 253430 567488 256943 567490
rect 253430 567432 256882 567488
rect 256938 567432 256943 567488
rect 253430 567430 256943 567432
rect 66897 567427 66963 567430
rect 189717 567427 189783 567430
rect 256877 567427 256943 567430
rect 94638 567218 94698 567256
rect 97901 567218 97967 567221
rect 94638 567216 97967 567218
rect 94638 567160 97906 567216
rect 97962 567160 97967 567216
rect 94638 567158 97967 567160
rect 97901 567155 97967 567158
rect 191373 567218 191439 567221
rect 193630 567218 193690 567256
rect 191373 567216 193690 567218
rect 191373 567160 191378 567216
rect 191434 567160 193690 567216
rect 191373 567158 193690 567160
rect 191373 567155 191439 567158
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67633 566674 67699 566677
rect 68878 566674 68938 566712
rect 67633 566672 68938 566674
rect 67633 566616 67638 566672
rect 67694 566616 68938 566672
rect 67633 566614 68938 566616
rect 67633 566611 67699 566614
rect 94638 565858 94698 565896
rect 95417 565858 95483 565861
rect 94638 565856 95483 565858
rect 94638 565800 95422 565856
rect 95478 565800 95483 565856
rect 94638 565798 95483 565800
rect 95417 565795 95483 565798
rect 166758 565796 166764 565860
rect 166828 565858 166834 565860
rect 193630 565858 193690 566440
rect 253430 566266 253490 566712
rect 255589 566266 255655 566269
rect 253430 566264 255655 566266
rect 253430 566208 255594 566264
rect 255650 566208 255655 566264
rect 253430 566206 255655 566208
rect 255589 566203 255655 566206
rect 255497 565994 255563 565997
rect 253430 565992 255563 565994
rect 253430 565936 255502 565992
rect 255558 565936 255563 565992
rect 253430 565934 255563 565936
rect 253430 565896 253490 565934
rect 255497 565931 255563 565934
rect 166828 565798 193690 565858
rect 166828 565796 166834 565798
rect 66437 564906 66503 564909
rect 68878 564906 68938 565352
rect 191281 565178 191347 565181
rect 193630 565178 193690 565352
rect 191281 565176 193690 565178
rect 191281 565120 191286 565176
rect 191342 565120 193690 565176
rect 191281 565118 193690 565120
rect 191281 565115 191347 565118
rect 191741 565042 191807 565045
rect 191741 565040 193690 565042
rect 191741 564984 191746 565040
rect 191802 564984 193690 565040
rect 191741 564982 193690 564984
rect 191741 564979 191807 564982
rect 66437 564904 68938 564906
rect 66437 564848 66442 564904
rect 66498 564848 68938 564904
rect 66437 564846 68938 564848
rect 66437 564843 66503 564846
rect 193630 564536 193690 564982
rect 253430 564770 253490 565080
rect 255497 564770 255563 564773
rect 253430 564768 255563 564770
rect 253430 564712 255502 564768
rect 255558 564712 255563 564768
rect 253430 564710 255563 564712
rect 255497 564707 255563 564710
rect 582833 564362 582899 564365
rect 583520 564362 584960 564452
rect 582833 564360 584960 564362
rect 582833 564304 582838 564360
rect 582894 564304 584960 564360
rect 582833 564302 584960 564304
rect 582833 564299 582899 564302
rect 65885 563410 65951 563413
rect 68878 563410 68938 563992
rect 94638 563682 94698 564264
rect 583520 564212 584960 564302
rect 95233 563682 95299 563685
rect 94638 563680 95299 563682
rect 94638 563624 95238 563680
rect 95294 563624 95299 563680
rect 94638 563622 95299 563624
rect 95233 563619 95299 563622
rect 191741 563682 191807 563685
rect 191741 563680 193690 563682
rect 191741 563624 191746 563680
rect 191802 563624 193690 563680
rect 191741 563622 193690 563624
rect 191741 563619 191807 563622
rect 193630 563448 193690 563622
rect 65885 563408 68938 563410
rect 65885 563352 65890 563408
rect 65946 563352 68938 563408
rect 65885 563350 68938 563352
rect 253430 563410 253490 563992
rect 260966 563410 260972 563412
rect 253430 563350 260972 563410
rect 65885 563347 65951 563350
rect 260966 563348 260972 563350
rect 261036 563348 261042 563412
rect 253430 563138 253490 563176
rect 263726 563138 263732 563140
rect 253430 563078 263732 563138
rect 263726 563076 263732 563078
rect 263796 563076 263802 563140
rect 67766 561988 67772 562052
rect 67836 562050 67842 562052
rect 68878 562050 68938 562632
rect 94638 562594 94698 562904
rect 97901 562594 97967 562597
rect 94638 562592 97967 562594
rect 94638 562536 97906 562592
rect 97962 562536 97967 562592
rect 94638 562534 97967 562536
rect 97901 562531 97967 562534
rect 190913 562186 190979 562189
rect 193630 562186 193690 562632
rect 190913 562184 193690 562186
rect 190913 562128 190918 562184
rect 190974 562128 193690 562184
rect 190913 562126 193690 562128
rect 190913 562123 190979 562126
rect 67836 561990 68938 562050
rect 67836 561988 67842 561990
rect 253430 561778 253490 562088
rect 255681 561778 255747 561781
rect 253430 561776 255747 561778
rect 253430 561720 255686 561776
rect 255742 561720 255747 561776
rect 253430 561718 255747 561720
rect 255681 561715 255747 561718
rect 66805 560690 66871 560693
rect 68878 560690 68938 561272
rect 94638 561098 94698 561544
rect 96797 561098 96863 561101
rect 97901 561098 97967 561101
rect 94638 561096 97967 561098
rect 94638 561040 96802 561096
rect 96858 561040 97906 561096
rect 97962 561040 97967 561096
rect 94638 561038 97967 561040
rect 96797 561035 96863 561038
rect 97901 561035 97967 561038
rect 190821 560962 190887 560965
rect 193630 560962 193690 561544
rect 190821 560960 193690 560962
rect 190821 560904 190826 560960
rect 190882 560904 193690 560960
rect 190821 560902 193690 560904
rect 190821 560899 190887 560902
rect 253430 560826 253490 561272
rect 255497 560826 255563 560829
rect 253430 560824 255563 560826
rect 253430 560768 255502 560824
rect 255558 560768 255563 560824
rect 253430 560766 255563 560768
rect 255497 560763 255563 560766
rect 66805 560688 68938 560690
rect 66805 560632 66810 560688
rect 66866 560632 68938 560688
rect 66805 560630 68938 560632
rect 66805 560627 66871 560630
rect 170806 560356 170812 560420
rect 170876 560418 170882 560420
rect 193630 560418 193690 560728
rect 170876 560358 193690 560418
rect 170876 560356 170882 560358
rect 66805 559330 66871 559333
rect 68878 559330 68938 559912
rect 94638 559602 94698 560184
rect 96889 559602 96955 559605
rect 94638 559600 96955 559602
rect 94638 559544 96894 559600
rect 96950 559544 96955 559600
rect 94638 559542 96955 559544
rect 96889 559539 96955 559542
rect 66805 559328 68938 559330
rect 66805 559272 66810 559328
rect 66866 559272 68938 559328
rect 66805 559270 68938 559272
rect 66805 559267 66871 559270
rect 191741 559194 191807 559197
rect 193630 559194 193690 559640
rect 253430 559602 253490 560184
rect 255589 559602 255655 559605
rect 253430 559600 255655 559602
rect 253430 559544 255594 559600
rect 255650 559544 255655 559600
rect 253430 559542 255655 559544
rect 255589 559539 255655 559542
rect 191741 559192 193690 559194
rect 191741 559136 191746 559192
rect 191802 559136 193690 559192
rect 191741 559134 193690 559136
rect 253430 559194 253490 559368
rect 255497 559194 255563 559197
rect 253430 559192 255563 559194
rect 253430 559136 255502 559192
rect 255558 559136 255563 559192
rect 253430 559134 255563 559136
rect 191741 559131 191807 559134
rect 255497 559131 255563 559134
rect 95141 558854 95207 558857
rect 94668 558852 95207 558854
rect 94668 558824 95146 558852
rect 94638 558796 95146 558824
rect 95202 558796 95207 558852
rect 94638 558794 95207 558796
rect 94638 558653 94698 558794
rect 95141 558791 95207 558794
rect 94638 558648 94747 558653
rect 94638 558592 94686 558648
rect 94742 558592 94747 558648
rect 94638 558590 94747 558592
rect 94681 558587 94747 558590
rect 66805 557970 66871 557973
rect 68878 557970 68938 558552
rect 186814 558180 186820 558244
rect 186884 558242 186890 558244
rect 193630 558242 193690 558824
rect 186884 558182 193690 558242
rect 186884 558180 186890 558182
rect 66805 557968 68938 557970
rect 66805 557912 66810 557968
rect 66866 557912 68938 557968
rect 66805 557910 68938 557912
rect 66805 557907 66871 557910
rect 191741 557834 191807 557837
rect 193630 557834 193690 558008
rect 253430 557970 253490 558280
rect 255589 557970 255655 557973
rect 253430 557968 255655 557970
rect 253430 557912 255594 557968
rect 255650 557912 255655 557968
rect 253430 557910 255655 557912
rect 255589 557907 255655 557910
rect 191741 557832 193690 557834
rect 191741 557776 191746 557832
rect 191802 557776 193690 557832
rect 191741 557774 193690 557776
rect 191741 557771 191807 557774
rect 67633 556610 67699 556613
rect 68878 556610 68938 557192
rect 94638 556882 94698 557464
rect 96705 556882 96771 556885
rect 97901 556882 97967 556885
rect 94638 556880 97967 556882
rect 94638 556824 96710 556880
rect 96766 556824 97906 556880
rect 97962 556824 97967 556880
rect 94638 556822 97967 556824
rect 96705 556819 96771 556822
rect 97901 556819 97967 556822
rect 67633 556608 68938 556610
rect 67633 556552 67638 556608
rect 67694 556552 68938 556608
rect 67633 556550 68938 556552
rect 67633 556547 67699 556550
rect 191741 556474 191807 556477
rect 193630 556474 193690 556920
rect 253430 556882 253490 557464
rect 255589 556882 255655 556885
rect 253430 556880 255655 556882
rect 253430 556824 255594 556880
rect 255650 556824 255655 556880
rect 253430 556822 255655 556824
rect 255589 556819 255655 556822
rect 191741 556472 193690 556474
rect 191741 556416 191746 556472
rect 191802 556416 193690 556472
rect 191741 556414 193690 556416
rect 191741 556411 191807 556414
rect 253430 556205 253490 556376
rect 253381 556200 253490 556205
rect 253381 556144 253386 556200
rect 253442 556144 253490 556200
rect 253381 556142 253490 556144
rect 253381 556139 253447 556142
rect 66529 555250 66595 555253
rect 68878 555250 68938 555832
rect 94638 555522 94698 556104
rect 95325 555522 95391 555525
rect 94638 555520 95391 555522
rect 94638 555464 95330 555520
rect 95386 555464 95391 555520
rect 94638 555462 95391 555464
rect 95325 555459 95391 555462
rect 193630 555250 193690 556104
rect 66529 555248 68938 555250
rect 66529 555192 66534 555248
rect 66590 555192 68938 555248
rect 66529 555190 68938 555192
rect 180750 555190 193690 555250
rect 66529 555187 66595 555190
rect 148174 554780 148180 554844
rect 148244 554842 148250 554844
rect 180750 554842 180810 555190
rect 191465 554978 191531 554981
rect 193630 554978 193690 555016
rect 191465 554976 193690 554978
rect 191465 554920 191470 554976
rect 191526 554920 193690 554976
rect 191465 554918 193690 554920
rect 253430 554978 253490 555560
rect 254117 554978 254183 554981
rect 253430 554976 254183 554978
rect 253430 554920 254122 554976
rect 254178 554920 254183 554976
rect 253430 554918 254183 554920
rect 191465 554915 191531 554918
rect 254117 554915 254183 554918
rect 148244 554782 180810 554842
rect 148244 554780 148250 554782
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 66897 553618 66963 553621
rect 68878 553618 68938 554200
rect 94638 554162 94698 554744
rect 96981 554162 97047 554165
rect 94638 554160 97047 554162
rect 94638 554104 96986 554160
rect 97042 554104 97047 554160
rect 94638 554102 97047 554104
rect 96981 554099 97047 554102
rect 116117 554026 116183 554029
rect 173157 554026 173223 554029
rect 66897 553616 68938 553618
rect 66897 553560 66902 553616
rect 66958 553560 68938 553616
rect 66897 553558 68938 553560
rect 103470 554024 173223 554026
rect 103470 553968 116122 554024
rect 116178 553968 173162 554024
rect 173218 553968 173223 554024
rect 103470 553966 173223 553968
rect 66897 553555 66963 553558
rect 96654 553420 96660 553484
rect 96724 553482 96730 553484
rect 103470 553482 103530 553966
rect 116117 553963 116183 553966
rect 173157 553963 173223 553966
rect 96724 553422 103530 553482
rect 189809 553482 189875 553485
rect 193630 553482 193690 554200
rect 253430 554162 253490 554744
rect 255681 554162 255747 554165
rect 253430 554160 255747 554162
rect 253430 554104 255686 554160
rect 255742 554104 255747 554160
rect 253430 554102 255747 554104
rect 255681 554099 255747 554102
rect 253430 553618 253490 553656
rect 255589 553618 255655 553621
rect 253430 553616 255655 553618
rect 253430 553560 255594 553616
rect 255650 553560 255655 553616
rect 253430 553558 255655 553560
rect 255589 553555 255655 553558
rect 189809 553480 193690 553482
rect 189809 553424 189814 553480
rect 189870 553424 193690 553480
rect 189809 553422 193690 553424
rect 96724 553420 96730 553422
rect 189809 553419 189875 553422
rect 67817 552258 67883 552261
rect 68878 552258 68938 552840
rect 94638 552802 94698 553384
rect 97901 552802 97967 552805
rect 94638 552800 97967 552802
rect 94638 552744 97906 552800
rect 97962 552744 97967 552800
rect 94638 552742 97967 552744
rect 97901 552739 97967 552742
rect 191097 552666 191163 552669
rect 193630 552666 193690 553112
rect 253430 552802 253490 552840
rect 255589 552802 255655 552805
rect 253430 552800 255655 552802
rect 253430 552744 255594 552800
rect 255650 552744 255655 552800
rect 253430 552742 255655 552744
rect 255589 552739 255655 552742
rect 191097 552664 193690 552666
rect 191097 552608 191102 552664
rect 191158 552608 193690 552664
rect 191097 552606 193690 552608
rect 191097 552603 191163 552606
rect 67817 552256 68938 552258
rect 67817 552200 67822 552256
rect 67878 552200 68938 552256
rect 67817 552198 68938 552200
rect 67817 552195 67883 552198
rect 158478 552196 158484 552260
rect 158548 552258 158554 552260
rect 193630 552258 193690 552296
rect 158548 552198 193690 552258
rect 158548 552196 158554 552198
rect 96613 552122 96679 552125
rect 97809 552122 97875 552125
rect 94638 552120 97875 552122
rect 94638 552064 96618 552120
rect 96674 552064 97814 552120
rect 97870 552064 97875 552120
rect 94638 552062 97875 552064
rect 94638 552024 94698 552062
rect 96613 552059 96679 552062
rect 97809 552059 97875 552062
rect 101397 551986 101463 551989
rect 104934 551986 104940 551988
rect 101397 551984 104940 551986
rect 101397 551928 101402 551984
rect 101458 551928 104940 551984
rect 101397 551926 104940 551928
rect 101397 551923 101463 551926
rect 104934 551924 104940 551926
rect 105004 551924 105010 551988
rect 253974 551782 253980 551784
rect 253460 551722 253980 551782
rect 253974 551720 253980 551722
rect 254044 551720 254050 551784
rect 69430 551172 69490 551480
rect 96654 551306 96660 551308
rect 94638 551246 96660 551306
rect 69422 551108 69428 551172
rect 69492 551108 69498 551172
rect 94638 550664 94698 551246
rect 96654 551244 96660 551246
rect 96724 551244 96730 551308
rect 191741 550762 191807 550765
rect 193630 550762 193690 551208
rect 583520 551020 584960 551260
rect 253430 550898 253490 550936
rect 255589 550898 255655 550901
rect 253430 550896 255655 550898
rect 253430 550840 255594 550896
rect 255650 550840 255655 550896
rect 253430 550838 255655 550840
rect 255589 550835 255655 550838
rect 191741 550760 193690 550762
rect 191741 550704 191746 550760
rect 191802 550704 193690 550760
rect 191741 550702 193690 550704
rect 191741 550699 191807 550702
rect 69430 549540 69490 550120
rect 191649 549810 191715 549813
rect 193630 549810 193690 550392
rect 255589 549946 255655 549949
rect 253430 549944 255655 549946
rect 253430 549888 255594 549944
rect 255650 549888 255655 549944
rect 253430 549886 255655 549888
rect 253430 549848 253490 549886
rect 255589 549883 255655 549886
rect 191649 549808 193690 549810
rect 191649 549752 191654 549808
rect 191710 549752 193690 549808
rect 191649 549750 193690 549752
rect 191649 549747 191715 549750
rect 69422 549476 69428 549540
rect 69492 549476 69498 549540
rect 101254 549402 101260 549404
rect 94638 549342 101260 549402
rect 94638 549304 94698 549342
rect 101254 549340 101260 549342
rect 101324 549340 101330 549404
rect 191741 549402 191807 549405
rect 191741 549400 193690 549402
rect 191741 549344 191746 549400
rect 191802 549344 193690 549400
rect 191741 549342 193690 549344
rect 191741 549339 191807 549342
rect 193630 549304 193690 549342
rect 65977 548314 66043 548317
rect 68878 548314 68938 548760
rect 65977 548312 68938 548314
rect 65977 548256 65982 548312
rect 66038 548256 68938 548312
rect 65977 548254 68938 548256
rect 190637 548314 190703 548317
rect 193630 548314 193690 548488
rect 253430 548450 253490 549032
rect 255589 548450 255655 548453
rect 253430 548448 255655 548450
rect 253430 548392 255594 548448
rect 255650 548392 255655 548448
rect 253430 548390 255655 548392
rect 255589 548387 255655 548390
rect 190637 548312 193690 548314
rect 190637 548256 190642 548312
rect 190698 548256 193690 548312
rect 190637 548254 193690 548256
rect 65977 548251 66043 548254
rect 190637 548251 190703 548254
rect 253430 547906 253490 547944
rect 255865 547906 255931 547909
rect 253430 547904 255931 547906
rect 253430 547848 255870 547904
rect 255926 547848 255931 547904
rect 253430 547846 255931 547848
rect 255865 547843 255931 547846
rect 66161 546818 66227 546821
rect 68878 546818 68938 547400
rect 94638 547090 94698 547672
rect 96838 547090 96844 547092
rect 94638 547030 96844 547090
rect 96838 547028 96844 547030
rect 96908 547028 96914 547092
rect 191557 547090 191623 547093
rect 193630 547090 193690 547672
rect 191557 547088 193690 547090
rect 191557 547032 191562 547088
rect 191618 547032 193690 547088
rect 191557 547030 193690 547032
rect 191557 547027 191623 547030
rect 66161 546816 68938 546818
rect 66161 546760 66166 546816
rect 66222 546760 68938 546816
rect 66161 546758 68938 546760
rect 253430 546818 253490 547128
rect 255497 546818 255563 546821
rect 253430 546816 255563 546818
rect 253430 546760 255502 546816
rect 255558 546760 255563 546816
rect 253430 546758 255563 546760
rect 66161 546755 66227 546758
rect 255497 546755 255563 546758
rect 191649 546546 191715 546549
rect 193630 546546 193690 546584
rect 191649 546544 193690 546546
rect 191649 546488 191654 546544
rect 191710 546488 193690 546544
rect 191649 546486 193690 546488
rect 191649 546483 191715 546486
rect 67357 545458 67423 545461
rect 68878 545458 68938 546040
rect 94638 545730 94698 546312
rect 253430 545866 253490 546312
rect 255497 545866 255563 545869
rect 253430 545864 255563 545866
rect 253430 545808 255502 545864
rect 255558 545808 255563 545864
rect 253430 545806 255563 545808
rect 255497 545803 255563 545806
rect 97073 545730 97139 545733
rect 94638 545728 97139 545730
rect 94638 545672 97078 545728
rect 97134 545672 97139 545728
rect 94638 545670 97139 545672
rect 97073 545667 97139 545670
rect 67357 545456 68938 545458
rect 67357 545400 67362 545456
rect 67418 545400 68938 545456
rect 67357 545398 68938 545400
rect 67357 545395 67423 545398
rect 191649 545322 191715 545325
rect 193630 545322 193690 545768
rect 191649 545320 193690 545322
rect 191649 545264 191654 545320
rect 191710 545264 193690 545320
rect 191649 545262 193690 545264
rect 191649 545259 191715 545262
rect 253430 545186 253490 545224
rect 254209 545186 254275 545189
rect 253430 545184 254275 545186
rect 253430 545128 254214 545184
rect 254270 545128 254275 545184
rect 253430 545126 254275 545128
rect 254209 545123 254275 545126
rect 66805 544098 66871 544101
rect 68878 544098 68938 544680
rect 94638 544370 94698 544952
rect 97533 544370 97599 544373
rect 94638 544368 97599 544370
rect 94638 544312 97538 544368
rect 97594 544312 97599 544368
rect 94638 544310 97599 544312
rect 97533 544307 97599 544310
rect 191005 544234 191071 544237
rect 193630 544234 193690 544680
rect 191005 544232 193690 544234
rect 191005 544176 191010 544232
rect 191066 544176 193690 544232
rect 191005 544174 193690 544176
rect 191005 544171 191071 544174
rect 66805 544096 68938 544098
rect 66805 544040 66810 544096
rect 66866 544040 68938 544096
rect 66805 544038 68938 544040
rect 191557 544098 191623 544101
rect 191557 544096 193690 544098
rect 191557 544040 191562 544096
rect 191618 544040 193690 544096
rect 191557 544038 193690 544040
rect 66805 544035 66871 544038
rect 191557 544035 191623 544038
rect 193630 543864 193690 544038
rect 253430 543826 253490 544408
rect 256601 543826 256667 543829
rect 253430 543824 256667 543826
rect 253430 543768 256606 543824
rect 256662 543768 256667 543824
rect 253430 543766 256667 543768
rect 256601 543763 256667 543766
rect 66253 543418 66319 543421
rect 67950 543418 67956 543420
rect 66253 543416 67956 543418
rect 66253 543360 66258 543416
rect 66314 543360 67956 543416
rect 66253 543358 67956 543360
rect 66253 543355 66319 543358
rect 67950 543356 67956 543358
rect 68020 543418 68026 543420
rect 68020 543358 68938 543418
rect 68020 543356 68026 543358
rect 68878 543320 68938 543358
rect 94638 543010 94698 543592
rect 97533 543010 97599 543013
rect 94638 543008 97599 543010
rect 94638 542952 97538 543008
rect 97594 542952 97599 543008
rect 94638 542950 97599 542952
rect 97533 542947 97599 542950
rect 253430 542874 253490 543320
rect 255589 542874 255655 542877
rect 253430 542872 255655 542874
rect 253430 542816 255594 542872
rect 255650 542816 255655 542872
rect 253430 542814 255655 542816
rect 255589 542811 255655 542814
rect 188470 542404 188476 542468
rect 188540 542466 188546 542468
rect 193630 542466 193690 542776
rect 188540 542406 193690 542466
rect 253430 542466 253490 542504
rect 255497 542466 255563 542469
rect 253430 542464 255563 542466
rect 253430 542408 255502 542464
rect 255558 542408 255563 542464
rect 253430 542406 255563 542408
rect 188540 542404 188546 542406
rect 255497 542403 255563 542406
rect 66253 541378 66319 541381
rect 68878 541378 68938 541960
rect 94638 541786 94698 542232
rect 96889 541786 96955 541789
rect 97901 541786 97967 541789
rect 94638 541784 97967 541786
rect 94638 541728 96894 541784
rect 96950 541728 97906 541784
rect 97962 541728 97967 541784
rect 94638 541726 97967 541728
rect 96889 541723 96955 541726
rect 97901 541723 97967 541726
rect 66253 541376 68938 541378
rect 66253 541320 66258 541376
rect 66314 541320 68938 541376
rect 66253 541318 68938 541320
rect 66253 541315 66319 541318
rect 170489 541106 170555 541109
rect 193630 541106 193690 541960
rect 253430 541109 253490 541416
rect 170489 541104 193690 541106
rect 170489 541048 170494 541104
rect 170550 541048 193690 541104
rect 170489 541046 193690 541048
rect 253381 541104 253490 541109
rect 253381 541048 253386 541104
rect 253442 541048 253490 541104
rect 253381 541046 253490 541048
rect 170489 541043 170555 541046
rect 253381 541043 253447 541046
rect -960 540684 480 540924
rect 66253 540018 66319 540021
rect 68878 540018 68938 540600
rect 94638 540290 94698 540872
rect 193630 540698 193690 540872
rect 180750 540638 193690 540698
rect 94773 540290 94839 540293
rect 94638 540288 94839 540290
rect 94638 540232 94778 540288
rect 94834 540232 94839 540288
rect 94638 540230 94839 540232
rect 94773 540227 94839 540230
rect 66253 540016 68938 540018
rect 66253 539960 66258 540016
rect 66314 539960 68938 540016
rect 66253 539958 68938 539960
rect 66253 539955 66319 539958
rect 72918 539548 72924 539612
rect 72988 539610 72994 539612
rect 73061 539610 73127 539613
rect 76741 539610 76807 539613
rect 72988 539608 76807 539610
rect 72988 539552 73066 539608
rect 73122 539552 76746 539608
rect 76802 539552 76807 539608
rect 72988 539550 76807 539552
rect 72988 539548 72994 539550
rect 73061 539547 73127 539550
rect 76741 539547 76807 539550
rect 161238 539548 161244 539612
rect 161308 539610 161314 539612
rect 180750 539610 180810 540638
rect 191649 540562 191715 540565
rect 191649 540560 193690 540562
rect 191649 540504 191654 540560
rect 191710 540504 193690 540560
rect 191649 540502 193690 540504
rect 191649 540499 191715 540502
rect 193630 540056 193690 540502
rect 253430 540154 253490 540600
rect 255497 540154 255563 540157
rect 253430 540152 255563 540154
rect 253430 540096 255502 540152
rect 255558 540096 255563 540152
rect 253430 540094 255563 540096
rect 255497 540091 255563 540094
rect 161308 539550 180810 539610
rect 161308 539548 161314 539550
rect 69657 539068 69723 539069
rect 69606 539004 69612 539068
rect 69676 539066 69723 539068
rect 69676 539064 69768 539066
rect 69718 539008 69768 539064
rect 69676 539006 69768 539008
rect 69676 539004 69723 539006
rect 69657 539003 69723 539004
rect 94638 538933 94698 539512
rect 253430 539474 253490 539512
rect 255497 539474 255563 539477
rect 253430 539472 255563 539474
rect 253430 539416 255502 539472
rect 255558 539416 255563 539472
rect 253430 539414 255563 539416
rect 255497 539411 255563 539414
rect 188429 539338 188495 539341
rect 255262 539338 255268 539340
rect 188429 539336 255268 539338
rect 188429 539280 188434 539336
rect 188490 539280 255268 539336
rect 188429 539278 255268 539280
rect 188429 539275 188495 539278
rect 255262 539276 255268 539278
rect 255332 539276 255338 539340
rect 251214 539004 251220 539068
rect 251284 539066 251290 539068
rect 251449 539066 251515 539069
rect 251284 539064 251515 539066
rect 251284 539008 251454 539064
rect 251510 539008 251515 539064
rect 251284 539006 251515 539008
rect 251284 539004 251290 539006
rect 251449 539003 251515 539006
rect 94589 538928 94698 538933
rect 94589 538872 94594 538928
rect 94650 538872 94698 538928
rect 94589 538870 94698 538872
rect 94589 538867 94655 538870
rect 67357 538794 67423 538797
rect 81985 538794 82051 538797
rect 67357 538792 82051 538794
rect 67357 538736 67362 538792
rect 67418 538736 81990 538792
rect 82046 538736 82051 538792
rect 67357 538734 82051 538736
rect 67357 538731 67423 538734
rect 81985 538731 82051 538734
rect 80053 538386 80119 538389
rect 80053 538384 122850 538386
rect 80053 538328 80058 538384
rect 80114 538328 122850 538384
rect 80053 538326 122850 538328
rect 80053 538323 80119 538326
rect 122790 538250 122850 538326
rect 135897 538250 135963 538253
rect 207381 538250 207447 538253
rect 122790 538248 207447 538250
rect 122790 538192 135902 538248
rect 135958 538192 207386 538248
rect 207442 538192 207447 538248
rect 122790 538190 207447 538192
rect 135897 538187 135963 538190
rect 207381 538187 207447 538190
rect 84009 538114 84075 538117
rect 202965 538114 203031 538117
rect 84009 538112 203031 538114
rect 84009 538056 84014 538112
rect 84070 538056 202970 538112
rect 203026 538056 203031 538112
rect 84009 538054 203031 538056
rect 84009 538051 84075 538054
rect 202965 538051 203031 538054
rect 582373 537842 582439 537845
rect 583520 537842 584960 537932
rect 582373 537840 584960 537842
rect 582373 537784 582378 537840
rect 582434 537784 584960 537840
rect 582373 537782 584960 537784
rect 582373 537779 582439 537782
rect 583520 537692 584960 537782
rect 143625 537434 143691 537437
rect 222101 537434 222167 537437
rect 143625 537432 222167 537434
rect 143625 537376 143630 537432
rect 143686 537376 222106 537432
rect 222162 537376 222167 537432
rect 143625 537374 222167 537376
rect 143625 537371 143691 537374
rect 222101 537371 222167 537374
rect 245101 537434 245167 537437
rect 253974 537434 253980 537436
rect 245101 537432 253980 537434
rect 245101 537376 245106 537432
rect 245162 537376 253980 537432
rect 245101 537374 253980 537376
rect 245101 537371 245167 537374
rect 253974 537372 253980 537374
rect 254044 537372 254050 537436
rect 93393 536754 93459 536757
rect 246757 536754 246823 536757
rect 285581 536754 285647 536757
rect 93393 536752 285647 536754
rect 93393 536696 93398 536752
rect 93454 536696 246762 536752
rect 246818 536696 285586 536752
rect 285642 536696 285647 536752
rect 93393 536694 285647 536696
rect 93393 536691 93459 536694
rect 246757 536691 246823 536694
rect 285581 536691 285647 536694
rect 69657 536212 69723 536213
rect 69606 536210 69612 536212
rect 69566 536150 69612 536210
rect 69676 536208 69723 536212
rect 69718 536152 69723 536208
rect 69606 536148 69612 536150
rect 69676 536148 69723 536152
rect 69657 536147 69723 536148
rect 189073 536210 189139 536213
rect 193581 536210 193647 536213
rect 189073 536208 193647 536210
rect 189073 536152 189078 536208
rect 189134 536152 193586 536208
rect 193642 536152 193647 536208
rect 189073 536150 193647 536152
rect 189073 536147 189139 536150
rect 193581 536147 193647 536150
rect 182909 536074 182975 536077
rect 194133 536074 194199 536077
rect 182909 536072 194199 536074
rect 182909 536016 182914 536072
rect 182970 536016 194138 536072
rect 194194 536016 194199 536072
rect 182909 536014 194199 536016
rect 182909 536011 182975 536014
rect 194133 536011 194199 536014
rect 285581 536074 285647 536077
rect 295425 536074 295491 536077
rect 285581 536072 295491 536074
rect 285581 536016 285586 536072
rect 285642 536016 295430 536072
rect 295486 536016 295491 536072
rect 285581 536014 295491 536016
rect 285581 536011 285647 536014
rect 295425 536011 295491 536014
rect 68921 535530 68987 535533
rect 72417 535530 72483 535533
rect 68921 535528 72483 535530
rect 68921 535472 68926 535528
rect 68982 535472 72422 535528
rect 72478 535472 72483 535528
rect 68921 535470 72483 535472
rect 68921 535467 68987 535470
rect 72417 535467 72483 535470
rect 88190 535468 88196 535532
rect 88260 535530 88266 535532
rect 88333 535530 88399 535533
rect 88260 535528 88399 535530
rect 88260 535472 88338 535528
rect 88394 535472 88399 535528
rect 88260 535470 88399 535472
rect 88260 535468 88266 535470
rect 88333 535467 88399 535470
rect 196014 535468 196020 535532
rect 196084 535530 196090 535532
rect 197261 535530 197327 535533
rect 196084 535528 197327 535530
rect 196084 535472 197266 535528
rect 197322 535472 197327 535528
rect 196084 535470 197327 535472
rect 196084 535468 196090 535470
rect 197261 535467 197327 535470
rect 206277 535530 206343 535533
rect 208117 535530 208183 535533
rect 206277 535528 208183 535530
rect 206277 535472 206282 535528
rect 206338 535472 208122 535528
rect 208178 535472 208183 535528
rect 206277 535470 208183 535472
rect 206277 535467 206343 535470
rect 208117 535467 208183 535470
rect 217409 535530 217475 535533
rect 219525 535530 219591 535533
rect 217409 535528 219591 535530
rect 217409 535472 217414 535528
rect 217470 535472 219530 535528
rect 219586 535472 219591 535528
rect 217409 535470 219591 535472
rect 217409 535467 217475 535470
rect 219525 535467 219591 535470
rect 222929 535530 222995 535533
rect 226517 535530 226583 535533
rect 222929 535528 226583 535530
rect 222929 535472 222934 535528
rect 222990 535472 226522 535528
rect 226578 535472 226583 535528
rect 222929 535470 226583 535472
rect 222929 535467 222995 535470
rect 226517 535467 226583 535470
rect 244917 535530 244983 535533
rect 246297 535530 246363 535533
rect 244917 535528 246363 535530
rect 244917 535472 244922 535528
rect 244978 535472 246302 535528
rect 246358 535472 246363 535528
rect 244917 535470 246363 535472
rect 244917 535467 244983 535470
rect 246297 535467 246363 535470
rect 65885 535394 65951 535397
rect 224677 535394 224743 535397
rect 65885 535392 224743 535394
rect 65885 535336 65890 535392
rect 65946 535336 224682 535392
rect 224738 535336 224743 535392
rect 65885 535334 224743 535336
rect 65885 535331 65951 535334
rect 224677 535331 224743 535334
rect 223665 534170 223731 534173
rect 224677 534170 224743 534173
rect 223665 534168 224743 534170
rect 223665 534112 223670 534168
rect 223726 534112 224682 534168
rect 224738 534112 224743 534168
rect 223665 534110 224743 534112
rect 223665 534107 223731 534110
rect 224677 534107 224743 534110
rect 181529 534034 181595 534037
rect 199837 534034 199903 534037
rect 181529 534032 199903 534034
rect 181529 533976 181534 534032
rect 181590 533976 199842 534032
rect 199898 533976 199903 534032
rect 181529 533974 199903 533976
rect 181529 533971 181595 533974
rect 199837 533971 199903 533974
rect 213085 533490 213151 533493
rect 200070 533488 213151 533490
rect 200070 533432 213090 533488
rect 213146 533432 213151 533488
rect 200070 533430 213151 533432
rect 57697 533354 57763 533357
rect 84285 533354 84351 533357
rect 57697 533352 84351 533354
rect 57697 533296 57702 533352
rect 57758 533296 84290 533352
rect 84346 533296 84351 533352
rect 57697 533294 84351 533296
rect 57697 533291 57763 533294
rect 84285 533291 84351 533294
rect 152457 533354 152523 533357
rect 200070 533354 200130 533430
rect 213085 533427 213151 533430
rect 152457 533352 200130 533354
rect 152457 533296 152462 533352
rect 152518 533296 200130 533352
rect 152457 533294 200130 533296
rect 238201 533354 238267 533357
rect 273437 533354 273503 533357
rect 238201 533352 273503 533354
rect 238201 533296 238206 533352
rect 238262 533296 273442 533352
rect 273498 533296 273503 533352
rect 238201 533294 273503 533296
rect 152457 533291 152523 533294
rect 238201 533291 238267 533294
rect 273437 533291 273503 533294
rect 204897 532130 204963 532133
rect 212625 532130 212691 532133
rect 204897 532128 212691 532130
rect 204897 532072 204902 532128
rect 204958 532072 212630 532128
rect 212686 532072 212691 532128
rect 204897 532070 212691 532072
rect 204897 532067 204963 532070
rect 212625 532067 212691 532070
rect 211797 531994 211863 531997
rect 238518 531994 238524 531996
rect 211797 531992 238524 531994
rect 211797 531936 211802 531992
rect 211858 531936 238524 531992
rect 211797 531934 238524 531936
rect 211797 531931 211863 531934
rect 238518 531932 238524 531934
rect 238588 531932 238594 531996
rect 187601 530770 187667 530773
rect 218646 530770 218652 530772
rect 187601 530768 218652 530770
rect 187601 530712 187606 530768
rect 187662 530712 218652 530768
rect 187601 530710 218652 530712
rect 187601 530707 187667 530710
rect 218646 530708 218652 530710
rect 218716 530708 218722 530772
rect 218789 530770 218855 530773
rect 230606 530770 230612 530772
rect 218789 530768 230612 530770
rect 218789 530712 218794 530768
rect 218850 530712 230612 530768
rect 218789 530710 230612 530712
rect 218789 530707 218855 530710
rect 230606 530708 230612 530710
rect 230676 530708 230682 530772
rect 69790 530572 69796 530636
rect 69860 530634 69866 530636
rect 82854 530634 82860 530636
rect 69860 530574 82860 530634
rect 69860 530572 69866 530574
rect 82854 530572 82860 530574
rect 82924 530572 82930 530636
rect 85757 530634 85823 530637
rect 111742 530634 111748 530636
rect 85757 530632 111748 530634
rect 85757 530576 85762 530632
rect 85818 530576 111748 530632
rect 85757 530574 111748 530576
rect 85757 530571 85823 530574
rect 111742 530572 111748 530574
rect 111812 530572 111818 530636
rect 133781 530634 133847 530637
rect 189073 530634 189139 530637
rect 133781 530632 189139 530634
rect 133781 530576 133786 530632
rect 133842 530576 189078 530632
rect 189134 530576 189139 530632
rect 133781 530574 189139 530576
rect 133781 530571 133847 530574
rect 189073 530571 189139 530574
rect 197997 530634 198063 530637
rect 203333 530634 203399 530637
rect 197997 530632 203399 530634
rect 197997 530576 198002 530632
rect 198058 530576 203338 530632
rect 203394 530576 203399 530632
rect 197997 530574 203399 530576
rect 197997 530571 198063 530574
rect 203333 530571 203399 530574
rect 229737 530634 229803 530637
rect 256785 530634 256851 530637
rect 229737 530632 256851 530634
rect 229737 530576 229742 530632
rect 229798 530576 256790 530632
rect 256846 530576 256851 530632
rect 229737 530574 256851 530576
rect 229737 530571 229803 530574
rect 256785 530571 256851 530574
rect 67725 529274 67791 529277
rect 96654 529274 96660 529276
rect 67725 529272 96660 529274
rect 67725 529216 67730 529272
rect 67786 529216 96660 529272
rect 67725 529214 96660 529216
rect 67725 529211 67791 529214
rect 96654 529212 96660 529214
rect 96724 529212 96730 529276
rect 64689 529138 64755 529141
rect 252461 529138 252527 529141
rect 261017 529138 261083 529141
rect 64689 529136 261083 529138
rect 64689 529080 64694 529136
rect 64750 529080 252466 529136
rect 252522 529080 261022 529136
rect 261078 529080 261083 529136
rect 64689 529078 261083 529080
rect 64689 529075 64755 529078
rect 252461 529075 252527 529078
rect 261017 529075 261083 529078
rect 243169 528594 243235 528597
rect 248454 528594 248460 528596
rect 243169 528592 248460 528594
rect 243169 528536 243174 528592
rect 243230 528536 248460 528592
rect 243169 528534 248460 528536
rect 243169 528531 243235 528534
rect 248454 528532 248460 528534
rect 248524 528532 248530 528596
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 145557 527778 145623 527781
rect 220077 527778 220143 527781
rect 145557 527776 220143 527778
rect 145557 527720 145562 527776
rect 145618 527720 220082 527776
rect 220138 527720 220143 527776
rect 145557 527718 220143 527720
rect 145557 527715 145623 527718
rect 220077 527715 220143 527718
rect 66110 526356 66116 526420
rect 66180 526418 66186 526420
rect 96705 526418 96771 526421
rect 66180 526416 96771 526418
rect 66180 526360 96710 526416
rect 96766 526360 96771 526416
rect 66180 526358 96771 526360
rect 66180 526356 66186 526358
rect 96705 526355 96771 526358
rect 219934 526356 219940 526420
rect 220004 526418 220010 526420
rect 231117 526418 231183 526421
rect 220004 526416 231183 526418
rect 220004 526360 231122 526416
rect 231178 526360 231183 526416
rect 220004 526358 231183 526360
rect 220004 526356 220010 526358
rect 231117 526355 231183 526358
rect 249885 526418 249951 526421
rect 259545 526418 259611 526421
rect 249885 526416 259611 526418
rect 249885 526360 249890 526416
rect 249946 526360 259550 526416
rect 259606 526360 259611 526416
rect 249885 526358 259611 526360
rect 249885 526355 249951 526358
rect 259545 526355 259611 526358
rect 582741 524514 582807 524517
rect 583520 524514 584960 524604
rect 582741 524512 584960 524514
rect 582741 524456 582746 524512
rect 582802 524456 584960 524512
rect 582741 524454 584960 524456
rect 582741 524451 582807 524454
rect 583520 524364 584960 524454
rect 159950 523636 159956 523700
rect 160020 523698 160026 523700
rect 173249 523698 173315 523701
rect 160020 523696 173315 523698
rect 160020 523640 173254 523696
rect 173310 523640 173315 523696
rect 160020 523638 173315 523640
rect 160020 523636 160026 523638
rect 173249 523635 173315 523638
rect 224953 523698 225019 523701
rect 249742 523698 249748 523700
rect 224953 523696 249748 523698
rect 224953 523640 224958 523696
rect 225014 523640 249748 523696
rect 224953 523638 249748 523640
rect 224953 523635 225019 523638
rect 249742 523636 249748 523638
rect 249812 523636 249818 523700
rect 204989 522474 205055 522477
rect 219566 522474 219572 522476
rect 204989 522472 219572 522474
rect 204989 522416 204994 522472
rect 205050 522416 219572 522472
rect 204989 522414 219572 522416
rect 204989 522411 205055 522414
rect 219566 522412 219572 522414
rect 219636 522412 219642 522476
rect 203517 522338 203583 522341
rect 229686 522338 229692 522340
rect 203517 522336 229692 522338
rect 203517 522280 203522 522336
rect 203578 522280 229692 522336
rect 203517 522278 229692 522280
rect 203517 522275 203583 522278
rect 229686 522276 229692 522278
rect 229756 522276 229762 522340
rect 67950 521596 67956 521660
rect 68020 521658 68026 521660
rect 68870 521658 68876 521660
rect 68020 521598 68876 521658
rect 68020 521596 68026 521598
rect 68870 521596 68876 521598
rect 68940 521658 68946 521660
rect 258349 521658 258415 521661
rect 68940 521656 258415 521658
rect 68940 521600 258354 521656
rect 258410 521600 258415 521656
rect 68940 521598 258415 521600
rect 68940 521596 68946 521598
rect 258349 521595 258415 521598
rect 77150 520916 77156 520980
rect 77220 520978 77226 520980
rect 95325 520978 95391 520981
rect 77220 520976 95391 520978
rect 77220 520920 95330 520976
rect 95386 520920 95391 520976
rect 77220 520918 95391 520920
rect 77220 520916 77226 520918
rect 95325 520915 95391 520918
rect 61837 519482 61903 519485
rect 96838 519482 96844 519484
rect 61837 519480 96844 519482
rect 61837 519424 61842 519480
rect 61898 519424 96844 519480
rect 61837 519422 96844 519424
rect 61837 519419 61903 519422
rect 96838 519420 96844 519422
rect 96908 519420 96914 519484
rect 232446 518876 232452 518940
rect 232516 518938 232522 518940
rect 239397 518938 239463 518941
rect 232516 518936 239463 518938
rect 232516 518880 239402 518936
rect 239458 518880 239463 518936
rect 232516 518878 239463 518880
rect 232516 518876 232522 518878
rect 239397 518875 239463 518878
rect 69606 516700 69612 516764
rect 69676 516762 69682 516764
rect 115197 516762 115263 516765
rect 69676 516760 115263 516762
rect 69676 516704 115202 516760
rect 115258 516704 115263 516760
rect 69676 516702 115263 516704
rect 69676 516700 69682 516702
rect 115197 516699 115263 516702
rect 150341 515402 150407 515405
rect 184054 515402 184060 515404
rect 150341 515400 184060 515402
rect 150341 515344 150346 515400
rect 150402 515344 184060 515400
rect 150341 515342 184060 515344
rect 150341 515339 150407 515342
rect 184054 515340 184060 515342
rect 184124 515340 184130 515404
rect 194593 515402 194659 515405
rect 244406 515402 244412 515404
rect 194593 515400 244412 515402
rect 194593 515344 194598 515400
rect 194654 515344 244412 515400
rect 194593 515342 244412 515344
rect 194593 515339 194659 515342
rect 244406 515340 244412 515342
rect 244476 515340 244482 515404
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 72734 512620 72740 512684
rect 72804 512682 72810 512684
rect 95233 512682 95299 512685
rect 72804 512680 95299 512682
rect 72804 512624 95238 512680
rect 95294 512624 95299 512680
rect 72804 512622 95299 512624
rect 72804 512620 72810 512622
rect 95233 512619 95299 512622
rect 166206 512620 166212 512684
rect 166276 512682 166282 512684
rect 197353 512682 197419 512685
rect 166276 512680 197419 512682
rect 166276 512624 197358 512680
rect 197414 512624 197419 512680
rect 166276 512622 197419 512624
rect 166276 512620 166282 512622
rect 197353 512619 197419 512622
rect 195329 511458 195395 511461
rect 211654 511458 211660 511460
rect 195329 511456 211660 511458
rect 195329 511400 195334 511456
rect 195390 511400 211660 511456
rect 195329 511398 211660 511400
rect 195329 511395 195395 511398
rect 211654 511396 211660 511398
rect 211724 511396 211730 511460
rect 230974 511396 230980 511460
rect 231044 511458 231050 511460
rect 245694 511458 245700 511460
rect 231044 511398 245700 511458
rect 231044 511396 231050 511398
rect 245694 511396 245700 511398
rect 245764 511396 245770 511460
rect 210734 511260 210740 511324
rect 210804 511322 210810 511324
rect 232497 511322 232563 511325
rect 210804 511320 232563 511322
rect 210804 511264 232502 511320
rect 232558 511264 232563 511320
rect 210804 511262 232563 511264
rect 210804 511260 210810 511262
rect 232497 511259 232563 511262
rect 582649 511322 582715 511325
rect 583520 511322 584960 511412
rect 582649 511320 584960 511322
rect 582649 511264 582654 511320
rect 582710 511264 584960 511320
rect 582649 511262 584960 511264
rect 582649 511259 582715 511262
rect 583520 511172 584960 511262
rect 214649 509826 214715 509829
rect 226374 509826 226380 509828
rect 214649 509824 226380 509826
rect 214649 509768 214654 509824
rect 214710 509768 226380 509824
rect 214649 509766 226380 509768
rect 214649 509763 214715 509766
rect 226374 509764 226380 509766
rect 226444 509764 226450 509828
rect 227713 509826 227779 509829
rect 253054 509826 253060 509828
rect 227713 509824 253060 509826
rect 227713 509768 227718 509824
rect 227774 509768 253060 509824
rect 227713 509766 253060 509768
rect 227713 509763 227779 509766
rect 253054 509764 253060 509766
rect 253124 509764 253130 509828
rect 222694 505684 222700 505748
rect 222764 505746 222770 505748
rect 244273 505746 244339 505749
rect 222764 505744 244339 505746
rect 222764 505688 244278 505744
rect 244334 505688 244339 505744
rect 222764 505686 244339 505688
rect 222764 505684 222770 505686
rect 244273 505683 244339 505686
rect 150934 502964 150940 503028
rect 151004 503026 151010 503028
rect 197997 503026 198063 503029
rect 151004 503024 198063 503026
rect 151004 502968 198002 503024
rect 198058 502968 198063 503024
rect 151004 502966 198063 502968
rect 151004 502964 151010 502966
rect 197997 502963 198063 502966
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 75678 500108 75684 500172
rect 75748 500170 75754 500172
rect 94589 500170 94655 500173
rect 75748 500168 94655 500170
rect 75748 500112 94594 500168
rect 94650 500112 94655 500168
rect 75748 500110 94655 500112
rect 75748 500108 75754 500110
rect 94589 500107 94655 500110
rect 158621 498810 158687 498813
rect 188470 498810 188476 498812
rect 158621 498808 188476 498810
rect 158621 498752 158626 498808
rect 158682 498752 188476 498808
rect 158621 498750 188476 498752
rect 158621 498747 158687 498750
rect 188470 498748 188476 498750
rect 188540 498748 188546 498812
rect 204846 498748 204852 498812
rect 204916 498810 204922 498812
rect 241697 498810 241763 498813
rect 204916 498808 241763 498810
rect 204916 498752 241702 498808
rect 241758 498752 241763 498808
rect 204916 498750 241763 498752
rect 204916 498748 204922 498750
rect 241697 498747 241763 498750
rect 583520 497844 584960 498084
rect 161054 497388 161060 497452
rect 161124 497450 161130 497452
rect 222929 497450 222995 497453
rect 161124 497448 222995 497450
rect 161124 497392 222934 497448
rect 222990 497392 222995 497448
rect 161124 497390 222995 497392
rect 161124 497388 161130 497390
rect 222929 497387 222995 497390
rect 244365 496634 244431 496637
rect 244590 496634 244596 496636
rect 244365 496632 244596 496634
rect 244365 496576 244370 496632
rect 244426 496576 244596 496632
rect 244365 496574 244596 496576
rect 244365 496571 244431 496574
rect 244590 496572 244596 496574
rect 244660 496572 244666 496636
rect 140589 489970 140655 489973
rect 223798 489970 223804 489972
rect 140589 489968 223804 489970
rect 140589 489912 140594 489968
rect 140650 489912 223804 489968
rect 140589 489910 223804 489912
rect 140589 489907 140655 489910
rect 223798 489908 223804 489910
rect 223868 489908 223874 489972
rect 173617 489154 173683 489157
rect 251214 489154 251220 489156
rect 173617 489152 251220 489154
rect 173617 489096 173622 489152
rect 173678 489096 251220 489152
rect 173617 489094 251220 489096
rect 173617 489091 173683 489094
rect 251214 489092 251220 489094
rect 251284 489092 251290 489156
rect -960 488596 480 488836
rect 168966 486508 168972 486572
rect 169036 486570 169042 486572
rect 214649 486570 214715 486573
rect 169036 486568 214715 486570
rect 169036 486512 214654 486568
rect 214710 486512 214715 486568
rect 169036 486510 214715 486512
rect 169036 486508 169042 486510
rect 214649 486507 214715 486510
rect 197118 486372 197124 486436
rect 197188 486434 197194 486436
rect 254526 486434 254532 486436
rect 197188 486374 254532 486434
rect 197188 486372 197194 486374
rect 254526 486372 254532 486374
rect 254596 486372 254602 486436
rect 183461 485074 183527 485077
rect 207657 485074 207723 485077
rect 183461 485072 207723 485074
rect 183461 485016 183466 485072
rect 183522 485016 207662 485072
rect 207718 485016 207723 485072
rect 183461 485014 207723 485016
rect 183461 485011 183527 485014
rect 207657 485011 207723 485014
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 252553 484396 252619 484397
rect 252502 484332 252508 484396
rect 252572 484394 252619 484396
rect 252572 484392 252664 484394
rect 252614 484336 252664 484392
rect 252572 484334 252664 484336
rect 252572 484332 252619 484334
rect 252553 484331 252619 484332
rect 235901 483850 235967 483853
rect 252686 483850 252692 483852
rect 235901 483848 252692 483850
rect 235901 483792 235906 483848
rect 235962 483792 252692 483848
rect 235901 483790 252692 483792
rect 235901 483787 235967 483790
rect 252686 483788 252692 483790
rect 252756 483788 252762 483852
rect 163497 483714 163563 483717
rect 237414 483714 237420 483716
rect 163497 483712 237420 483714
rect 163497 483656 163502 483712
rect 163558 483656 237420 483712
rect 163497 483654 237420 483656
rect 163497 483651 163563 483654
rect 237414 483652 237420 483654
rect 237484 483652 237490 483716
rect 88977 482898 89043 482901
rect 89294 482898 89300 482900
rect 88977 482896 89300 482898
rect 88977 482840 88982 482896
rect 89038 482840 89300 482896
rect 88977 482838 89300 482840
rect 88977 482835 89043 482838
rect 89294 482836 89300 482838
rect 89364 482836 89370 482900
rect 196709 482218 196775 482221
rect 220854 482218 220860 482220
rect 196709 482216 220860 482218
rect 196709 482160 196714 482216
rect 196770 482160 220860 482216
rect 196709 482158 220860 482160
rect 196709 482155 196775 482158
rect 220854 482156 220860 482158
rect 220924 482156 220930 482220
rect 157149 481810 157215 481813
rect 249926 481810 249932 481812
rect 157149 481808 249932 481810
rect 157149 481752 157154 481808
rect 157210 481752 249932 481808
rect 157149 481750 249932 481752
rect 157149 481747 157215 481750
rect 249926 481748 249932 481750
rect 249996 481748 250002 481812
rect 88977 481674 89043 481677
rect 210509 481674 210575 481677
rect 88977 481672 210575 481674
rect 88977 481616 88982 481672
rect 89038 481616 210514 481672
rect 210570 481616 210575 481672
rect 88977 481614 210575 481616
rect 88977 481611 89043 481614
rect 210509 481611 210575 481614
rect 252461 481674 252527 481677
rect 285622 481674 285628 481676
rect 252461 481672 285628 481674
rect 252461 481616 252466 481672
rect 252522 481616 285628 481672
rect 252461 481614 285628 481616
rect 252461 481611 252527 481614
rect 285622 481612 285628 481614
rect 285692 481612 285698 481676
rect 240777 481540 240843 481541
rect 240726 481476 240732 481540
rect 240796 481538 240843 481540
rect 240796 481536 240888 481538
rect 240838 481480 240888 481536
rect 240796 481478 240888 481480
rect 240796 481476 240843 481478
rect 240777 481475 240843 481476
rect 202229 480858 202295 480861
rect 252461 480858 252527 480861
rect 202229 480856 252527 480858
rect 202229 480800 202234 480856
rect 202290 480800 252466 480856
rect 252522 480800 252527 480856
rect 202229 480798 252527 480800
rect 202229 480795 202295 480798
rect 252461 480795 252527 480798
rect 231853 478138 231919 478141
rect 262438 478138 262444 478140
rect 231853 478136 262444 478138
rect 231853 478080 231858 478136
rect 231914 478080 262444 478136
rect 231853 478078 262444 478080
rect 231853 478075 231919 478078
rect 262438 478076 262444 478078
rect 262508 478076 262514 478140
rect 178718 476716 178724 476780
rect 178788 476778 178794 476780
rect 217317 476778 217383 476781
rect 178788 476776 217383 476778
rect 178788 476720 217322 476776
rect 217378 476720 217383 476776
rect 178788 476718 217383 476720
rect 178788 476716 178794 476718
rect 217317 476715 217383 476718
rect 151077 476234 151143 476237
rect 151629 476234 151695 476237
rect 239489 476234 239555 476237
rect 151077 476232 239555 476234
rect 151077 476176 151082 476232
rect 151138 476176 151634 476232
rect 151690 476176 239494 476232
rect 239550 476176 239555 476232
rect 151077 476174 239555 476176
rect 151077 476171 151143 476174
rect 151629 476171 151695 476174
rect 239489 476171 239555 476174
rect 249374 476172 249380 476236
rect 249444 476234 249450 476236
rect 253289 476234 253355 476237
rect 249444 476232 253355 476234
rect 249444 476176 253294 476232
rect 253350 476176 253355 476232
rect 249444 476174 253355 476176
rect 249444 476172 249450 476174
rect 253289 476171 253355 476174
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 169569 475554 169635 475557
rect 192569 475554 192635 475557
rect 169569 475552 192635 475554
rect 169569 475496 169574 475552
rect 169630 475496 192574 475552
rect 192630 475496 192635 475552
rect 169569 475494 192635 475496
rect 169569 475491 169635 475494
rect 192569 475491 192635 475494
rect 187550 475356 187556 475420
rect 187620 475418 187626 475420
rect 218789 475418 218855 475421
rect 187620 475416 218855 475418
rect 187620 475360 218794 475416
rect 218850 475360 218855 475416
rect 187620 475358 218855 475360
rect 187620 475356 187626 475358
rect 218789 475355 218855 475358
rect 230473 475418 230539 475421
rect 258165 475418 258231 475421
rect 230473 475416 258231 475418
rect 230473 475360 230478 475416
rect 230534 475360 258170 475416
rect 258226 475360 258231 475416
rect 230473 475358 258231 475360
rect 230473 475355 230539 475358
rect 258165 475355 258231 475358
rect 180425 474194 180491 474197
rect 186814 474194 186820 474196
rect 180425 474192 186820 474194
rect 180425 474136 180430 474192
rect 180486 474136 186820 474192
rect 180425 474134 186820 474136
rect 180425 474131 180491 474134
rect 186814 474132 186820 474134
rect 186884 474132 186890 474196
rect 109033 474058 109099 474061
rect 109677 474058 109743 474061
rect 248597 474058 248663 474061
rect 249057 474058 249123 474061
rect 109033 474056 249123 474058
rect 109033 474000 109038 474056
rect 109094 474000 109682 474056
rect 109738 474000 248602 474056
rect 248658 474000 249062 474056
rect 249118 474000 249123 474056
rect 109033 473998 249123 474000
rect 109033 473995 109099 473998
rect 109677 473995 109743 473998
rect 248597 473995 248663 473998
rect 249057 473995 249123 473998
rect 181478 471820 181484 471884
rect 181548 471882 181554 471884
rect 189809 471882 189875 471885
rect 181548 471880 189875 471882
rect 181548 471824 189814 471880
rect 189870 471824 189875 471880
rect 181548 471822 189875 471824
rect 181548 471820 181554 471822
rect 189809 471819 189875 471822
rect 237373 471882 237439 471885
rect 238017 471882 238083 471885
rect 237373 471880 238083 471882
rect 237373 471824 237378 471880
rect 237434 471824 238022 471880
rect 238078 471824 238083 471880
rect 237373 471822 238083 471824
rect 237373 471819 237439 471822
rect 238017 471819 238083 471822
rect 582465 471474 582531 471477
rect 583520 471474 584960 471564
rect 582465 471472 584960 471474
rect 582465 471416 582470 471472
rect 582526 471416 584960 471472
rect 582465 471414 584960 471416
rect 582465 471411 582531 471414
rect 173566 471276 173572 471340
rect 173636 471338 173642 471340
rect 211797 471338 211863 471341
rect 173636 471336 211863 471338
rect 173636 471280 211802 471336
rect 211858 471280 211863 471336
rect 583520 471324 584960 471414
rect 173636 471278 211863 471280
rect 173636 471276 173642 471278
rect 211797 471275 211863 471278
rect 158713 471202 158779 471205
rect 159357 471202 159423 471205
rect 239397 471202 239463 471205
rect 158713 471200 239463 471202
rect 158713 471144 158718 471200
rect 158774 471144 159362 471200
rect 159418 471144 239402 471200
rect 239458 471144 239463 471200
rect 158713 471142 239463 471144
rect 158713 471139 158779 471142
rect 159357 471139 159423 471142
rect 239397 471139 239463 471142
rect 237373 470658 237439 470661
rect 294045 470658 294111 470661
rect 237373 470656 294111 470658
rect 237373 470600 237378 470656
rect 237434 470600 294050 470656
rect 294106 470600 294111 470656
rect 237373 470598 294111 470600
rect 237373 470595 237439 470598
rect 294045 470595 294111 470598
rect 187509 469842 187575 469845
rect 216673 469842 216739 469845
rect 187509 469840 216739 469842
rect 187509 469784 187514 469840
rect 187570 469784 216678 469840
rect 216734 469784 216739 469840
rect 187509 469782 216739 469784
rect 187509 469779 187575 469782
rect 216673 469779 216739 469782
rect 165521 469298 165587 469301
rect 173157 469298 173223 469301
rect 165521 469296 173223 469298
rect 165521 469240 165526 469296
rect 165582 469240 173162 469296
rect 173218 469240 173223 469296
rect 165521 469238 173223 469240
rect 165521 469235 165587 469238
rect 173157 469235 173223 469238
rect 173750 469236 173756 469300
rect 173820 469298 173826 469300
rect 180006 469298 180012 469300
rect 173820 469238 180012 469298
rect 173820 469236 173826 469238
rect 180006 469236 180012 469238
rect 180076 469236 180082 469300
rect 162526 468420 162532 468484
rect 162596 468482 162602 468484
rect 177389 468482 177455 468485
rect 162596 468480 177455 468482
rect 162596 468424 177394 468480
rect 177450 468424 177455 468480
rect 162596 468422 177455 468424
rect 162596 468420 162602 468422
rect 177389 468419 177455 468422
rect 177573 468482 177639 468485
rect 206277 468482 206343 468485
rect 177573 468480 206343 468482
rect 177573 468424 177578 468480
rect 177634 468424 206282 468480
rect 206338 468424 206343 468480
rect 177573 468422 206343 468424
rect 177573 468419 177639 468422
rect 206277 468419 206343 468422
rect 187693 468074 187759 468077
rect 227713 468074 227779 468077
rect 187693 468072 227779 468074
rect 187693 468016 187698 468072
rect 187754 468016 227718 468072
rect 227774 468016 227779 468072
rect 187693 468014 227779 468016
rect 187693 468011 187759 468014
rect 227713 468011 227779 468014
rect 68921 467940 68987 467941
rect 68870 467938 68876 467940
rect 68830 467878 68876 467938
rect 68940 467938 68987 467940
rect 187785 467938 187851 467941
rect 68940 467936 187851 467938
rect 68982 467880 187790 467936
rect 187846 467880 187851 467936
rect 68870 467876 68876 467878
rect 68940 467878 187851 467880
rect 68940 467876 68987 467878
rect 68921 467875 68987 467876
rect 187785 467875 187851 467878
rect 212625 467938 212691 467941
rect 213269 467938 213335 467941
rect 287237 467938 287303 467941
rect 212625 467936 287303 467938
rect 212625 467880 212630 467936
rect 212686 467880 213274 467936
rect 213330 467880 287242 467936
rect 287298 467880 287303 467936
rect 212625 467878 287303 467880
rect 212625 467875 212691 467878
rect 213269 467875 213335 467878
rect 287237 467875 287303 467878
rect 190310 467060 190316 467124
rect 190380 467122 190386 467124
rect 203006 467122 203012 467124
rect 190380 467062 203012 467122
rect 190380 467060 190386 467062
rect 203006 467060 203012 467062
rect 203076 467060 203082 467124
rect 66110 466516 66116 466580
rect 66180 466578 66186 466580
rect 153929 466578 153995 466581
rect 66180 466576 153995 466578
rect 66180 466520 153934 466576
rect 153990 466520 153995 466576
rect 66180 466518 153995 466520
rect 66180 466516 66186 466518
rect 153929 466515 153995 466518
rect 155217 466578 155283 466581
rect 255262 466578 255268 466580
rect 155217 466576 255268 466578
rect 155217 466520 155222 466576
rect 155278 466520 255268 466576
rect 155217 466518 255268 466520
rect 155217 466515 155283 466518
rect 255262 466516 255268 466518
rect 255332 466516 255338 466580
rect 170990 465836 170996 465900
rect 171060 465898 171066 465900
rect 201534 465898 201540 465900
rect 171060 465838 201540 465898
rect 171060 465836 171066 465838
rect 201534 465836 201540 465838
rect 201604 465836 201610 465900
rect 218697 465898 218763 465901
rect 236494 465898 236500 465900
rect 218697 465896 236500 465898
rect 218697 465840 218702 465896
rect 218758 465840 236500 465896
rect 218697 465838 236500 465840
rect 218697 465835 218763 465838
rect 236494 465836 236500 465838
rect 236564 465836 236570 465900
rect 67766 465700 67772 465764
rect 67836 465762 67842 465764
rect 91318 465762 91324 465764
rect 67836 465702 91324 465762
rect 67836 465700 67842 465702
rect 91318 465700 91324 465702
rect 91388 465700 91394 465764
rect 151261 465762 151327 465765
rect 187601 465762 187667 465765
rect 151261 465760 187667 465762
rect 151261 465704 151266 465760
rect 151322 465704 187606 465760
rect 187662 465704 187667 465760
rect 151261 465702 187667 465704
rect 151261 465699 151327 465702
rect 187601 465699 187667 465702
rect 197353 465762 197419 465765
rect 223982 465762 223988 465764
rect 197353 465760 223988 465762
rect 197353 465704 197358 465760
rect 197414 465704 223988 465760
rect 197353 465702 223988 465704
rect 197353 465699 197419 465702
rect 223982 465700 223988 465702
rect 224052 465700 224058 465764
rect 232497 465626 232563 465629
rect 233233 465626 233299 465629
rect 232497 465624 233299 465626
rect 232497 465568 232502 465624
rect 232558 465568 233238 465624
rect 233294 465568 233299 465624
rect 232497 465566 233299 465568
rect 232497 465563 232563 465566
rect 233233 465563 233299 465566
rect 233233 465218 233299 465221
rect 299473 465218 299539 465221
rect 233233 465216 299539 465218
rect 233233 465160 233238 465216
rect 233294 465160 299478 465216
rect 299534 465160 299539 465216
rect 233233 465158 299539 465160
rect 233233 465155 233299 465158
rect 299473 465155 299539 465158
rect 204161 464538 204227 464541
rect 215334 464538 215340 464540
rect 204161 464536 215340 464538
rect 204161 464480 204166 464536
rect 204222 464480 215340 464536
rect 204161 464478 215340 464480
rect 204161 464475 204227 464478
rect 215334 464476 215340 464478
rect 215404 464476 215410 464540
rect 176510 464340 176516 464404
rect 176580 464402 176586 464404
rect 205081 464402 205147 464405
rect 176580 464400 205147 464402
rect 176580 464344 205086 464400
rect 205142 464344 205147 464400
rect 176580 464342 205147 464344
rect 176580 464340 176586 464342
rect 205081 464339 205147 464342
rect 215477 464402 215543 464405
rect 223798 464402 223804 464404
rect 215477 464400 223804 464402
rect 215477 464344 215482 464400
rect 215538 464344 223804 464400
rect 215477 464342 223804 464344
rect 215477 464339 215543 464342
rect 223798 464340 223804 464342
rect 223868 464340 223874 464404
rect 146201 463722 146267 463725
rect 216765 463722 216831 463725
rect 146201 463720 216831 463722
rect 146201 463664 146206 463720
rect 146262 463664 216770 463720
rect 216826 463664 216831 463720
rect 146201 463662 216831 463664
rect 146201 463659 146267 463662
rect 216765 463659 216831 463662
rect 224953 463722 225019 463725
rect 226241 463722 226307 463725
rect 280153 463722 280219 463725
rect 224953 463720 280219 463722
rect 224953 463664 224958 463720
rect 225014 463664 226246 463720
rect 226302 463664 280158 463720
rect 280214 463664 280219 463720
rect 224953 463662 280219 463664
rect 224953 463659 225019 463662
rect 226241 463659 226307 463662
rect 280153 463659 280219 463662
rect 115197 463586 115263 463589
rect 235993 463586 236059 463589
rect 115197 463584 236059 463586
rect 115197 463528 115202 463584
rect 115258 463528 235998 463584
rect 236054 463528 236059 463584
rect 115197 463526 236059 463528
rect 115197 463523 115263 463526
rect 235993 463523 236059 463526
rect 241605 463586 241671 463589
rect 242157 463586 242223 463589
rect 241605 463584 242223 463586
rect 241605 463528 241610 463584
rect 241666 463528 242162 463584
rect 242218 463528 242223 463584
rect 241605 463526 242223 463528
rect 241605 463523 241671 463526
rect 242157 463523 242223 463526
rect 66161 462906 66227 462909
rect 104198 462906 104204 462908
rect 66161 462904 104204 462906
rect 66161 462848 66166 462904
rect 66222 462848 104204 462904
rect 66161 462846 104204 462848
rect 66161 462843 66227 462846
rect 104198 462844 104204 462846
rect 104268 462844 104274 462908
rect 177614 462844 177620 462908
rect 177684 462906 177690 462908
rect 207054 462906 207060 462908
rect 177684 462846 207060 462906
rect 177684 462844 177690 462846
rect 207054 462844 207060 462846
rect 207124 462844 207130 462908
rect 239489 462906 239555 462909
rect 254209 462906 254275 462909
rect 239489 462904 254275 462906
rect 239489 462848 239494 462904
rect 239550 462848 254214 462904
rect 254270 462848 254275 462904
rect 239489 462846 254275 462848
rect 239489 462843 239555 462846
rect 254209 462843 254275 462846
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 241605 462362 241671 462365
rect 299565 462362 299631 462365
rect 241605 462360 299631 462362
rect 241605 462304 241610 462360
rect 241666 462304 299570 462360
rect 299626 462304 299631 462360
rect 241605 462302 299631 462304
rect 241605 462299 241671 462302
rect 299565 462299 299631 462302
rect 201585 462226 201651 462229
rect 202229 462226 202295 462229
rect 201585 462224 202295 462226
rect 201585 462168 201590 462224
rect 201646 462168 202234 462224
rect 202290 462168 202295 462224
rect 201585 462166 202295 462168
rect 201585 462163 201651 462166
rect 202229 462163 202295 462166
rect 234613 462226 234679 462229
rect 235901 462226 235967 462229
rect 234613 462224 235967 462226
rect 234613 462168 234618 462224
rect 234674 462168 235906 462224
rect 235962 462168 235967 462224
rect 234613 462166 235967 462168
rect 234613 462163 234679 462166
rect 235901 462163 235967 462166
rect 187785 461682 187851 461685
rect 208393 461682 208459 461685
rect 187785 461680 208459 461682
rect 187785 461624 187790 461680
rect 187846 461624 208398 461680
rect 208454 461624 208459 461680
rect 187785 461622 208459 461624
rect 187785 461619 187851 461622
rect 208393 461619 208459 461622
rect 158529 461546 158595 461549
rect 195329 461546 195395 461549
rect 158529 461544 195395 461546
rect 158529 461488 158534 461544
rect 158590 461488 195334 461544
rect 195390 461488 195395 461544
rect 158529 461486 195395 461488
rect 158529 461483 158595 461486
rect 195329 461483 195395 461486
rect 202321 461546 202387 461549
rect 222837 461546 222903 461549
rect 202321 461544 222903 461546
rect 202321 461488 202326 461544
rect 202382 461488 222842 461544
rect 222898 461488 222903 461544
rect 202321 461486 222903 461488
rect 202321 461483 202387 461486
rect 222837 461483 222903 461486
rect 75729 461002 75795 461005
rect 201585 461002 201651 461005
rect 75729 461000 201651 461002
rect 75729 460944 75734 461000
rect 75790 460944 201590 461000
rect 201646 460944 201651 461000
rect 75729 460942 201651 460944
rect 75729 460939 75795 460942
rect 201585 460939 201651 460942
rect 235901 461002 235967 461005
rect 269389 461002 269455 461005
rect 235901 461000 269455 461002
rect 235901 460944 235906 461000
rect 235962 460944 269394 461000
rect 269450 460944 269455 461000
rect 235901 460942 269455 460944
rect 235901 460939 235967 460942
rect 269389 460939 269455 460942
rect 74533 460186 74599 460189
rect 152917 460186 152983 460189
rect 188429 460186 188495 460189
rect 74533 460184 188495 460186
rect 74533 460128 74538 460184
rect 74594 460128 152922 460184
rect 152978 460128 188434 460184
rect 188490 460128 188495 460184
rect 74533 460126 188495 460128
rect 74533 460123 74599 460126
rect 152917 460123 152983 460126
rect 188429 460123 188495 460126
rect 184197 459914 184263 459917
rect 218053 459914 218119 459917
rect 218697 459914 218763 459917
rect 184197 459912 218763 459914
rect 184197 459856 184202 459912
rect 184258 459856 218058 459912
rect 218114 459856 218702 459912
rect 218758 459856 218763 459912
rect 184197 459854 218763 459856
rect 184197 459851 184263 459854
rect 218053 459851 218119 459854
rect 218697 459851 218763 459854
rect 215937 459778 216003 459781
rect 288433 459778 288499 459781
rect 215937 459776 288499 459778
rect 215937 459720 215942 459776
rect 215998 459720 288438 459776
rect 288494 459720 288499 459776
rect 215937 459718 288499 459720
rect 215937 459715 216003 459718
rect 288433 459715 288499 459718
rect 187693 459642 187759 459645
rect 273529 459642 273595 459645
rect 187693 459640 273595 459642
rect 187693 459584 187698 459640
rect 187754 459584 273534 459640
rect 273590 459584 273595 459640
rect 187693 459582 273595 459584
rect 187693 459579 187759 459582
rect 273529 459579 273595 459582
rect 188838 459036 188844 459100
rect 188908 459098 188914 459100
rect 196617 459098 196683 459101
rect 188908 459096 196683 459098
rect 188908 459040 196622 459096
rect 196678 459040 196683 459096
rect 188908 459038 196683 459040
rect 188908 459036 188914 459038
rect 196617 459035 196683 459038
rect 201401 459098 201467 459101
rect 233182 459098 233188 459100
rect 201401 459096 233188 459098
rect 201401 459040 201406 459096
rect 201462 459040 233188 459096
rect 201401 459038 233188 459040
rect 201401 459035 201467 459038
rect 233182 459036 233188 459038
rect 233252 459036 233258 459100
rect 195053 458962 195119 458965
rect 234654 458962 234660 458964
rect 195053 458960 234660 458962
rect 195053 458904 195058 458960
rect 195114 458904 234660 458960
rect 195053 458902 234660 458904
rect 195053 458899 195119 458902
rect 234654 458900 234660 458902
rect 234724 458900 234730 458964
rect 184790 458764 184796 458828
rect 184860 458826 184866 458828
rect 204989 458826 205055 458829
rect 184860 458824 205055 458826
rect 184860 458768 204994 458824
rect 205050 458768 205055 458824
rect 184860 458766 205055 458768
rect 184860 458764 184866 458766
rect 204989 458763 205055 458766
rect 232129 458826 232195 458829
rect 233141 458826 233207 458829
rect 277485 458826 277551 458829
rect 277761 458826 277827 458829
rect 232129 458824 277827 458826
rect 232129 458768 232134 458824
rect 232190 458768 233146 458824
rect 233202 458768 277490 458824
rect 277546 458768 277766 458824
rect 277822 458768 277827 458824
rect 232129 458766 277827 458768
rect 232129 458763 232195 458766
rect 233141 458763 233207 458766
rect 277485 458763 277551 458766
rect 277761 458763 277827 458766
rect 237465 458282 237531 458285
rect 238109 458282 238175 458285
rect 298185 458282 298251 458285
rect 237465 458280 298251 458282
rect 237465 458224 237470 458280
rect 237526 458224 238114 458280
rect 238170 458224 298190 458280
rect 298246 458224 298251 458280
rect 237465 458222 298251 458224
rect 237465 458219 237531 458222
rect 238109 458219 238175 458222
rect 298185 458219 298251 458222
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 80053 457466 80119 457469
rect 114318 457466 114324 457468
rect 80053 457464 114324 457466
rect 80053 457408 80058 457464
rect 80114 457408 114324 457464
rect 80053 457406 114324 457408
rect 80053 457403 80119 457406
rect 114318 457404 114324 457406
rect 114388 457404 114394 457468
rect 240777 457466 240843 457469
rect 255589 457466 255655 457469
rect 240777 457464 255655 457466
rect 240777 457408 240782 457464
rect 240838 457408 255594 457464
rect 255650 457408 255655 457464
rect 240777 457406 255655 457408
rect 240777 457403 240843 457406
rect 255589 457403 255655 457406
rect 118601 456922 118667 456925
rect 223665 456922 223731 456925
rect 118601 456920 223731 456922
rect 118601 456864 118606 456920
rect 118662 456864 223670 456920
rect 223726 456864 223731 456920
rect 118601 456862 223731 456864
rect 118601 456859 118667 456862
rect 223665 456859 223731 456862
rect 231209 456922 231275 456925
rect 289813 456922 289879 456925
rect 231209 456920 289879 456922
rect 231209 456864 231214 456920
rect 231270 456864 289818 456920
rect 289874 456864 289879 456920
rect 231209 456862 289879 456864
rect 231209 456859 231275 456862
rect 289813 456859 289879 456862
rect 180558 456316 180564 456380
rect 180628 456378 180634 456380
rect 196709 456378 196775 456381
rect 180628 456376 196775 456378
rect 180628 456320 196714 456376
rect 196770 456320 196775 456376
rect 180628 456318 196775 456320
rect 180628 456316 180634 456318
rect 196709 456315 196775 456318
rect 191649 456242 191715 456245
rect 228214 456242 228220 456244
rect 191649 456240 228220 456242
rect 191649 456184 191654 456240
rect 191710 456184 228220 456240
rect 191649 456182 228220 456184
rect 191649 456179 191715 456182
rect 228214 456180 228220 456182
rect 228284 456180 228290 456244
rect 151169 456106 151235 456109
rect 187693 456106 187759 456109
rect 151169 456104 187759 456106
rect 151169 456048 151174 456104
rect 151230 456048 187698 456104
rect 187754 456048 187759 456104
rect 151169 456046 187759 456048
rect 151169 456043 151235 456046
rect 187693 456043 187759 456046
rect 191557 456106 191623 456109
rect 247718 456106 247724 456108
rect 191557 456104 247724 456106
rect 191557 456048 191562 456104
rect 191618 456048 247724 456104
rect 191557 456046 247724 456048
rect 191557 456043 191623 456046
rect 247718 456044 247724 456046
rect 247788 456044 247794 456108
rect 232589 455562 232655 455565
rect 287329 455562 287395 455565
rect 288341 455562 288407 455565
rect 232589 455560 288407 455562
rect 232589 455504 232594 455560
rect 232650 455504 287334 455560
rect 287390 455504 288346 455560
rect 288402 455504 288407 455560
rect 232589 455502 288407 455504
rect 232589 455499 232655 455502
rect 287329 455499 287395 455502
rect 288341 455499 288407 455502
rect 250294 455364 250300 455428
rect 250364 455426 250370 455428
rect 252093 455426 252159 455429
rect 250364 455424 252159 455426
rect 250364 455368 252098 455424
rect 252154 455368 252159 455424
rect 250364 455366 252159 455368
rect 250364 455364 250370 455366
rect 252093 455363 252159 455366
rect 73153 454746 73219 454749
rect 112294 454746 112300 454748
rect 73153 454744 112300 454746
rect 73153 454688 73158 454744
rect 73214 454688 112300 454744
rect 73153 454686 112300 454688
rect 73153 454683 73219 454686
rect 112294 454684 112300 454686
rect 112364 454684 112370 454748
rect 181897 454746 181963 454749
rect 204897 454746 204963 454749
rect 181897 454744 204963 454746
rect 181897 454688 181902 454744
rect 181958 454688 204902 454744
rect 204958 454688 204963 454744
rect 181897 454686 204963 454688
rect 181897 454683 181963 454686
rect 204897 454683 204963 454686
rect 222101 454202 222167 454205
rect 265617 454202 265683 454205
rect 222101 454200 265683 454202
rect 222101 454144 222106 454200
rect 222162 454144 265622 454200
rect 265678 454144 265683 454200
rect 222101 454142 265683 454144
rect 222101 454139 222167 454142
rect 265617 454139 265683 454142
rect 147581 454066 147647 454069
rect 197905 454066 197971 454069
rect 147581 454064 197971 454066
rect 147581 454008 147586 454064
rect 147642 454008 197910 454064
rect 197966 454008 197971 454064
rect 147581 454006 197971 454008
rect 147581 454003 147647 454006
rect 197905 454003 197971 454006
rect 223665 454066 223731 454069
rect 284334 454066 284340 454068
rect 223665 454064 284340 454066
rect 223665 454008 223670 454064
rect 223726 454008 284340 454064
rect 223665 454006 284340 454008
rect 223665 454003 223731 454006
rect 284334 454004 284340 454006
rect 284404 454004 284410 454068
rect 172513 453930 172579 453933
rect 173566 453930 173572 453932
rect 172513 453928 173572 453930
rect 172513 453872 172518 453928
rect 172574 453872 173572 453928
rect 172513 453870 173572 453872
rect 172513 453867 172579 453870
rect 173566 453868 173572 453870
rect 173636 453868 173642 453932
rect 173566 453732 173572 453796
rect 173636 453794 173642 453796
rect 176101 453794 176167 453797
rect 173636 453792 176167 453794
rect 173636 453736 176106 453792
rect 176162 453736 176167 453792
rect 173636 453734 176167 453736
rect 173636 453732 173642 453734
rect 176101 453731 176167 453734
rect 74441 452978 74507 452981
rect 200849 452978 200915 452981
rect 201401 452978 201467 452981
rect 74441 452976 201467 452978
rect 74441 452920 74446 452976
rect 74502 452920 200854 452976
rect 200910 452920 201406 452976
rect 201462 452920 201467 452976
rect 74441 452918 201467 452920
rect 74441 452915 74507 452918
rect 200849 452915 200915 452918
rect 201401 452915 201467 452918
rect 251541 452978 251607 452981
rect 261017 452978 261083 452981
rect 251541 452976 261083 452978
rect 251541 452920 251546 452976
rect 251602 452920 261022 452976
rect 261078 452920 261083 452976
rect 251541 452918 261083 452920
rect 251541 452915 251607 452918
rect 261017 452915 261083 452918
rect 119337 452842 119403 452845
rect 233233 452842 233299 452845
rect 119337 452840 233299 452842
rect 119337 452784 119342 452840
rect 119398 452784 233238 452840
rect 233294 452784 233299 452840
rect 119337 452782 233299 452784
rect 119337 452779 119403 452782
rect 233233 452779 233299 452782
rect 238845 452842 238911 452845
rect 244917 452842 244983 452845
rect 278773 452842 278839 452845
rect 238845 452840 278839 452842
rect 238845 452784 238850 452840
rect 238906 452784 244922 452840
rect 244978 452784 278778 452840
rect 278834 452784 278839 452840
rect 238845 452782 278839 452784
rect 238845 452779 238911 452782
rect 244917 452779 244983 452782
rect 278773 452779 278839 452782
rect 188429 452706 188495 452709
rect 195605 452706 195671 452709
rect 203149 452706 203215 452709
rect 273437 452706 273503 452709
rect 188429 452704 195671 452706
rect 188429 452648 188434 452704
rect 188490 452648 195610 452704
rect 195666 452648 195671 452704
rect 188429 452646 195671 452648
rect 188429 452643 188495 452646
rect 195605 452643 195671 452646
rect 203014 452704 273503 452706
rect 203014 452648 203154 452704
rect 203210 452648 273442 452704
rect 273498 452648 273503 452704
rect 203014 452646 273503 452648
rect 176653 452570 176719 452573
rect 177297 452570 177363 452573
rect 176653 452568 177363 452570
rect 176653 452512 176658 452568
rect 176714 452512 177302 452568
rect 177358 452512 177363 452568
rect 176653 452510 177363 452512
rect 176653 452507 176719 452510
rect 177297 452507 177363 452510
rect 186221 452570 186287 452573
rect 203014 452570 203074 452646
rect 203149 452643 203215 452646
rect 273437 452643 273503 452646
rect 186221 452568 203074 452570
rect 186221 452512 186226 452568
rect 186282 452512 203074 452568
rect 186221 452510 203074 452512
rect 251081 452570 251147 452573
rect 287053 452570 287119 452573
rect 288525 452570 288591 452573
rect 251081 452568 288591 452570
rect 251081 452512 251086 452568
rect 251142 452512 287058 452568
rect 287114 452512 288530 452568
rect 288586 452512 288591 452568
rect 251081 452510 288591 452512
rect 186221 452507 186287 452510
rect 251081 452507 251147 452510
rect 287053 452507 287119 452510
rect 288525 452507 288591 452510
rect 184749 452434 184815 452437
rect 187141 452434 187207 452437
rect 273253 452436 273319 452437
rect 273253 452434 273300 452436
rect 184749 452432 187207 452434
rect 184749 452376 184754 452432
rect 184810 452376 187146 452432
rect 187202 452376 187207 452432
rect 184749 452374 187207 452376
rect 273208 452432 273300 452434
rect 273208 452376 273258 452432
rect 273208 452374 273300 452376
rect 184749 452371 184815 452374
rect 187141 452371 187207 452374
rect 273253 452372 273300 452374
rect 273364 452372 273370 452436
rect 273253 452371 273319 452372
rect 67449 451890 67515 451893
rect 176653 451890 176719 451893
rect 67449 451888 176719 451890
rect 67449 451832 67454 451888
rect 67510 451832 176658 451888
rect 176714 451832 176719 451888
rect 67449 451830 176719 451832
rect 67449 451827 67515 451830
rect 176653 451827 176719 451830
rect 228725 451618 228791 451621
rect 270677 451618 270743 451621
rect 228725 451616 270743 451618
rect 228725 451560 228730 451616
rect 228786 451560 270682 451616
rect 270738 451560 270743 451616
rect 228725 451558 270743 451560
rect 228725 451555 228791 451558
rect 270677 451555 270743 451558
rect 186313 451482 186379 451485
rect 187141 451482 187207 451485
rect 250621 451482 250687 451485
rect 186313 451480 250687 451482
rect 186313 451424 186318 451480
rect 186374 451424 187146 451480
rect 187202 451424 250626 451480
rect 250682 451424 250687 451480
rect 186313 451422 250687 451424
rect 186313 451419 186379 451422
rect 187141 451419 187207 451422
rect 250621 451419 250687 451422
rect 204069 451346 204135 451349
rect 273069 451346 273135 451349
rect 204069 451344 273135 451346
rect 204069 451288 204074 451344
rect 204130 451288 273074 451344
rect 273130 451288 273135 451344
rect 204069 451286 273135 451288
rect 204069 451283 204135 451286
rect 273069 451283 273135 451286
rect 166349 451210 166415 451213
rect 238845 451210 238911 451213
rect 166349 451208 238911 451210
rect 166349 451152 166354 451208
rect 166410 451152 238850 451208
rect 238906 451152 238911 451208
rect 166349 451150 238911 451152
rect 166349 451147 166415 451150
rect 238845 451147 238911 451150
rect 233877 450666 233943 450669
rect 247166 450666 247172 450668
rect 233877 450664 247172 450666
rect 233877 450608 233882 450664
rect 233938 450608 247172 450664
rect 233877 450606 247172 450608
rect 233877 450603 233943 450606
rect 247166 450604 247172 450606
rect 247236 450604 247242 450668
rect 106273 450530 106339 450533
rect 166349 450530 166415 450533
rect 106273 450528 166415 450530
rect 106273 450472 106278 450528
rect 106334 450472 166354 450528
rect 166410 450472 166415 450528
rect 106273 450470 166415 450472
rect 106273 450467 106339 450470
rect 166349 450467 166415 450470
rect 244273 450530 244339 450533
rect 287053 450530 287119 450533
rect 244273 450528 287119 450530
rect 244273 450472 244278 450528
rect 244334 450472 287058 450528
rect 287114 450472 287119 450528
rect 244273 450470 287119 450472
rect 244273 450467 244339 450470
rect 287053 450467 287119 450470
rect 193070 450332 193076 450396
rect 193140 450394 193146 450396
rect 199377 450394 199443 450397
rect 193140 450392 199443 450394
rect 193140 450336 199382 450392
rect 199438 450336 199443 450392
rect 193140 450334 199443 450336
rect 193140 450332 193146 450334
rect 199377 450331 199443 450334
rect 195237 449986 195303 449989
rect 245745 449988 245811 449989
rect 193262 449984 195303 449986
rect 193262 449928 195242 449984
rect 195298 449928 195303 449984
rect 193262 449926 195303 449928
rect 113817 449850 113883 449853
rect 116577 449850 116643 449853
rect 113817 449848 116643 449850
rect 113817 449792 113822 449848
rect 113878 449792 116582 449848
rect 116638 449792 116643 449848
rect 113817 449790 116643 449792
rect 113817 449787 113883 449790
rect 116577 449787 116643 449790
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 177798 449380 177804 449444
rect 177868 449442 177874 449444
rect 193262 449442 193322 449926
rect 195237 449923 195303 449926
rect 245694 449924 245700 449988
rect 245764 449986 245811 449988
rect 249609 449986 249675 449989
rect 267917 449986 267983 449989
rect 245764 449984 245856 449986
rect 245806 449928 245856 449984
rect 245764 449926 245856 449928
rect 249609 449984 267983 449986
rect 249609 449928 249614 449984
rect 249670 449928 267922 449984
rect 267978 449928 267983 449984
rect 249609 449926 267983 449928
rect 245764 449924 245811 449926
rect 245745 449923 245811 449924
rect 249609 449923 249675 449926
rect 267917 449923 267983 449926
rect 247033 449714 247099 449717
rect 247718 449714 247724 449716
rect 247033 449712 247724 449714
rect 247033 449656 247038 449712
rect 247094 449656 247724 449712
rect 247033 449654 247724 449656
rect 247033 449651 247099 449654
rect 247718 449652 247724 449654
rect 247788 449652 247794 449716
rect 177868 449382 193322 449442
rect 177868 449380 177874 449382
rect 190453 449170 190519 449173
rect 190453 449168 193660 449170
rect 190453 449112 190458 449168
rect 190514 449112 193660 449168
rect 190453 449110 193660 449112
rect 190453 449107 190519 449110
rect 255589 448898 255655 448901
rect 253460 448896 255655 448898
rect 253460 448840 255594 448896
rect 255650 448840 255655 448896
rect 253460 448838 255655 448840
rect 255589 448835 255655 448838
rect 253933 448764 253999 448765
rect 253933 448762 253980 448764
rect 253888 448760 253980 448762
rect 253888 448704 253938 448760
rect 253888 448702 253980 448704
rect 253933 448700 253980 448702
rect 254044 448700 254050 448764
rect 253933 448699 253999 448700
rect 70853 448628 70919 448629
rect 70853 448624 70900 448628
rect 70964 448626 70970 448628
rect 254025 448626 254091 448629
rect 254526 448626 254532 448628
rect 70853 448568 70858 448624
rect 70853 448564 70900 448568
rect 70964 448566 71010 448626
rect 254025 448624 254532 448626
rect 254025 448568 254030 448624
rect 254086 448568 254532 448624
rect 254025 448566 254532 448568
rect 70964 448564 70970 448566
rect 70853 448563 70919 448564
rect 254025 448563 254091 448566
rect 254526 448564 254532 448566
rect 254596 448564 254602 448628
rect 191782 448428 191788 448492
rect 191852 448490 191858 448492
rect 191925 448490 191991 448493
rect 191852 448488 191991 448490
rect 191852 448432 191930 448488
rect 191986 448432 191991 448488
rect 191852 448430 191991 448432
rect 191852 448428 191858 448430
rect 191925 448427 191991 448430
rect 69606 447748 69612 447812
rect 69676 447810 69682 447812
rect 191557 447810 191623 447813
rect 69676 447808 193660 447810
rect 69676 447752 191562 447808
rect 191618 447752 193660 447808
rect 69676 447750 193660 447752
rect 69676 447748 69682 447750
rect 191557 447747 191623 447750
rect 254209 447538 254275 447541
rect 254485 447538 254551 447541
rect 253460 447536 254551 447538
rect 253460 447480 254214 447536
rect 254270 447480 254490 447536
rect 254546 447480 254551 447536
rect 253460 447478 254551 447480
rect 254209 447475 254275 447478
rect 254485 447475 254551 447478
rect 253054 446796 253060 446860
rect 253124 446796 253130 446860
rect 183369 446586 183435 446589
rect 193070 446586 193076 446588
rect 183369 446584 193076 446586
rect 183369 446528 183374 446584
rect 183430 446528 193076 446584
rect 183369 446526 193076 446528
rect 183369 446523 183435 446526
rect 193070 446524 193076 446526
rect 193140 446524 193146 446588
rect 191557 446450 191623 446453
rect 253062 446450 253122 446796
rect 261109 446450 261175 446453
rect 191557 446448 193660 446450
rect 191557 446392 191562 446448
rect 191618 446392 193660 446448
rect 191557 446390 193660 446392
rect 253062 446448 261175 446450
rect 253062 446392 261114 446448
rect 261170 446392 261175 446448
rect 253062 446390 261175 446392
rect 191557 446387 191623 446390
rect 261109 446387 261175 446390
rect 255497 446178 255563 446181
rect 253460 446176 255563 446178
rect 253460 446120 255502 446176
rect 255558 446120 255563 446176
rect 253460 446118 255563 446120
rect 255497 446115 255563 446118
rect 191557 445090 191623 445093
rect 191557 445088 193660 445090
rect 191557 445032 191562 445088
rect 191618 445032 193660 445088
rect 191557 445030 193660 445032
rect 191557 445027 191623 445030
rect 255589 444818 255655 444821
rect 253460 444816 255655 444818
rect 253460 444760 255594 444816
rect 255650 444760 255655 444816
rect 253460 444758 255655 444760
rect 255589 444755 255655 444758
rect 583520 444668 584960 444908
rect 176009 444274 176075 444277
rect 176510 444274 176516 444276
rect 176009 444272 176516 444274
rect 176009 444216 176014 444272
rect 176070 444216 176516 444272
rect 176009 444214 176516 444216
rect 176009 444211 176075 444214
rect 176510 444212 176516 444214
rect 176580 444212 176586 444276
rect 193029 443730 193095 443733
rect 193029 443728 193660 443730
rect 193029 443672 193034 443728
rect 193090 443672 193660 443728
rect 193029 443670 193660 443672
rect 193029 443667 193095 443670
rect 176326 443532 176332 443596
rect 176396 443594 176402 443596
rect 191833 443594 191899 443597
rect 176396 443592 191899 443594
rect 176396 443536 191838 443592
rect 191894 443536 191899 443592
rect 176396 443534 191899 443536
rect 176396 443532 176402 443534
rect 191833 443531 191899 443534
rect 255497 443458 255563 443461
rect 253460 443456 255563 443458
rect 253460 443400 255502 443456
rect 255558 443400 255563 443456
rect 253460 443398 255563 443400
rect 255497 443395 255563 443398
rect 191373 442098 191439 442101
rect 255681 442098 255747 442101
rect 191373 442096 193660 442098
rect 191373 442040 191378 442096
rect 191434 442040 193660 442096
rect 191373 442038 193660 442040
rect 253460 442096 255747 442098
rect 253460 442040 255686 442096
rect 255742 442040 255747 442096
rect 253460 442038 255747 442040
rect 191373 442035 191439 442038
rect 255681 442035 255747 442038
rect 269757 441690 269823 441693
rect 277342 441690 277348 441692
rect 269757 441688 277348 441690
rect 269757 441632 269762 441688
rect 269818 441632 277348 441688
rect 269757 441630 277348 441632
rect 269757 441627 269823 441630
rect 277342 441628 277348 441630
rect 277412 441628 277418 441692
rect 252870 440948 252876 441012
rect 252940 440948 252946 441012
rect 50981 440874 51047 440877
rect 83733 440874 83799 440877
rect 50981 440872 83799 440874
rect 50981 440816 50986 440872
rect 51042 440816 83738 440872
rect 83794 440816 83799 440872
rect 50981 440814 83799 440816
rect 50981 440811 51047 440814
rect 83733 440811 83799 440814
rect 190637 440738 190703 440741
rect 190637 440736 193660 440738
rect 190637 440680 190642 440736
rect 190698 440680 193660 440736
rect 190637 440678 193660 440680
rect 190637 440675 190703 440678
rect 252878 440436 252938 440948
rect 63125 439514 63191 439517
rect 155677 439514 155743 439517
rect 63125 439512 155743 439514
rect 63125 439456 63130 439512
rect 63186 439456 155682 439512
rect 155738 439456 155743 439512
rect 63125 439454 155743 439456
rect 63125 439451 63191 439454
rect 155677 439451 155743 439454
rect 191649 439378 191715 439381
rect 191649 439376 193660 439378
rect 191649 439320 191654 439376
rect 191710 439320 193660 439376
rect 191649 439318 193660 439320
rect 191649 439315 191715 439318
rect 255497 439106 255563 439109
rect 253460 439104 255563 439106
rect 253460 439048 255502 439104
rect 255558 439048 255563 439104
rect 253460 439046 255563 439048
rect 255497 439043 255563 439046
rect 69657 438834 69723 438837
rect 188429 438834 188495 438837
rect 69657 438832 188495 438834
rect 69657 438776 69662 438832
rect 69718 438776 188434 438832
rect 188490 438776 188495 438832
rect 69657 438774 188495 438776
rect 69657 438771 69723 438774
rect 188429 438771 188495 438774
rect 98361 438154 98427 438157
rect 119337 438154 119403 438157
rect 98361 438152 119403 438154
rect 98361 438096 98366 438152
rect 98422 438096 119342 438152
rect 119398 438096 119403 438152
rect 98361 438094 119403 438096
rect 98361 438091 98427 438094
rect 119337 438091 119403 438094
rect 163446 438092 163452 438156
rect 163516 438154 163522 438156
rect 172513 438154 172579 438157
rect 163516 438152 172579 438154
rect 163516 438096 172518 438152
rect 172574 438096 172579 438152
rect 163516 438094 172579 438096
rect 163516 438092 163522 438094
rect 172513 438091 172579 438094
rect 190637 438018 190703 438021
rect 190637 438016 193660 438018
rect 190637 437960 190642 438016
rect 190698 437960 193660 438016
rect 190637 437958 193660 437960
rect 190637 437955 190703 437958
rect 255497 437746 255563 437749
rect 253460 437744 255563 437746
rect 253460 437688 255502 437744
rect 255558 437688 255563 437744
rect 253460 437686 255563 437688
rect 255497 437683 255563 437686
rect 255262 437548 255268 437612
rect 255332 437610 255338 437612
rect 255497 437610 255563 437613
rect 255332 437608 255563 437610
rect 255332 437552 255502 437608
rect 255558 437552 255563 437608
rect 255332 437550 255563 437552
rect 255332 437548 255338 437550
rect 255497 437547 255563 437550
rect 89345 436794 89411 436797
rect 118601 436794 118667 436797
rect 118785 436794 118851 436797
rect 89345 436792 118851 436794
rect -960 436508 480 436748
rect 89345 436736 89350 436792
rect 89406 436736 118606 436792
rect 118662 436736 118790 436792
rect 118846 436736 118851 436792
rect 89345 436734 118851 436736
rect 89345 436731 89411 436734
rect 118601 436731 118667 436734
rect 118785 436731 118851 436734
rect 153929 436794 153995 436797
rect 191557 436794 191623 436797
rect 153929 436792 191623 436794
rect 153929 436736 153934 436792
rect 153990 436736 191562 436792
rect 191618 436736 191623 436792
rect 153929 436734 191623 436736
rect 153929 436731 153995 436734
rect 191557 436731 191623 436734
rect 191649 436658 191715 436661
rect 191649 436656 193660 436658
rect 191649 436600 191654 436656
rect 191710 436600 193660 436656
rect 191649 436598 193660 436600
rect 191649 436595 191715 436598
rect 73470 436460 73476 436524
rect 73540 436522 73546 436524
rect 80329 436522 80395 436525
rect 73540 436520 80395 436522
rect 73540 436464 80334 436520
rect 80390 436464 80395 436520
rect 73540 436462 80395 436464
rect 73540 436460 73546 436462
rect 80329 436459 80395 436462
rect 79174 436324 79180 436388
rect 79244 436386 79250 436388
rect 88425 436386 88491 436389
rect 255497 436386 255563 436389
rect 79244 436384 88491 436386
rect 79244 436328 88430 436384
rect 88486 436328 88491 436384
rect 79244 436326 88491 436328
rect 253460 436384 255563 436386
rect 253460 436328 255502 436384
rect 255558 436328 255563 436384
rect 253460 436326 255563 436328
rect 79244 436324 79250 436326
rect 88425 436323 88491 436326
rect 255497 436323 255563 436326
rect 75126 436188 75132 436252
rect 75196 436250 75202 436252
rect 80053 436250 80119 436253
rect 75196 436248 80119 436250
rect 75196 436192 80058 436248
rect 80114 436192 80119 436248
rect 75196 436190 80119 436192
rect 75196 436188 75202 436190
rect 80053 436187 80119 436190
rect 81014 436188 81020 436252
rect 81084 436250 81090 436252
rect 89897 436250 89963 436253
rect 81084 436248 89963 436250
rect 81084 436192 89902 436248
rect 89958 436192 89963 436248
rect 81084 436190 89963 436192
rect 81084 436188 81090 436190
rect 89897 436187 89963 436190
rect 71078 436052 71084 436116
rect 71148 436114 71154 436116
rect 75453 436114 75519 436117
rect 71148 436112 75519 436114
rect 71148 436056 75458 436112
rect 75514 436056 75519 436112
rect 71148 436054 75519 436056
rect 71148 436052 71154 436054
rect 75453 436051 75519 436054
rect 94446 436052 94452 436116
rect 94516 436114 94522 436116
rect 96705 436114 96771 436117
rect 96981 436114 97047 436117
rect 94516 436112 97047 436114
rect 94516 436056 96710 436112
rect 96766 436056 96986 436112
rect 97042 436056 97047 436112
rect 94516 436054 97047 436056
rect 94516 436052 94522 436054
rect 96705 436051 96771 436054
rect 96981 436051 97047 436054
rect 106038 436052 106044 436116
rect 106108 436114 106114 436116
rect 107653 436114 107719 436117
rect 106108 436112 107719 436114
rect 106108 436056 107658 436112
rect 107714 436056 107719 436112
rect 106108 436054 107719 436056
rect 106108 436052 106114 436054
rect 107653 436051 107719 436054
rect 66069 435298 66135 435301
rect 178033 435298 178099 435301
rect 66069 435296 178099 435298
rect 66069 435240 66074 435296
rect 66130 435240 178038 435296
rect 178094 435240 178099 435296
rect 66069 435238 178099 435240
rect 66069 435235 66135 435238
rect 178033 435235 178099 435238
rect 191557 435298 191623 435301
rect 191557 435296 193660 435298
rect 191557 435240 191562 435296
rect 191618 435240 193660 435296
rect 191557 435238 193660 435240
rect 191557 435235 191623 435238
rect 255497 435026 255563 435029
rect 253460 435024 255563 435026
rect 253460 434968 255502 435024
rect 255558 434968 255563 435024
rect 253460 434966 255563 434968
rect 255497 434963 255563 434966
rect 52269 434754 52335 434757
rect 68369 434754 68435 434757
rect 52269 434752 68435 434754
rect 52269 434696 52274 434752
rect 52330 434696 68374 434752
rect 68430 434696 68435 434752
rect 52269 434694 68435 434696
rect 52269 434691 52335 434694
rect 68369 434691 68435 434694
rect 102726 434556 102732 434620
rect 102796 434618 102802 434620
rect 104893 434618 104959 434621
rect 102796 434616 104959 434618
rect 102796 434560 104898 434616
rect 104954 434560 104959 434616
rect 102796 434558 104959 434560
rect 102796 434556 102802 434558
rect 104893 434555 104959 434558
rect 69289 434348 69355 434349
rect 69238 434346 69244 434348
rect 69198 434286 69244 434346
rect 69308 434344 69355 434348
rect 69350 434288 69355 434344
rect 69238 434284 69244 434286
rect 69308 434284 69355 434288
rect 95182 434284 95188 434348
rect 95252 434346 95258 434348
rect 95693 434346 95759 434349
rect 100201 434348 100267 434349
rect 100150 434346 100156 434348
rect 95252 434344 95759 434346
rect 95252 434288 95698 434344
rect 95754 434288 95759 434344
rect 95252 434286 95759 434288
rect 100110 434286 100156 434346
rect 100220 434344 100267 434348
rect 100262 434288 100267 434344
rect 95252 434284 95258 434286
rect 69289 434283 69355 434284
rect 95693 434283 95759 434286
rect 100150 434284 100156 434286
rect 100220 434284 100267 434288
rect 100201 434283 100267 434284
rect 92749 434212 92815 434213
rect 92749 434208 92796 434212
rect 92860 434210 92866 434212
rect 92749 434152 92754 434208
rect 92749 434148 92796 434152
rect 92860 434150 92906 434210
rect 92860 434148 92866 434150
rect 92749 434147 92815 434148
rect 80646 434012 80652 434076
rect 80716 434074 80722 434076
rect 80973 434074 81039 434077
rect 80716 434072 81039 434074
rect 80716 434016 80978 434072
rect 81034 434016 81039 434072
rect 80716 434014 81039 434016
rect 80716 434012 80722 434014
rect 80973 434011 81039 434014
rect 67950 433876 67956 433940
rect 68020 433938 68026 433940
rect 191465 433938 191531 433941
rect 68020 433936 193690 433938
rect 68020 433880 191470 433936
rect 191526 433880 193690 433936
rect 68020 433878 193690 433880
rect 68020 433876 68026 433878
rect 191465 433875 191531 433878
rect 77477 433802 77543 433805
rect 78213 433802 78279 433805
rect 78438 433802 78444 433804
rect 77477 433800 78444 433802
rect 77477 433744 77482 433800
rect 77538 433744 78218 433800
rect 78274 433744 78444 433800
rect 77477 433742 78444 433744
rect 77477 433739 77543 433742
rect 78213 433739 78279 433742
rect 78438 433740 78444 433742
rect 78508 433740 78514 433804
rect 85849 433802 85915 433805
rect 86718 433802 86724 433804
rect 85849 433800 86724 433802
rect 85849 433744 85854 433800
rect 85910 433744 86724 433800
rect 85849 433742 86724 433744
rect 85849 433739 85915 433742
rect 86718 433740 86724 433742
rect 86788 433740 86794 433804
rect 98494 433740 98500 433804
rect 98564 433802 98570 433804
rect 101213 433802 101279 433805
rect 98564 433800 101279 433802
rect 98564 433744 101218 433800
rect 101274 433744 101279 433800
rect 98564 433742 101279 433744
rect 98564 433740 98570 433742
rect 101213 433739 101279 433742
rect 74809 433668 74875 433669
rect 74758 433604 74764 433668
rect 74828 433666 74875 433668
rect 74828 433664 74920 433666
rect 74870 433608 74920 433664
rect 74828 433606 74920 433608
rect 74828 433604 74875 433606
rect 75862 433604 75868 433668
rect 75932 433666 75938 433668
rect 76189 433666 76255 433669
rect 75932 433664 76255 433666
rect 75932 433608 76194 433664
rect 76250 433608 76255 433664
rect 75932 433606 76255 433608
rect 75932 433604 75938 433606
rect 74809 433603 74875 433604
rect 76189 433603 76255 433606
rect 78121 433666 78187 433669
rect 81893 433668 81959 433669
rect 78254 433666 78260 433668
rect 78121 433664 78260 433666
rect 78121 433608 78126 433664
rect 78182 433608 78260 433664
rect 78121 433606 78260 433608
rect 78121 433603 78187 433606
rect 78254 433604 78260 433606
rect 78324 433604 78330 433668
rect 81893 433666 81940 433668
rect 81848 433664 81940 433666
rect 81848 433608 81898 433664
rect 81848 433606 81940 433608
rect 81893 433604 81940 433606
rect 82004 433604 82010 433668
rect 82486 433604 82492 433668
rect 82556 433666 82562 433668
rect 82905 433666 82971 433669
rect 82556 433664 82971 433666
rect 82556 433608 82910 433664
rect 82966 433608 82971 433664
rect 82556 433606 82971 433608
rect 82556 433604 82562 433606
rect 81893 433603 81959 433604
rect 82905 433603 82971 433606
rect 83038 433604 83044 433668
rect 83108 433666 83114 433668
rect 83825 433666 83891 433669
rect 84561 433668 84627 433669
rect 83108 433664 83891 433666
rect 83108 433608 83830 433664
rect 83886 433608 83891 433664
rect 83108 433606 83891 433608
rect 83108 433604 83114 433606
rect 83825 433603 83891 433606
rect 84510 433604 84516 433668
rect 84580 433666 84627 433668
rect 84580 433664 84672 433666
rect 84622 433608 84672 433664
rect 84580 433606 84672 433608
rect 84580 433604 84627 433606
rect 85798 433604 85804 433668
rect 85868 433666 85874 433668
rect 85941 433666 86007 433669
rect 85868 433664 86007 433666
rect 85868 433608 85946 433664
rect 86002 433608 86007 433664
rect 85868 433606 86007 433608
rect 85868 433604 85874 433606
rect 84561 433603 84627 433604
rect 85941 433603 86007 433606
rect 87086 433604 87092 433668
rect 87156 433666 87162 433668
rect 87229 433666 87295 433669
rect 87156 433664 87295 433666
rect 87156 433608 87234 433664
rect 87290 433608 87295 433664
rect 87156 433606 87295 433608
rect 87156 433604 87162 433606
rect 87229 433603 87295 433606
rect 89662 433604 89668 433668
rect 89732 433666 89738 433668
rect 89989 433666 90055 433669
rect 89732 433664 90055 433666
rect 89732 433608 89994 433664
rect 90050 433608 90055 433664
rect 89732 433606 90055 433608
rect 89732 433604 89738 433606
rect 89989 433603 90055 433606
rect 90214 433604 90220 433668
rect 90284 433666 90290 433668
rect 90725 433666 90791 433669
rect 91553 433668 91619 433669
rect 93025 433668 93091 433669
rect 91502 433666 91508 433668
rect 90284 433664 90791 433666
rect 90284 433608 90730 433664
rect 90786 433608 90791 433664
rect 90284 433606 90791 433608
rect 91462 433606 91508 433666
rect 91572 433664 91619 433668
rect 92974 433666 92980 433668
rect 91614 433608 91619 433664
rect 90284 433604 90290 433606
rect 90725 433603 90791 433606
rect 91502 433604 91508 433606
rect 91572 433604 91619 433608
rect 92934 433606 92980 433666
rect 93044 433664 93091 433668
rect 93086 433608 93091 433664
rect 92974 433604 92980 433606
rect 93044 433604 93091 433608
rect 97942 433604 97948 433668
rect 98012 433666 98018 433668
rect 98453 433666 98519 433669
rect 98012 433664 98519 433666
rect 98012 433608 98458 433664
rect 98514 433608 98519 433664
rect 98012 433606 98519 433608
rect 98012 433604 98018 433606
rect 91553 433603 91619 433604
rect 93025 433603 93091 433604
rect 98453 433603 98519 433606
rect 99833 433666 99899 433669
rect 100661 433668 100727 433669
rect 99966 433666 99972 433668
rect 99833 433664 99972 433666
rect 99833 433608 99838 433664
rect 99894 433608 99972 433664
rect 99833 433606 99972 433608
rect 99833 433603 99899 433606
rect 99966 433604 99972 433606
rect 100036 433604 100042 433668
rect 100661 433664 100708 433668
rect 100772 433666 100778 433668
rect 100661 433608 100666 433664
rect 100661 433604 100708 433608
rect 100772 433606 100818 433666
rect 100772 433604 100778 433606
rect 106406 433604 106412 433668
rect 106476 433666 106482 433668
rect 106733 433666 106799 433669
rect 106476 433664 106799 433666
rect 106476 433608 106738 433664
rect 106794 433608 106799 433664
rect 106476 433606 106799 433608
rect 106476 433604 106482 433606
rect 100661 433603 100727 433604
rect 106733 433603 106799 433606
rect 109493 433668 109559 433669
rect 109493 433664 109540 433668
rect 109604 433666 109610 433668
rect 109493 433608 109498 433664
rect 109493 433604 109540 433608
rect 109604 433606 109650 433666
rect 109604 433604 109610 433606
rect 111006 433604 111012 433668
rect 111076 433666 111082 433668
rect 111701 433666 111767 433669
rect 111076 433664 111767 433666
rect 111076 433608 111706 433664
rect 111762 433608 111767 433664
rect 193630 433636 193690 433878
rect 255497 433666 255563 433669
rect 253460 433664 255563 433666
rect 111076 433606 111767 433608
rect 253460 433608 255502 433664
rect 255558 433608 255563 433664
rect 253460 433606 255563 433608
rect 111076 433604 111082 433606
rect 109493 433603 109559 433604
rect 111701 433603 111767 433606
rect 255497 433603 255563 433606
rect 66805 433394 66871 433397
rect 115749 433394 115815 433397
rect 66805 433392 68908 433394
rect 66805 433336 66810 433392
rect 66866 433336 68908 433392
rect 66805 433334 68908 433336
rect 112700 433392 115815 433394
rect 112700 433336 115754 433392
rect 115810 433336 115815 433392
rect 112700 433334 115815 433336
rect 66805 433331 66871 433334
rect 115749 433331 115815 433334
rect 143257 433258 143323 433261
rect 148174 433258 148180 433260
rect 143257 433256 148180 433258
rect 143257 433200 143262 433256
rect 143318 433200 148180 433256
rect 143257 433198 148180 433200
rect 143257 433195 143323 433198
rect 148174 433196 148180 433198
rect 148244 433196 148250 433260
rect 69422 433060 69428 433124
rect 69492 433060 69498 433124
rect 65977 432578 66043 432581
rect 69430 432578 69490 433060
rect 65977 432576 69490 432578
rect 65977 432520 65982 432576
rect 66038 432548 69490 432576
rect 66038 432520 69460 432548
rect 65977 432518 69460 432520
rect 65977 432515 66043 432518
rect 115841 432306 115907 432309
rect 112700 432304 115907 432306
rect 112700 432248 115846 432304
rect 115902 432248 115907 432304
rect 112700 432246 115907 432248
rect 115841 432243 115907 432246
rect 191649 432306 191715 432309
rect 191649 432304 193660 432306
rect 191649 432248 191654 432304
rect 191710 432248 193660 432304
rect 191649 432246 193660 432248
rect 191649 432243 191715 432246
rect 255957 432034 256023 432037
rect 253460 432032 256023 432034
rect 253460 431976 255962 432032
rect 256018 431976 256023 432032
rect 253460 431974 256023 431976
rect 255957 431971 256023 431974
rect 582741 431626 582807 431629
rect 583520 431626 584960 431716
rect 582741 431624 584960 431626
rect 582741 431568 582746 431624
rect 582802 431568 584960 431624
rect 582741 431566 584960 431568
rect 582741 431563 582807 431566
rect 67541 431490 67607 431493
rect 67541 431488 68908 431490
rect 67541 431432 67546 431488
rect 67602 431432 68908 431488
rect 583520 431476 584960 431566
rect 67541 431430 68908 431432
rect 67541 431427 67607 431430
rect 115565 431218 115631 431221
rect 112700 431216 115631 431218
rect 112700 431160 115570 431216
rect 115626 431160 115631 431216
rect 112700 431158 115631 431160
rect 115565 431155 115631 431158
rect 191741 430946 191807 430949
rect 191741 430944 193660 430946
rect 191741 430888 191746 430944
rect 191802 430888 193660 430944
rect 191741 430886 193660 430888
rect 191741 430883 191807 430886
rect 253054 430884 253060 430948
rect 253124 430946 253130 430948
rect 253974 430946 253980 430948
rect 253124 430886 253980 430946
rect 253124 430884 253130 430886
rect 253974 430884 253980 430886
rect 254044 430884 254050 430948
rect 255405 430674 255471 430677
rect 253460 430672 255471 430674
rect 253460 430616 255410 430672
rect 255466 430616 255471 430672
rect 253460 430614 255471 430616
rect 255405 430611 255471 430614
rect 66161 430402 66227 430405
rect 66161 430400 68908 430402
rect 66161 430344 66166 430400
rect 66222 430344 68908 430400
rect 66161 430342 68908 430344
rect 66161 430339 66227 430342
rect 114829 430130 114895 430133
rect 112700 430128 114895 430130
rect 112700 430072 114834 430128
rect 114890 430072 114895 430128
rect 112700 430070 114895 430072
rect 114829 430067 114895 430070
rect 253565 429858 253631 429861
rect 253430 429856 253631 429858
rect 253430 429800 253570 429856
rect 253626 429800 253631 429856
rect 253430 429798 253631 429800
rect 191005 429586 191071 429589
rect 191005 429584 193660 429586
rect 191005 429528 191010 429584
rect 191066 429528 193660 429584
rect 191005 429526 193660 429528
rect 191005 429523 191071 429526
rect 66621 429314 66687 429317
rect 115749 429314 115815 429317
rect 66621 429312 68908 429314
rect 66621 429256 66626 429312
rect 66682 429256 68908 429312
rect 66621 429254 68908 429256
rect 112700 429312 115815 429314
rect 112700 429256 115754 429312
rect 115810 429256 115815 429312
rect 112700 429254 115815 429256
rect 66621 429251 66687 429254
rect 115749 429251 115815 429254
rect 143349 429314 143415 429317
rect 148174 429314 148180 429316
rect 143349 429312 148180 429314
rect 143349 429256 143354 429312
rect 143410 429256 148180 429312
rect 143349 429254 148180 429256
rect 143349 429251 143415 429254
rect 148174 429252 148180 429254
rect 148244 429252 148250 429316
rect 253430 429284 253490 429798
rect 253565 429795 253631 429798
rect 67725 428226 67791 428229
rect 113214 428226 113220 428228
rect 67725 428224 68908 428226
rect 67725 428168 67730 428224
rect 67786 428168 68908 428224
rect 67725 428166 68908 428168
rect 112700 428166 113220 428226
rect 67725 428163 67791 428166
rect 113214 428164 113220 428166
rect 113284 428226 113290 428228
rect 115841 428226 115907 428229
rect 113284 428224 115907 428226
rect 113284 428168 115846 428224
rect 115902 428168 115907 428224
rect 113284 428166 115907 428168
rect 113284 428164 113290 428166
rect 115841 428163 115907 428166
rect 190821 428226 190887 428229
rect 190821 428224 193660 428226
rect 190821 428168 190826 428224
rect 190882 428168 193660 428224
rect 190821 428166 193660 428168
rect 190821 428163 190887 428166
rect 254209 427954 254275 427957
rect 253460 427952 254275 427954
rect 253460 427896 254214 427952
rect 254270 427896 254275 427952
rect 253460 427894 254275 427896
rect 254209 427891 254275 427894
rect 66805 427410 66871 427413
rect 66805 427408 68908 427410
rect 66805 427352 66810 427408
rect 66866 427352 68908 427408
rect 66805 427350 68908 427352
rect 66805 427347 66871 427350
rect 114502 427138 114508 427140
rect 112700 427078 114508 427138
rect 114502 427076 114508 427078
rect 114572 427076 114578 427140
rect 170806 427076 170812 427140
rect 170876 427138 170882 427140
rect 177297 427138 177363 427141
rect 170876 427136 177363 427138
rect 170876 427080 177302 427136
rect 177358 427080 177363 427136
rect 170876 427078 177363 427080
rect 170876 427076 170882 427078
rect 177297 427075 177363 427078
rect 190821 426866 190887 426869
rect 190821 426864 193660 426866
rect 190821 426808 190826 426864
rect 190882 426808 193660 426864
rect 190821 426806 193660 426808
rect 190821 426803 190887 426806
rect 255405 426594 255471 426597
rect 253460 426592 255471 426594
rect 253460 426536 255410 426592
rect 255466 426536 255471 426592
rect 253460 426534 255471 426536
rect 255405 426531 255471 426534
rect 68878 425642 68938 426292
rect 113265 426050 113331 426053
rect 115841 426050 115907 426053
rect 112700 426048 115907 426050
rect 112700 425992 113270 426048
rect 113326 425992 115846 426048
rect 115902 425992 115907 426048
rect 112700 425990 115907 425992
rect 113265 425987 113331 425990
rect 115841 425987 115907 425990
rect 64830 425582 68938 425642
rect 56501 425098 56567 425101
rect 63125 425098 63191 425101
rect 64830 425098 64890 425582
rect 191741 425506 191807 425509
rect 191741 425504 193660 425506
rect 191741 425448 191746 425504
rect 191802 425448 193660 425504
rect 191741 425446 193660 425448
rect 191741 425443 191807 425446
rect 66621 425234 66687 425237
rect 255497 425234 255563 425237
rect 66621 425232 68908 425234
rect 66621 425176 66626 425232
rect 66682 425176 68908 425232
rect 66621 425174 68908 425176
rect 253460 425232 255563 425234
rect 253460 425176 255502 425232
rect 255558 425176 255563 425232
rect 253460 425174 255563 425176
rect 66621 425171 66687 425174
rect 255497 425171 255563 425174
rect 56501 425096 64890 425098
rect 56501 425040 56506 425096
rect 56562 425040 63130 425096
rect 63186 425040 64890 425096
rect 56501 425038 64890 425040
rect 56501 425035 56567 425038
rect 63125 425035 63191 425038
rect 113817 424962 113883 424965
rect 112700 424960 113883 424962
rect 112700 424904 113822 424960
rect 113878 424904 113883 424960
rect 112700 424902 113883 424904
rect 113817 424899 113883 424902
rect 66805 424146 66871 424149
rect 115841 424146 115907 424149
rect 66805 424144 68908 424146
rect 66805 424088 66810 424144
rect 66866 424088 68908 424144
rect 66805 424086 68908 424088
rect 112700 424144 115907 424146
rect 112700 424088 115846 424144
rect 115902 424088 115907 424144
rect 112700 424086 115907 424088
rect 66805 424083 66871 424086
rect 115841 424083 115907 424086
rect 191741 423874 191807 423877
rect 191741 423872 193660 423874
rect 191741 423816 191746 423872
rect 191802 423816 193660 423872
rect 191741 423814 193660 423816
rect 191741 423811 191807 423814
rect 168189 423738 168255 423741
rect 172094 423738 172100 423740
rect 168189 423736 172100 423738
rect -960 423602 480 423692
rect 168189 423680 168194 423736
rect 168250 423680 172100 423736
rect 168189 423678 172100 423680
rect 168189 423675 168255 423678
rect 172094 423676 172100 423678
rect 172164 423676 172170 423740
rect 3417 423602 3483 423605
rect 255497 423602 255563 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect 253460 423600 255563 423602
rect 253460 423544 255502 423600
rect 255558 423544 255563 423600
rect 253460 423542 255563 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 255497 423539 255563 423542
rect 66110 423268 66116 423332
rect 66180 423330 66186 423332
rect 66253 423330 66319 423333
rect 66180 423328 68908 423330
rect 66180 423272 66258 423328
rect 66314 423272 68908 423328
rect 66180 423270 68908 423272
rect 66180 423268 66186 423270
rect 66253 423267 66319 423270
rect 115841 423058 115907 423061
rect 112700 423056 115907 423058
rect 112700 423000 115846 423056
rect 115902 423000 115907 423056
rect 112700 422998 115907 423000
rect 115841 422995 115907 422998
rect 191005 422514 191071 422517
rect 191005 422512 193660 422514
rect 191005 422456 191010 422512
rect 191066 422456 193660 422512
rect 191005 422454 193660 422456
rect 191005 422451 191071 422454
rect 67173 422242 67239 422245
rect 67950 422242 67956 422244
rect 67173 422240 67956 422242
rect 67173 422184 67178 422240
rect 67234 422184 67956 422240
rect 67173 422182 67956 422184
rect 67173 422179 67239 422182
rect 67950 422180 67956 422182
rect 68020 422242 68026 422244
rect 255497 422242 255563 422245
rect 68020 422182 68908 422242
rect 253460 422240 255563 422242
rect 253460 422184 255502 422240
rect 255558 422184 255563 422240
rect 253460 422182 255563 422184
rect 68020 422180 68026 422182
rect 255497 422179 255563 422182
rect 115197 421970 115263 421973
rect 112700 421968 115263 421970
rect 112700 421912 115202 421968
rect 115258 421912 115263 421968
rect 112700 421910 115263 421912
rect 115197 421907 115263 421910
rect 66897 421154 66963 421157
rect 191741 421154 191807 421157
rect 66897 421152 68908 421154
rect 66897 421096 66902 421152
rect 66958 421096 68908 421152
rect 66897 421094 68908 421096
rect 191741 421152 193660 421154
rect 191741 421096 191746 421152
rect 191802 421096 193660 421152
rect 191741 421094 193660 421096
rect 66897 421091 66963 421094
rect 191741 421091 191807 421094
rect 113173 420882 113239 420885
rect 255497 420882 255563 420885
rect 112700 420880 113239 420882
rect 112700 420824 113178 420880
rect 113234 420824 113239 420880
rect 112700 420822 113239 420824
rect 253460 420880 255563 420882
rect 253460 420824 255502 420880
rect 255558 420824 255563 420880
rect 253460 420822 255563 420824
rect 113173 420819 113239 420822
rect 255497 420819 255563 420822
rect 67357 420066 67423 420069
rect 114645 420066 114711 420069
rect 67357 420064 68908 420066
rect 67357 420008 67362 420064
rect 67418 420008 68908 420064
rect 67357 420006 68908 420008
rect 112700 420064 114711 420066
rect 112700 420008 114650 420064
rect 114706 420008 114711 420064
rect 112700 420006 114711 420008
rect 67357 420003 67423 420006
rect 114645 420003 114711 420006
rect 192477 419794 192543 419797
rect 192477 419792 193660 419794
rect 192477 419736 192482 419792
rect 192538 419736 193660 419792
rect 192477 419734 193660 419736
rect 192477 419731 192543 419734
rect 155585 419658 155651 419661
rect 155718 419658 155724 419660
rect 155585 419656 155724 419658
rect 155585 419600 155590 419656
rect 155646 419600 155724 419656
rect 155585 419598 155724 419600
rect 155585 419595 155651 419598
rect 155718 419596 155724 419598
rect 155788 419596 155794 419660
rect 172278 419596 172284 419660
rect 172348 419658 172354 419660
rect 177573 419658 177639 419661
rect 172348 419656 177639 419658
rect 172348 419600 177578 419656
rect 177634 419600 177639 419656
rect 172348 419598 177639 419600
rect 172348 419596 172354 419598
rect 177573 419595 177639 419598
rect 255405 419522 255471 419525
rect 253460 419520 255471 419522
rect 253460 419464 255410 419520
rect 255466 419464 255471 419520
rect 253460 419462 255471 419464
rect 255405 419459 255471 419462
rect 66621 418978 66687 418981
rect 113357 418978 113423 418981
rect 115841 418978 115907 418981
rect 66621 418976 68908 418978
rect 66621 418920 66626 418976
rect 66682 418920 68908 418976
rect 66621 418918 68908 418920
rect 112700 418976 115907 418978
rect 112700 418920 113362 418976
rect 113418 418920 115846 418976
rect 115902 418920 115907 418976
rect 112700 418918 115907 418920
rect 66621 418915 66687 418918
rect 113357 418915 113423 418918
rect 115841 418915 115907 418918
rect 191741 418434 191807 418437
rect 191741 418432 193660 418434
rect 191741 418376 191746 418432
rect 191802 418376 193660 418432
rect 191741 418374 193660 418376
rect 191741 418371 191807 418374
rect 287094 418236 287100 418300
rect 287164 418298 287170 418300
rect 287421 418298 287487 418301
rect 287164 418296 287487 418298
rect 287164 418240 287426 418296
rect 287482 418240 287487 418296
rect 287164 418238 287487 418240
rect 287164 418236 287170 418238
rect 287421 418235 287487 418238
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 66989 418162 67055 418165
rect 255405 418162 255471 418165
rect 66989 418160 68908 418162
rect 66989 418104 66994 418160
rect 67050 418104 68908 418160
rect 66989 418102 68908 418104
rect 253460 418160 255471 418162
rect 253460 418104 255410 418160
rect 255466 418104 255471 418160
rect 583520 418148 584960 418238
rect 253460 418102 255471 418104
rect 66989 418099 67055 418102
rect 255405 418099 255471 418102
rect 114553 417890 114619 417893
rect 112700 417888 114619 417890
rect 112700 417832 114558 417888
rect 114614 417832 114619 417888
rect 112700 417830 114619 417832
rect 114553 417827 114619 417830
rect 154389 417482 154455 417485
rect 188286 417482 188292 417484
rect 154389 417480 188292 417482
rect 154389 417424 154394 417480
rect 154450 417424 188292 417480
rect 154389 417422 188292 417424
rect 154389 417419 154455 417422
rect 188286 417420 188292 417422
rect 188356 417420 188362 417484
rect 67449 417074 67515 417077
rect 191741 417074 191807 417077
rect 67449 417072 68908 417074
rect 67449 417016 67454 417072
rect 67510 417016 68908 417072
rect 67449 417014 68908 417016
rect 191741 417072 193660 417074
rect 191741 417016 191746 417072
rect 191802 417016 193660 417072
rect 191741 417014 193660 417016
rect 67449 417011 67515 417014
rect 191741 417011 191807 417014
rect 115841 416802 115907 416805
rect 255405 416802 255471 416805
rect 112700 416800 115907 416802
rect 112700 416744 115846 416800
rect 115902 416744 115907 416800
rect 112700 416742 115907 416744
rect 253460 416800 255471 416802
rect 253460 416744 255410 416800
rect 255466 416744 255471 416800
rect 253460 416742 255471 416744
rect 115841 416739 115907 416742
rect 255405 416739 255471 416742
rect 280286 416740 280292 416804
rect 280356 416802 280362 416804
rect 280429 416802 280495 416805
rect 280356 416800 280495 416802
rect 280356 416744 280434 416800
rect 280490 416744 280495 416800
rect 280356 416742 280495 416744
rect 280356 416740 280362 416742
rect 280429 416739 280495 416742
rect 66805 415986 66871 415989
rect 66805 415984 68908 415986
rect 66805 415928 66810 415984
rect 66866 415928 68908 415984
rect 66805 415926 68908 415928
rect 66805 415923 66871 415926
rect 115841 415714 115907 415717
rect 112700 415712 115907 415714
rect 112700 415656 115846 415712
rect 115902 415656 115907 415712
rect 112700 415654 115907 415656
rect 115841 415651 115907 415654
rect 190637 415442 190703 415445
rect 190637 415440 193660 415442
rect 190637 415384 190642 415440
rect 190698 415384 193660 415440
rect 190637 415382 193660 415384
rect 190637 415379 190703 415382
rect 254526 415170 254532 415172
rect 253460 415110 254532 415170
rect 254526 415108 254532 415110
rect 254596 415170 254602 415172
rect 255313 415170 255379 415173
rect 254596 415168 255379 415170
rect 254596 415112 255318 415168
rect 255374 415112 255379 415168
rect 254596 415110 255379 415112
rect 254596 415108 254602 415110
rect 255313 415107 255379 415110
rect 66805 414898 66871 414901
rect 115841 414898 115907 414901
rect 66805 414896 68908 414898
rect 66805 414840 66810 414896
rect 66866 414840 68908 414896
rect 66805 414838 68908 414840
rect 112700 414896 115907 414898
rect 112700 414840 115846 414896
rect 115902 414840 115907 414896
rect 112700 414838 115907 414840
rect 66805 414835 66871 414838
rect 115841 414835 115907 414838
rect 65885 414082 65951 414085
rect 191465 414082 191531 414085
rect 65885 414080 68908 414082
rect 65885 414024 65890 414080
rect 65946 414024 68908 414080
rect 65885 414022 68908 414024
rect 191465 414080 193660 414082
rect 191465 414024 191470 414080
rect 191526 414024 193660 414080
rect 191465 414022 193660 414024
rect 65885 414019 65951 414022
rect 191465 414019 191531 414022
rect 114737 413946 114803 413949
rect 113130 413944 114803 413946
rect 113130 413888 114742 413944
rect 114798 413888 114803 413944
rect 113130 413886 114803 413888
rect 113130 413810 113190 413886
rect 114737 413883 114803 413886
rect 144637 413946 144703 413949
rect 150934 413946 150940 413948
rect 144637 413944 150940 413946
rect 144637 413888 144642 413944
rect 144698 413888 150940 413944
rect 144637 413886 150940 413888
rect 144637 413883 144703 413886
rect 150934 413884 150940 413886
rect 151004 413884 151010 413948
rect 255405 413810 255471 413813
rect 112700 413750 113190 413810
rect 253460 413808 255471 413810
rect 253460 413752 255410 413808
rect 255466 413752 255471 413808
rect 253460 413750 255471 413752
rect 255405 413747 255471 413750
rect 66621 412994 66687 412997
rect 66621 412992 68908 412994
rect 66621 412936 66626 412992
rect 66682 412936 68908 412992
rect 66621 412934 68908 412936
rect 66621 412931 66687 412934
rect 115749 412722 115815 412725
rect 112700 412720 115815 412722
rect 112700 412664 115754 412720
rect 115810 412664 115815 412720
rect 112700 412662 115815 412664
rect 115749 412659 115815 412662
rect 191741 412722 191807 412725
rect 191741 412720 193660 412722
rect 191741 412664 191746 412720
rect 191802 412664 193660 412720
rect 191741 412662 193660 412664
rect 191741 412659 191807 412662
rect 255405 412450 255471 412453
rect 253460 412448 255471 412450
rect 253460 412392 255410 412448
rect 255466 412392 255471 412448
rect 253460 412390 255471 412392
rect 255405 412387 255471 412390
rect 66897 411906 66963 411909
rect 66897 411904 68908 411906
rect 66897 411848 66902 411904
rect 66958 411848 68908 411904
rect 66897 411846 68908 411848
rect 66897 411843 66963 411846
rect 115013 411634 115079 411637
rect 112700 411632 115079 411634
rect 112700 411576 115018 411632
rect 115074 411576 115079 411632
rect 112700 411574 115079 411576
rect 115013 411571 115079 411574
rect 192845 411362 192911 411365
rect 193121 411362 193187 411365
rect 192845 411360 193660 411362
rect 192845 411304 192850 411360
rect 192906 411304 193126 411360
rect 193182 411304 193660 411360
rect 192845 411302 193660 411304
rect 192845 411299 192911 411302
rect 193121 411299 193187 411302
rect 255497 411090 255563 411093
rect 253460 411088 255563 411090
rect 253460 411032 255502 411088
rect 255558 411032 255563 411088
rect 253460 411030 255563 411032
rect 255497 411027 255563 411030
rect 66805 410818 66871 410821
rect 66805 410816 68908 410818
rect 66805 410760 66810 410816
rect 66866 410760 68908 410816
rect 66805 410758 68908 410760
rect 66805 410755 66871 410758
rect -960 410546 480 410636
rect 2773 410546 2839 410549
rect 115565 410546 115631 410549
rect -960 410544 2839 410546
rect -960 410488 2778 410544
rect 2834 410488 2839 410544
rect -960 410486 2839 410488
rect 112700 410544 115631 410546
rect 112700 410488 115570 410544
rect 115626 410488 115631 410544
rect 112700 410486 115631 410488
rect -960 410396 480 410486
rect 2773 410483 2839 410486
rect 115565 410483 115631 410486
rect 190453 410002 190519 410005
rect 190453 410000 193660 410002
rect 190453 409944 190458 410000
rect 190514 409944 193660 410000
rect 190453 409942 193660 409944
rect 190453 409939 190519 409942
rect 67633 409730 67699 409733
rect 115841 409730 115907 409733
rect 255405 409730 255471 409733
rect 67633 409728 68908 409730
rect 67633 409672 67638 409728
rect 67694 409672 68908 409728
rect 67633 409670 68908 409672
rect 112700 409728 115907 409730
rect 112700 409672 115846 409728
rect 115902 409672 115907 409728
rect 112700 409670 115907 409672
rect 253460 409728 255471 409730
rect 253460 409672 255410 409728
rect 255466 409672 255471 409728
rect 253460 409670 255471 409672
rect 67633 409667 67699 409670
rect 115841 409667 115907 409670
rect 255405 409667 255471 409670
rect 123569 409186 123635 409189
rect 151721 409186 151787 409189
rect 188429 409186 188495 409189
rect 123569 409184 188495 409186
rect 123569 409128 123574 409184
rect 123630 409128 151726 409184
rect 151782 409128 188434 409184
rect 188490 409128 188495 409184
rect 123569 409126 188495 409128
rect 123569 409123 123635 409126
rect 151721 409123 151787 409126
rect 188429 409123 188495 409126
rect 66805 408914 66871 408917
rect 66805 408912 68908 408914
rect 66805 408856 66810 408912
rect 66866 408856 68908 408912
rect 66805 408854 68908 408856
rect 66805 408851 66871 408854
rect 115841 408642 115907 408645
rect 112700 408640 115907 408642
rect 112700 408584 115846 408640
rect 115902 408584 115907 408640
rect 112700 408582 115907 408584
rect 115841 408579 115907 408582
rect 191741 408642 191807 408645
rect 191741 408640 193660 408642
rect 191741 408584 191746 408640
rect 191802 408584 193660 408640
rect 191741 408582 193660 408584
rect 191741 408579 191807 408582
rect 255405 408370 255471 408373
rect 253460 408368 255471 408370
rect 253460 408312 255410 408368
rect 255466 408312 255471 408368
rect 253460 408310 255471 408312
rect 255405 408307 255471 408310
rect 66897 407826 66963 407829
rect 66897 407824 68908 407826
rect 66897 407768 66902 407824
rect 66958 407768 68908 407824
rect 66897 407766 68908 407768
rect 66897 407763 66963 407766
rect 112670 407146 112730 407524
rect 113081 407146 113147 407149
rect 112670 407144 113147 407146
rect 112670 407088 113086 407144
rect 113142 407088 113147 407144
rect 112670 407086 113147 407088
rect 113081 407083 113147 407086
rect 191741 407010 191807 407013
rect 255497 407010 255563 407013
rect 191741 407008 193660 407010
rect 191741 406952 191746 407008
rect 191802 406952 193660 407008
rect 191741 406950 193660 406952
rect 253460 407008 255563 407010
rect 253460 406952 255502 407008
rect 255558 406952 255563 407008
rect 253460 406950 255563 406952
rect 191741 406947 191807 406950
rect 255497 406947 255563 406950
rect 66805 406738 66871 406741
rect 66805 406736 68908 406738
rect 66805 406680 66810 406736
rect 66866 406680 68908 406736
rect 66805 406678 68908 406680
rect 66805 406675 66871 406678
rect 114461 406466 114527 406469
rect 115197 406466 115263 406469
rect 112700 406464 115263 406466
rect 112700 406408 114466 406464
rect 114522 406408 115202 406464
rect 115258 406408 115263 406464
rect 112700 406406 115263 406408
rect 114461 406403 114527 406406
rect 115197 406403 115263 406406
rect 181478 406268 181484 406332
rect 181548 406330 181554 406332
rect 191966 406330 191972 406332
rect 181548 406270 191972 406330
rect 181548 406268 181554 406270
rect 191966 406268 191972 406270
rect 192036 406268 192042 406332
rect 67265 405650 67331 405653
rect 115841 405650 115907 405653
rect 67265 405648 68908 405650
rect 67265 405592 67270 405648
rect 67326 405592 68908 405648
rect 67265 405590 68908 405592
rect 112700 405648 115907 405650
rect 112700 405592 115846 405648
rect 115902 405592 115907 405648
rect 112700 405590 115907 405592
rect 67265 405587 67331 405590
rect 115841 405587 115907 405590
rect 191649 405650 191715 405653
rect 191649 405648 193660 405650
rect 191649 405592 191654 405648
rect 191710 405592 193660 405648
rect 191649 405590 193660 405592
rect 191649 405587 191715 405590
rect 254117 405378 254183 405381
rect 253460 405376 254183 405378
rect 253460 405320 254122 405376
rect 254178 405320 254183 405376
rect 253460 405318 254183 405320
rect 254117 405315 254183 405318
rect 582649 404970 582715 404973
rect 583520 404970 584960 405060
rect 582649 404968 584960 404970
rect 582649 404912 582654 404968
rect 582710 404912 584960 404968
rect 582649 404910 584960 404912
rect 582649 404907 582715 404910
rect 583520 404820 584960 404910
rect 66805 404562 66871 404565
rect 115841 404562 115907 404565
rect 66805 404560 68908 404562
rect 66805 404504 66810 404560
rect 66866 404504 68908 404560
rect 66805 404502 68908 404504
rect 112700 404560 115907 404562
rect 112700 404504 115846 404560
rect 115902 404504 115907 404560
rect 112700 404502 115907 404504
rect 66805 404499 66871 404502
rect 115841 404499 115907 404502
rect 191741 404290 191807 404293
rect 191741 404288 193660 404290
rect 191741 404232 191746 404288
rect 191802 404232 193660 404288
rect 191741 404230 193660 404232
rect 191741 404227 191807 404230
rect 256877 404018 256943 404021
rect 253460 404016 256943 404018
rect 253460 403960 256882 404016
rect 256938 403960 256943 404016
rect 253460 403958 256943 403960
rect 256877 403955 256943 403958
rect 66069 403746 66135 403749
rect 66069 403744 68908 403746
rect 66069 403688 66074 403744
rect 66130 403688 68908 403744
rect 66069 403686 68908 403688
rect 66069 403683 66135 403686
rect 180425 403610 180491 403613
rect 184933 403610 184999 403613
rect 180425 403608 184999 403610
rect 180425 403552 180430 403608
rect 180486 403552 184938 403608
rect 184994 403552 184999 403608
rect 180425 403550 184999 403552
rect 180425 403547 180491 403550
rect 184933 403547 184999 403550
rect 115841 403474 115907 403477
rect 112700 403472 115907 403474
rect 112700 403416 115846 403472
rect 115902 403416 115907 403472
rect 112700 403414 115907 403416
rect 115841 403411 115907 403414
rect 193121 402930 193187 402933
rect 193121 402928 193660 402930
rect 193121 402872 193126 402928
rect 193182 402872 193660 402928
rect 193121 402870 193660 402872
rect 193121 402867 193187 402870
rect 66662 402596 66668 402660
rect 66732 402658 66738 402660
rect 67817 402658 67883 402661
rect 66732 402656 68908 402658
rect 66732 402600 67822 402656
rect 67878 402600 68908 402656
rect 66732 402598 68908 402600
rect 66732 402596 66738 402598
rect 67817 402595 67883 402598
rect 112110 402596 112116 402660
rect 112180 402596 112186 402660
rect 254710 402658 254716 402660
rect 253460 402598 254716 402658
rect 254710 402596 254716 402598
rect 254780 402658 254786 402660
rect 255313 402658 255379 402661
rect 254780 402656 255379 402658
rect 254780 402600 255318 402656
rect 255374 402600 255379 402656
rect 254780 402598 255379 402600
rect 254780 402596 254786 402598
rect 112118 402386 112178 402596
rect 255313 402595 255379 402598
rect 113449 402386 113515 402389
rect 112118 402384 113515 402386
rect 112118 402356 113454 402384
rect 112148 402328 113454 402356
rect 113510 402328 113515 402384
rect 112148 402326 113515 402328
rect 113449 402323 113515 402326
rect 162577 401706 162643 401709
rect 162710 401706 162716 401708
rect 162577 401704 162716 401706
rect 162577 401648 162582 401704
rect 162638 401648 162716 401704
rect 162577 401646 162716 401648
rect 162577 401643 162643 401646
rect 162710 401644 162716 401646
rect 162780 401644 162786 401708
rect 163497 401706 163563 401709
rect 162902 401704 163563 401706
rect 162902 401648 163502 401704
rect 163558 401648 163563 401704
rect 162902 401646 163563 401648
rect 66805 401570 66871 401573
rect 66805 401568 68908 401570
rect 66805 401512 66810 401568
rect 66866 401512 68908 401568
rect 66805 401510 68908 401512
rect 66805 401507 66871 401510
rect 162710 401508 162716 401572
rect 162780 401570 162786 401572
rect 162902 401570 162962 401646
rect 163497 401643 163563 401646
rect 162780 401510 162962 401570
rect 191557 401570 191623 401573
rect 191557 401568 193660 401570
rect 191557 401512 191562 401568
rect 191618 401512 193660 401568
rect 191557 401510 193660 401512
rect 162780 401508 162786 401510
rect 191557 401507 191623 401510
rect 115749 401298 115815 401301
rect 255405 401298 255471 401301
rect 112700 401296 115815 401298
rect 112700 401240 115754 401296
rect 115810 401240 115815 401296
rect 112700 401238 115815 401240
rect 253460 401296 255471 401298
rect 253460 401240 255410 401296
rect 255466 401240 255471 401296
rect 253460 401238 255471 401240
rect 115749 401235 115815 401238
rect 255405 401235 255471 401238
rect 67357 400482 67423 400485
rect 115565 400482 115631 400485
rect 67357 400480 68908 400482
rect 67357 400424 67362 400480
rect 67418 400424 68908 400480
rect 67357 400422 68908 400424
rect 112700 400480 115631 400482
rect 112700 400424 115570 400480
rect 115626 400424 115631 400480
rect 112700 400422 115631 400424
rect 67357 400419 67423 400422
rect 115565 400419 115631 400422
rect 113030 400148 113036 400212
rect 113100 400210 113106 400212
rect 148961 400210 149027 400213
rect 113100 400208 149027 400210
rect 113100 400152 148966 400208
rect 149022 400152 149027 400208
rect 113100 400150 149027 400152
rect 113100 400148 113106 400150
rect 148961 400147 149027 400150
rect 180609 400210 180675 400213
rect 181897 400210 181963 400213
rect 180609 400208 181963 400210
rect 180609 400152 180614 400208
rect 180670 400152 181902 400208
rect 181958 400152 181963 400208
rect 180609 400150 181963 400152
rect 180609 400147 180675 400150
rect 181897 400147 181963 400150
rect 191741 400210 191807 400213
rect 191741 400208 193660 400210
rect 191741 400152 191746 400208
rect 191802 400152 193660 400208
rect 191741 400150 193660 400152
rect 191741 400147 191807 400150
rect 255405 399938 255471 399941
rect 253460 399936 255471 399938
rect 253460 399880 255410 399936
rect 255466 399880 255471 399936
rect 253460 399878 255471 399880
rect 255405 399875 255471 399878
rect 66805 399666 66871 399669
rect 66805 399664 68908 399666
rect 66805 399608 66810 399664
rect 66866 399608 68908 399664
rect 66805 399606 68908 399608
rect 66805 399603 66871 399606
rect 115841 399394 115907 399397
rect 112700 399392 115907 399394
rect 112700 399336 115846 399392
rect 115902 399336 115907 399392
rect 112700 399334 115907 399336
rect 115841 399331 115907 399334
rect 66529 398578 66595 398581
rect 191741 398578 191807 398581
rect 255405 398578 255471 398581
rect 66529 398576 68908 398578
rect 66529 398520 66534 398576
rect 66590 398520 68908 398576
rect 66529 398518 68908 398520
rect 191741 398576 193660 398578
rect 191741 398520 191746 398576
rect 191802 398520 193660 398576
rect 191741 398518 193660 398520
rect 253460 398576 255471 398578
rect 253460 398520 255410 398576
rect 255466 398520 255471 398576
rect 253460 398518 255471 398520
rect 66529 398515 66595 398518
rect 191741 398515 191807 398518
rect 255405 398515 255471 398518
rect 115841 398306 115907 398309
rect 112700 398304 115907 398306
rect 112700 398248 115846 398304
rect 115902 398248 115907 398304
rect 112700 398246 115907 398248
rect 115841 398243 115907 398246
rect 184790 397972 184796 398036
rect 184860 398034 184866 398036
rect 193305 398034 193371 398037
rect 184860 398032 193371 398034
rect 184860 397976 193310 398032
rect 193366 397976 193371 398032
rect 184860 397974 193371 397976
rect 184860 397972 184866 397974
rect 193305 397971 193371 397974
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 67081 397490 67147 397493
rect 67449 397490 67515 397493
rect 67081 397488 68908 397490
rect 67081 397432 67086 397488
rect 67142 397432 67454 397488
rect 67510 397432 68908 397488
rect 67081 397430 68908 397432
rect 67081 397427 67147 397430
rect 67449 397427 67515 397430
rect 65977 397354 66043 397357
rect 66294 397354 66300 397356
rect 65977 397352 66300 397354
rect 65977 397296 65982 397352
rect 66038 397296 66300 397352
rect 65977 397294 66300 397296
rect 65977 397291 66043 397294
rect 66294 397292 66300 397294
rect 66364 397292 66370 397356
rect 115565 397218 115631 397221
rect 112700 397216 115631 397218
rect 112700 397160 115570 397216
rect 115626 397160 115631 397216
rect 112700 397158 115631 397160
rect 115565 397155 115631 397158
rect 67541 396402 67607 396405
rect 114318 396402 114324 396404
rect 67541 396400 68908 396402
rect 67541 396344 67546 396400
rect 67602 396344 68908 396400
rect 67541 396342 68908 396344
rect 112700 396342 114324 396402
rect 67541 396339 67607 396342
rect 114318 396340 114324 396342
rect 114388 396402 114394 396404
rect 115105 396402 115171 396405
rect 114388 396400 115171 396402
rect 114388 396344 115110 396400
rect 115166 396344 115171 396400
rect 114388 396342 115171 396344
rect 114388 396340 114394 396342
rect 115105 396339 115171 396342
rect 189717 396130 189783 396133
rect 193630 396130 193690 397188
rect 254025 396946 254091 396949
rect 252908 396944 254091 396946
rect 252908 396916 254030 396944
rect 252878 396888 254030 396916
rect 254086 396888 254091 396944
rect 252878 396886 254091 396888
rect 252878 396812 252938 396886
rect 254025 396883 254091 396886
rect 252870 396748 252876 396812
rect 252940 396748 252946 396812
rect 189717 396128 193690 396130
rect 189717 396072 189722 396128
rect 189778 396072 193690 396128
rect 189717 396070 193690 396072
rect 189717 396067 189783 396070
rect 67265 395314 67331 395317
rect 115841 395314 115907 395317
rect 67265 395312 68908 395314
rect 67265 395256 67270 395312
rect 67326 395256 68908 395312
rect 67265 395254 68908 395256
rect 112700 395312 115907 395314
rect 112700 395256 115846 395312
rect 115902 395256 115907 395312
rect 112700 395254 115907 395256
rect 67265 395251 67331 395254
rect 115841 395251 115907 395254
rect 155953 394770 156019 394773
rect 193630 394770 193690 395828
rect 254025 395586 254091 395589
rect 253460 395584 254091 395586
rect 253460 395528 254030 395584
rect 254086 395528 254091 395584
rect 253460 395526 254091 395528
rect 254025 395523 254091 395526
rect 258901 395314 258967 395317
rect 276422 395314 276428 395316
rect 258901 395312 276428 395314
rect 258901 395256 258906 395312
rect 258962 395256 276428 395312
rect 258901 395254 276428 395256
rect 258901 395251 258967 395254
rect 276422 395252 276428 395254
rect 276492 395252 276498 395316
rect 155953 394768 193690 394770
rect 155953 394712 155958 394768
rect 156014 394712 193690 394768
rect 155953 394710 193690 394712
rect 155953 394707 156019 394710
rect 67725 394498 67791 394501
rect 191005 394498 191071 394501
rect 67725 394496 68908 394498
rect 67725 394440 67730 394496
rect 67786 394440 68908 394496
rect 67725 394438 68908 394440
rect 191005 394496 193660 394498
rect 191005 394440 191010 394496
rect 191066 394440 193660 394496
rect 191005 394438 193660 394440
rect 67725 394435 67791 394438
rect 191005 394435 191071 394438
rect 115841 394226 115907 394229
rect 255497 394226 255563 394229
rect 112700 394224 115907 394226
rect 112700 394168 115846 394224
rect 115902 394168 115907 394224
rect 112700 394166 115907 394168
rect 253460 394224 255563 394226
rect 253460 394168 255502 394224
rect 255558 394168 255563 394224
rect 253460 394166 255563 394168
rect 115841 394163 115907 394166
rect 255497 394163 255563 394166
rect 112846 393892 112852 393956
rect 112916 393954 112922 393956
rect 181989 393954 182055 393957
rect 186773 393954 186839 393957
rect 112916 393952 186839 393954
rect 112916 393896 181994 393952
rect 182050 393896 186778 393952
rect 186834 393896 186839 393952
rect 112916 393894 186839 393896
rect 112916 393892 112922 393894
rect 181989 393891 182055 393894
rect 186773 393891 186839 393894
rect 65977 393410 66043 393413
rect 180609 393410 180675 393413
rect 180742 393410 180748 393412
rect 65977 393408 68908 393410
rect 65977 393352 65982 393408
rect 66038 393352 68908 393408
rect 65977 393350 68908 393352
rect 180609 393408 180748 393410
rect 180609 393352 180614 393408
rect 180670 393352 180748 393408
rect 180609 393350 180748 393352
rect 65977 393347 66043 393350
rect 180609 393347 180675 393350
rect 180742 393348 180748 393350
rect 180812 393348 180818 393412
rect 115841 393138 115907 393141
rect 180701 393140 180767 393141
rect 180701 393138 180748 393140
rect 112700 393136 115907 393138
rect 112700 393080 115846 393136
rect 115902 393080 115907 393136
rect 112700 393078 115907 393080
rect 180656 393136 180748 393138
rect 180812 393138 180818 393140
rect 191925 393138 191991 393141
rect 180656 393080 180706 393136
rect 180656 393078 180748 393080
rect 115841 393075 115907 393078
rect 180701 393076 180748 393078
rect 180812 393078 180894 393138
rect 191925 393136 193660 393138
rect 191925 393080 191930 393136
rect 191986 393080 193660 393136
rect 191925 393078 193660 393080
rect 180812 393076 180818 393078
rect 180701 393075 180767 393076
rect 191925 393075 191991 393078
rect 254301 392866 254367 392869
rect 253460 392864 254367 392866
rect 253460 392808 254306 392864
rect 254362 392808 254367 392864
rect 253460 392806 254367 392808
rect 254301 392803 254367 392806
rect 137829 392594 137895 392597
rect 145557 392594 145623 392597
rect 137829 392592 145623 392594
rect 137829 392536 137834 392592
rect 137890 392536 145562 392592
rect 145618 392536 145623 392592
rect 137829 392534 145623 392536
rect 137829 392531 137895 392534
rect 145557 392531 145623 392534
rect 66805 392322 66871 392325
rect 66805 392320 68908 392322
rect 66805 392264 66810 392320
rect 66866 392264 68908 392320
rect 66805 392262 68908 392264
rect 66805 392259 66871 392262
rect 115841 392050 115907 392053
rect 112700 392048 115907 392050
rect 112700 391992 115846 392048
rect 115902 391992 115907 392048
rect 112700 391990 115907 391992
rect 115841 391987 115907 391990
rect 253933 392050 253999 392053
rect 254710 392050 254716 392052
rect 253933 392048 254716 392050
rect 253933 391992 253938 392048
rect 253994 391992 254716 392048
rect 253933 391990 254716 391992
rect 253933 391987 253999 391990
rect 254710 391988 254716 391990
rect 254780 391988 254786 392052
rect 191741 391778 191807 391781
rect 191741 391776 193660 391778
rect 191741 391720 191746 391776
rect 191802 391720 193660 391776
rect 191741 391718 193660 391720
rect 191741 391715 191807 391718
rect 111926 391580 111932 391644
rect 111996 391642 112002 391644
rect 113030 391642 113036 391644
rect 111996 391582 113036 391642
rect 111996 391580 112002 391582
rect 113030 391580 113036 391582
rect 113100 391580 113106 391644
rect 583520 391628 584960 391868
rect 63401 391506 63467 391509
rect 114502 391506 114508 391508
rect 63401 391504 80070 391506
rect 63401 391448 63406 391504
rect 63462 391448 80070 391504
rect 63401 391446 80070 391448
rect 63401 391443 63467 391446
rect 69430 390690 69490 391204
rect 80010 391098 80070 391446
rect 108990 391446 114508 391506
rect 80010 391038 85130 391098
rect 72417 390962 72483 390965
rect 72734 390962 72740 390964
rect 72417 390960 72740 390962
rect 72417 390904 72422 390960
rect 72478 390904 72740 390960
rect 72417 390902 72740 390904
rect 72417 390899 72483 390902
rect 72734 390900 72740 390902
rect 72804 390900 72810 390964
rect 84377 390962 84443 390965
rect 84510 390962 84516 390964
rect 84377 390960 84516 390962
rect 84377 390904 84382 390960
rect 84438 390904 84516 390960
rect 84377 390902 84516 390904
rect 84377 390899 84443 390902
rect 84510 390900 84516 390902
rect 84580 390900 84586 390964
rect 85070 390962 85130 391038
rect 87137 390962 87203 390965
rect 87873 390962 87939 390965
rect 85070 390960 87939 390962
rect 85070 390904 87142 390960
rect 87198 390904 87878 390960
rect 87934 390904 87939 390960
rect 85070 390902 87939 390904
rect 87137 390899 87203 390902
rect 87873 390899 87939 390902
rect 99649 390962 99715 390965
rect 104249 390964 104315 390965
rect 100150 390962 100156 390964
rect 99649 390960 100156 390962
rect 99649 390904 99654 390960
rect 99710 390904 100156 390960
rect 99649 390902 100156 390904
rect 99649 390899 99715 390902
rect 100150 390900 100156 390902
rect 100220 390900 100226 390964
rect 104198 390900 104204 390964
rect 104268 390962 104315 390964
rect 104268 390960 104360 390962
rect 104310 390904 104360 390960
rect 104268 390902 104360 390904
rect 104268 390900 104315 390902
rect 104934 390900 104940 390964
rect 105004 390962 105010 390964
rect 105261 390962 105327 390965
rect 105004 390960 105327 390962
rect 105004 390904 105266 390960
rect 105322 390904 105327 390960
rect 105004 390902 105327 390904
rect 105004 390900 105010 390902
rect 104249 390899 104315 390900
rect 105261 390899 105327 390902
rect 105905 390962 105971 390965
rect 108990 390962 109050 391446
rect 114502 391444 114508 391446
rect 114572 391444 114578 391508
rect 112670 391098 112730 391204
rect 112897 391098 112963 391101
rect 112670 391096 112963 391098
rect 112670 391040 112902 391096
rect 112958 391040 112963 391096
rect 112670 391038 112963 391040
rect 112897 391035 112963 391038
rect 192477 391098 192543 391101
rect 193397 391098 193463 391101
rect 192477 391096 193463 391098
rect 192477 391040 192482 391096
rect 192538 391040 193402 391096
rect 193458 391040 193463 391096
rect 192477 391038 193463 391040
rect 192477 391035 192543 391038
rect 193397 391035 193463 391038
rect 111977 390964 112043 390965
rect 105905 390960 109050 390962
rect 105905 390904 105910 390960
rect 105966 390904 109050 390960
rect 105905 390902 109050 390904
rect 105905 390899 105971 390902
rect 111926 390900 111932 390964
rect 111996 390962 112043 390964
rect 155677 390962 155743 390965
rect 156597 390962 156663 390965
rect 111996 390960 112088 390962
rect 112038 390904 112088 390960
rect 111996 390902 112088 390904
rect 112302 390960 156663 390962
rect 112302 390904 155682 390960
rect 155738 390904 156602 390960
rect 156658 390904 156663 390960
rect 112302 390902 156663 390904
rect 111996 390900 112043 390902
rect 111977 390899 112043 390900
rect 79910 390764 79916 390828
rect 79980 390826 79986 390828
rect 80145 390826 80211 390829
rect 80973 390826 81039 390829
rect 79980 390824 81039 390826
rect 79980 390768 80150 390824
rect 80206 390768 80978 390824
rect 81034 390768 81039 390824
rect 79980 390766 81039 390768
rect 79980 390764 79986 390766
rect 80145 390763 80211 390766
rect 80973 390763 81039 390766
rect 82854 390764 82860 390828
rect 82924 390826 82930 390828
rect 83181 390826 83247 390829
rect 82924 390824 83247 390826
rect 82924 390768 83186 390824
rect 83242 390768 83247 390824
rect 82924 390766 83247 390768
rect 82924 390764 82930 390766
rect 83181 390763 83247 390766
rect 103789 390826 103855 390829
rect 112302 390826 112362 390902
rect 155677 390899 155743 390902
rect 156597 390899 156663 390902
rect 180149 390962 180215 390965
rect 212441 390962 212507 390965
rect 180149 390960 212507 390962
rect 180149 390904 180154 390960
rect 180210 390904 212446 390960
rect 212502 390904 212507 390960
rect 180149 390902 212507 390904
rect 180149 390899 180215 390902
rect 212441 390899 212507 390902
rect 249701 390962 249767 390965
rect 252878 390962 252938 391476
rect 249701 390960 252938 390962
rect 249701 390904 249706 390960
rect 249762 390904 252938 390960
rect 249701 390902 252938 390904
rect 249701 390899 249767 390902
rect 103789 390824 112362 390826
rect 103789 390768 103794 390824
rect 103850 390768 112362 390824
rect 103789 390766 112362 390768
rect 112897 390826 112963 390829
rect 182817 390826 182883 390829
rect 112897 390824 182883 390826
rect 112897 390768 112902 390824
rect 112958 390768 182822 390824
rect 182878 390768 182883 390824
rect 112897 390766 182883 390768
rect 103789 390763 103855 390766
rect 112897 390763 112963 390766
rect 182817 390763 182883 390766
rect 158437 390690 158503 390693
rect 192017 390692 192083 390693
rect 191966 390690 191972 390692
rect 69430 390688 158503 390690
rect 69430 390632 158442 390688
rect 158498 390632 158503 390688
rect 69430 390630 158503 390632
rect 191926 390630 191972 390690
rect 192036 390688 192083 390692
rect 192078 390632 192083 390688
rect 158437 390627 158503 390630
rect 191966 390628 191972 390630
rect 192036 390628 192083 390632
rect 192017 390627 192083 390628
rect 82169 390554 82235 390557
rect 84694 390554 84700 390556
rect 82169 390552 84700 390554
rect 82169 390496 82174 390552
rect 82230 390496 84700 390552
rect 82169 390494 84700 390496
rect 82169 390491 82235 390494
rect 84694 390492 84700 390494
rect 84764 390554 84770 390556
rect 112846 390554 112852 390556
rect 84764 390494 112852 390554
rect 84764 390492 84770 390494
rect 112846 390492 112852 390494
rect 112916 390492 112922 390556
rect 284385 390554 284451 390557
rect 582741 390554 582807 390557
rect 284385 390552 582807 390554
rect 284385 390496 284390 390552
rect 284446 390496 582746 390552
rect 582802 390496 582807 390552
rect 284385 390494 582807 390496
rect 284385 390491 284451 390494
rect 582741 390491 582807 390494
rect 77201 390420 77267 390421
rect 77150 390418 77156 390420
rect 77110 390358 77156 390418
rect 77220 390416 77267 390420
rect 77262 390360 77267 390416
rect 77150 390356 77156 390358
rect 77220 390356 77267 390360
rect 91318 390356 91324 390420
rect 91388 390418 91394 390420
rect 92013 390418 92079 390421
rect 91388 390416 92079 390418
rect 91388 390360 92018 390416
rect 92074 390360 92079 390416
rect 91388 390358 92079 390360
rect 91388 390356 91394 390358
rect 77201 390355 77267 390356
rect 92013 390355 92079 390358
rect 96654 390356 96660 390420
rect 96724 390418 96730 390420
rect 96981 390418 97047 390421
rect 96724 390416 97047 390418
rect 96724 390360 96986 390416
rect 97042 390360 97047 390416
rect 96724 390358 97047 390360
rect 96724 390356 96730 390358
rect 96981 390355 97047 390358
rect 108297 389874 108363 389877
rect 118693 389874 118759 389877
rect 108297 389872 118759 389874
rect 108297 389816 108302 389872
rect 108358 389816 118698 389872
rect 118754 389816 118759 389872
rect 108297 389814 118759 389816
rect 108297 389811 108363 389814
rect 118693 389811 118759 389814
rect 154389 389874 154455 389877
rect 188521 389874 188587 389877
rect 154389 389872 188587 389874
rect 154389 389816 154394 389872
rect 154450 389816 188526 389872
rect 188582 389816 188587 389872
rect 154389 389814 188587 389816
rect 154389 389811 154455 389814
rect 188521 389811 188587 389814
rect 190310 389812 190316 389876
rect 190380 389874 190386 389876
rect 204345 389874 204411 389877
rect 190380 389872 204411 389874
rect 190380 389816 204350 389872
rect 204406 389816 204411 389872
rect 190380 389814 204411 389816
rect 190380 389812 190386 389814
rect 204345 389811 204411 389814
rect 250437 389466 250503 389469
rect 254025 389466 254091 389469
rect 250437 389464 254091 389466
rect 250437 389408 250442 389464
rect 250498 389408 254030 389464
rect 254086 389408 254091 389464
rect 250437 389406 254091 389408
rect 250437 389403 250503 389406
rect 254025 389403 254091 389406
rect 88190 389268 88196 389332
rect 88260 389330 88266 389332
rect 106733 389330 106799 389333
rect 230565 389330 230631 389333
rect 249742 389330 249748 389332
rect 88260 389328 109050 389330
rect 88260 389272 106738 389328
rect 106794 389272 109050 389328
rect 88260 389270 109050 389272
rect 88260 389268 88266 389270
rect 106733 389267 106799 389270
rect 57789 389194 57855 389197
rect 99281 389194 99347 389197
rect 57789 389192 99347 389194
rect 57789 389136 57794 389192
rect 57850 389136 99286 389192
rect 99342 389136 99347 389192
rect 57789 389134 99347 389136
rect 108990 389194 109050 389270
rect 230565 389328 249748 389330
rect 230565 389272 230570 389328
rect 230626 389272 249748 389328
rect 230565 389270 249748 389272
rect 230565 389267 230631 389270
rect 249742 389268 249748 389270
rect 249812 389268 249818 389332
rect 251030 389268 251036 389332
rect 251100 389330 251106 389332
rect 254209 389330 254275 389333
rect 251100 389328 254275 389330
rect 251100 389272 254214 389328
rect 254270 389272 254275 389328
rect 251100 389270 254275 389272
rect 251100 389268 251106 389270
rect 254209 389267 254275 389270
rect 123569 389194 123635 389197
rect 108990 389192 123635 389194
rect 108990 389136 123574 389192
rect 123630 389136 123635 389192
rect 108990 389134 123635 389136
rect 57789 389131 57855 389134
rect 99281 389131 99347 389134
rect 123569 389131 123635 389134
rect 181989 389194 182055 389197
rect 187693 389194 187759 389197
rect 181989 389192 187759 389194
rect 181989 389136 181994 389192
rect 182050 389136 187698 389192
rect 187754 389136 187759 389192
rect 181989 389134 187759 389136
rect 181989 389131 182055 389134
rect 187693 389131 187759 389134
rect 204805 389194 204871 389197
rect 284385 389194 284451 389197
rect 204805 389192 284451 389194
rect 204805 389136 204810 389192
rect 204866 389136 284390 389192
rect 284446 389136 284451 389192
rect 204805 389134 284451 389136
rect 204805 389131 204871 389134
rect 284385 389131 284451 389134
rect 105721 389058 105787 389061
rect 106089 389058 106155 389061
rect 105721 389056 106155 389058
rect 105721 389000 105726 389056
rect 105782 389000 106094 389056
rect 106150 389000 106155 389056
rect 105721 388998 106155 389000
rect 105721 388995 105787 388998
rect 106089 388995 106155 388998
rect 244222 388996 244228 389060
rect 244292 389058 244298 389060
rect 244733 389058 244799 389061
rect 248597 389060 248663 389061
rect 248597 389058 248644 389060
rect 244292 389056 244799 389058
rect 244292 389000 244738 389056
rect 244794 389000 244799 389056
rect 244292 388998 244799 389000
rect 248552 389056 248644 389058
rect 248708 389058 248714 389060
rect 249374 389058 249380 389060
rect 248552 389000 248602 389056
rect 248552 388998 248644 389000
rect 244292 388996 244298 388998
rect 244733 388995 244799 388998
rect 248597 388996 248644 388998
rect 248708 388998 249380 389058
rect 248708 388996 248714 388998
rect 249374 388996 249380 388998
rect 249444 388996 249450 389060
rect 249517 389058 249583 389061
rect 263593 389058 263659 389061
rect 249517 389056 263659 389058
rect 249517 389000 249522 389056
rect 249578 389000 263598 389056
rect 263654 389000 263659 389056
rect 249517 388998 263659 389000
rect 248597 388995 248663 388996
rect 249517 388995 249583 388998
rect 263593 388995 263659 388998
rect 72734 388860 72740 388924
rect 72804 388922 72810 388924
rect 173525 388922 173591 388925
rect 72804 388920 173591 388922
rect 72804 388864 173530 388920
rect 173586 388864 173591 388920
rect 72804 388862 173591 388864
rect 72804 388860 72810 388862
rect 173525 388859 173591 388862
rect 77201 388786 77267 388789
rect 169702 388786 169708 388788
rect 77201 388784 169708 388786
rect 77201 388728 77206 388784
rect 77262 388728 169708 388784
rect 77201 388726 169708 388728
rect 77201 388723 77267 388726
rect 169702 388724 169708 388726
rect 169772 388724 169778 388788
rect 100753 388650 100819 388653
rect 101254 388650 101260 388652
rect 100753 388648 101260 388650
rect 100753 388592 100758 388648
rect 100814 388592 101260 388648
rect 100753 388590 101260 388592
rect 100753 388587 100819 388590
rect 101254 388588 101260 388590
rect 101324 388650 101330 388652
rect 236637 388650 236703 388653
rect 237189 388650 237255 388653
rect 101324 388648 237255 388650
rect 101324 388592 236642 388648
rect 236698 388592 237194 388648
rect 237250 388592 237255 388648
rect 101324 388590 237255 388592
rect 101324 388588 101330 388590
rect 236637 388587 236703 388590
rect 237189 388587 237255 388590
rect 77385 388514 77451 388517
rect 78254 388514 78260 388516
rect 77385 388512 78260 388514
rect 77385 388456 77390 388512
rect 77446 388456 78260 388512
rect 77385 388454 78260 388456
rect 77385 388451 77451 388454
rect 78254 388452 78260 388454
rect 78324 388452 78330 388516
rect 80237 388514 80303 388517
rect 80646 388514 80652 388516
rect 80237 388512 80652 388514
rect 80237 388456 80242 388512
rect 80298 388456 80652 388512
rect 80237 388454 80652 388456
rect 80237 388451 80303 388454
rect 80646 388452 80652 388454
rect 80716 388452 80722 388516
rect 81433 388514 81499 388517
rect 247217 388516 247283 388517
rect 82486 388514 82492 388516
rect 81433 388512 82492 388514
rect 81433 388456 81438 388512
rect 81494 388456 82492 388512
rect 81433 388454 82492 388456
rect 81433 388451 81499 388454
rect 82486 388452 82492 388454
rect 82556 388452 82562 388516
rect 247166 388514 247172 388516
rect 247126 388454 247172 388514
rect 247236 388512 247283 388516
rect 247278 388456 247283 388512
rect 247166 388452 247172 388454
rect 247236 388452 247283 388456
rect 247217 388451 247283 388452
rect 83958 388316 83964 388380
rect 84028 388378 84034 388380
rect 85021 388378 85087 388381
rect 84028 388376 85087 388378
rect 84028 388320 85026 388376
rect 85082 388320 85087 388376
rect 84028 388318 85087 388320
rect 84028 388316 84034 388318
rect 85021 388315 85087 388318
rect 245561 388378 245627 388381
rect 262397 388378 262463 388381
rect 245561 388376 262463 388378
rect 245561 388320 245566 388376
rect 245622 388320 262402 388376
rect 262458 388320 262463 388376
rect 245561 388318 262463 388320
rect 245561 388315 245627 388318
rect 262397 388315 262463 388318
rect 96654 387772 96660 387836
rect 96724 387834 96730 387836
rect 97533 387834 97599 387837
rect 96724 387832 97599 387834
rect 96724 387776 97538 387832
rect 97594 387776 97599 387832
rect 96724 387774 97599 387776
rect 96724 387772 96730 387774
rect 97533 387771 97599 387774
rect 73061 387698 73127 387701
rect 75126 387698 75132 387700
rect 73061 387696 75132 387698
rect 73061 387640 73066 387696
rect 73122 387640 75132 387696
rect 73061 387638 75132 387640
rect 73061 387635 73127 387638
rect 75126 387636 75132 387638
rect 75196 387636 75202 387700
rect 173525 387698 173591 387701
rect 173801 387698 173867 387701
rect 191833 387698 191899 387701
rect 173525 387696 191899 387698
rect 173525 387640 173530 387696
rect 173586 387640 173806 387696
rect 173862 387640 191838 387696
rect 191894 387640 191899 387696
rect 173525 387638 191899 387640
rect 173525 387635 173591 387638
rect 173801 387635 173867 387638
rect 191833 387635 191899 387638
rect 192017 387698 192083 387701
rect 195237 387698 195303 387701
rect 192017 387696 195303 387698
rect 192017 387640 192022 387696
rect 192078 387640 195242 387696
rect 195298 387640 195303 387696
rect 192017 387638 195303 387640
rect 192017 387635 192083 387638
rect 195237 387635 195303 387638
rect 197353 387698 197419 387701
rect 198181 387698 198247 387701
rect 280245 387698 280311 387701
rect 281441 387698 281507 387701
rect 197353 387696 281507 387698
rect 197353 387640 197358 387696
rect 197414 387640 198186 387696
rect 198242 387640 280250 387696
rect 280306 387640 281446 387696
rect 281502 387640 281507 387696
rect 197353 387638 281507 387640
rect 197353 387635 197419 387638
rect 198181 387635 198247 387638
rect 280245 387635 280311 387638
rect 281441 387635 281507 387638
rect 178033 387562 178099 387565
rect 178769 387562 178835 387565
rect 178033 387560 178835 387562
rect 178033 387504 178038 387560
rect 178094 387504 178774 387560
rect 178830 387504 178835 387560
rect 178033 387502 178835 387504
rect 178033 387499 178099 387502
rect 178769 387499 178835 387502
rect 180057 387562 180123 387565
rect 180609 387562 180675 387565
rect 213453 387562 213519 387565
rect 180057 387560 213519 387562
rect 180057 387504 180062 387560
rect 180118 387504 180614 387560
rect 180670 387504 213458 387560
rect 213514 387504 213519 387560
rect 180057 387502 213519 387504
rect 180057 387499 180123 387502
rect 180609 387499 180675 387502
rect 213453 387499 213519 387502
rect 191833 387426 191899 387429
rect 197353 387426 197419 387429
rect 191833 387424 197419 387426
rect 191833 387368 191838 387424
rect 191894 387368 197358 387424
rect 197414 387368 197419 387424
rect 191833 387366 197419 387368
rect 191833 387363 191899 387366
rect 197353 387363 197419 387366
rect 83549 387290 83615 387293
rect 89662 387290 89668 387292
rect 83549 387288 89668 387290
rect 83549 387232 83554 387288
rect 83610 387232 89668 387288
rect 83549 387230 89668 387232
rect 83549 387227 83615 387230
rect 89662 387228 89668 387230
rect 89732 387228 89738 387292
rect 86861 387154 86927 387157
rect 117957 387154 118023 387157
rect 86861 387152 118023 387154
rect 86861 387096 86866 387152
rect 86922 387096 117962 387152
rect 118018 387096 118023 387152
rect 86861 387094 118023 387096
rect 86861 387091 86927 387094
rect 117957 387091 118023 387094
rect 48129 387018 48195 387021
rect 178033 387018 178099 387021
rect 48129 387016 178099 387018
rect 48129 386960 48134 387016
rect 48190 386960 178038 387016
rect 178094 386960 178099 387016
rect 48129 386958 178099 386960
rect 48129 386955 48195 386958
rect 178033 386955 178099 386958
rect 238017 387018 238083 387021
rect 247718 387018 247724 387020
rect 238017 387016 247724 387018
rect 238017 386960 238022 387016
rect 238078 386960 247724 387016
rect 238017 386958 247724 386960
rect 238017 386955 238083 386958
rect 247718 386956 247724 386958
rect 247788 386956 247794 387020
rect 67265 386338 67331 386341
rect 139393 386338 139459 386341
rect 67265 386336 139459 386338
rect 67265 386280 67270 386336
rect 67326 386280 139398 386336
rect 139454 386280 139459 386336
rect 67265 386278 139459 386280
rect 67265 386275 67331 386278
rect 139393 386275 139459 386278
rect 169702 386276 169708 386340
rect 169772 386338 169778 386340
rect 170806 386338 170812 386340
rect 169772 386278 170812 386338
rect 169772 386276 169778 386278
rect 170806 386276 170812 386278
rect 170876 386338 170882 386340
rect 204805 386338 204871 386341
rect 170876 386336 204871 386338
rect 170876 386280 204810 386336
rect 204866 386280 204871 386336
rect 170876 386278 204871 386280
rect 170876 386276 170882 386278
rect 204805 386275 204871 386278
rect 188429 386202 188495 386205
rect 244917 386202 244983 386205
rect 188429 386200 244983 386202
rect 188429 386144 188434 386200
rect 188490 386144 244922 386200
rect 244978 386144 244983 386200
rect 188429 386142 244983 386144
rect 188429 386139 188495 386142
rect 244917 386139 244983 386142
rect 167637 386066 167703 386069
rect 201125 386066 201191 386069
rect 167637 386064 201191 386066
rect 167637 386008 167642 386064
rect 167698 386008 201130 386064
rect 201186 386008 201191 386064
rect 167637 386006 201191 386008
rect 167637 386003 167703 386006
rect 201125 386003 201191 386006
rect 203517 386066 203583 386069
rect 283097 386066 283163 386069
rect 203517 386064 283163 386066
rect 203517 386008 203522 386064
rect 203578 386008 283102 386064
rect 283158 386008 283163 386064
rect 203517 386006 283163 386008
rect 203517 386003 203583 386006
rect 283097 386003 283163 386006
rect 89621 385794 89687 385797
rect 100702 385794 100708 385796
rect 89621 385792 100708 385794
rect 89621 385736 89626 385792
rect 89682 385736 100708 385792
rect 89621 385734 100708 385736
rect 89621 385731 89687 385734
rect 100702 385732 100708 385734
rect 100772 385732 100778 385796
rect 101949 385794 102015 385797
rect 113265 385794 113331 385797
rect 101949 385792 113331 385794
rect 101949 385736 101954 385792
rect 102010 385736 113270 385792
rect 113326 385736 113331 385792
rect 101949 385734 113331 385736
rect 101949 385731 102015 385734
rect 113265 385731 113331 385734
rect 80881 385658 80947 385661
rect 104157 385658 104223 385661
rect 116117 385658 116183 385661
rect 80881 385656 116183 385658
rect 80881 385600 80886 385656
rect 80942 385600 104162 385656
rect 104218 385600 116122 385656
rect 116178 385600 116183 385656
rect 80881 385598 116183 385600
rect 80881 385595 80947 385598
rect 104157 385595 104223 385598
rect 116117 385595 116183 385598
rect 209589 385658 209655 385661
rect 284385 385658 284451 385661
rect 209589 385656 284451 385658
rect 209589 385600 209594 385656
rect 209650 385600 284390 385656
rect 284446 385600 284451 385656
rect 209589 385598 284451 385600
rect 209589 385595 209655 385598
rect 284385 385595 284451 385598
rect 72417 385114 72483 385117
rect 74758 385114 74764 385116
rect 72417 385112 74764 385114
rect 72417 385056 72422 385112
rect 72478 385056 74764 385112
rect 72417 385054 74764 385056
rect 72417 385051 72483 385054
rect 74758 385052 74764 385054
rect 74828 385052 74834 385116
rect 71681 384978 71747 384981
rect 141969 384978 142035 384981
rect 71681 384976 142035 384978
rect 71681 384920 71686 384976
rect 71742 384920 141974 384976
rect 142030 384920 142035 384976
rect 71681 384918 142035 384920
rect 71681 384915 71747 384918
rect 141969 384915 142035 384918
rect 181529 384978 181595 384981
rect 252461 384978 252527 384981
rect 181529 384976 252527 384978
rect 181529 384920 181534 384976
rect 181590 384920 252466 384976
rect 252522 384920 252527 384976
rect 181529 384918 252527 384920
rect 181529 384915 181595 384918
rect 252461 384915 252527 384918
rect 224861 384842 224927 384845
rect 261109 384842 261175 384845
rect 224861 384840 261175 384842
rect 224861 384784 224866 384840
rect 224922 384784 261114 384840
rect 261170 384784 261175 384840
rect 224861 384782 261175 384784
rect 224861 384779 224927 384782
rect 261109 384779 261175 384782
rect -960 384284 480 384524
rect 141969 384434 142035 384437
rect 188797 384434 188863 384437
rect 199101 384434 199167 384437
rect 141969 384432 199167 384434
rect 141969 384376 141974 384432
rect 142030 384376 188802 384432
rect 188858 384376 199106 384432
rect 199162 384376 199167 384432
rect 141969 384374 199167 384376
rect 141969 384371 142035 384374
rect 188797 384371 188863 384374
rect 199101 384371 199167 384374
rect 91277 384298 91343 384301
rect 162117 384298 162183 384301
rect 91277 384296 162183 384298
rect 91277 384240 91282 384296
rect 91338 384240 162122 384296
rect 162178 384240 162183 384296
rect 91277 384238 162183 384240
rect 91277 384235 91343 384238
rect 161289 383754 161355 383757
rect 161430 383754 161490 384238
rect 162117 384235 162183 384238
rect 186957 384298 187023 384301
rect 220077 384298 220143 384301
rect 186957 384296 220143 384298
rect 186957 384240 186962 384296
rect 187018 384240 220082 384296
rect 220138 384240 220143 384296
rect 186957 384238 220143 384240
rect 186957 384235 187023 384238
rect 220077 384235 220143 384238
rect 180742 383828 180748 383892
rect 180812 383828 180818 383892
rect 180750 383757 180810 383828
rect 180701 383754 180810 383757
rect 161289 383752 161490 383754
rect 161289 383696 161294 383752
rect 161350 383696 161490 383752
rect 161289 383694 161490 383696
rect 180656 383752 180810 383754
rect 180656 383696 180706 383752
rect 180762 383696 180810 383752
rect 180656 383694 180810 383696
rect 161289 383691 161355 383694
rect 180701 383691 180767 383694
rect 67449 383618 67515 383621
rect 128997 383618 129063 383621
rect 180701 383618 180767 383621
rect 180926 383618 180932 383620
rect 67449 383616 129063 383618
rect 67449 383560 67454 383616
rect 67510 383560 129002 383616
rect 129058 383560 129063 383616
rect 67449 383558 129063 383560
rect 180656 383616 180932 383618
rect 180656 383560 180706 383616
rect 180762 383560 180932 383616
rect 180656 383558 180932 383560
rect 67449 383555 67515 383558
rect 128997 383555 129063 383558
rect 180701 383555 180767 383558
rect 180926 383556 180932 383558
rect 180996 383556 181002 383620
rect 188521 383618 188587 383621
rect 265157 383618 265223 383621
rect 188521 383616 265223 383618
rect 188521 383560 188526 383616
rect 188582 383560 265162 383616
rect 265218 383560 265223 383616
rect 188521 383558 265223 383560
rect 188521 383555 188587 383558
rect 265157 383555 265223 383558
rect 171041 383482 171107 383485
rect 216673 383482 216739 383485
rect 171041 383480 216739 383482
rect 171041 383424 171046 383480
rect 171102 383424 216678 383480
rect 216734 383424 216739 383480
rect 171041 383422 216739 383424
rect 171041 383419 171150 383422
rect 216673 383419 216739 383422
rect 93761 382938 93827 382941
rect 102726 382938 102732 382940
rect 93761 382936 102732 382938
rect 93761 382880 93766 382936
rect 93822 382880 102732 382936
rect 93761 382878 102732 382880
rect 93761 382875 93827 382878
rect 102726 382876 102732 382878
rect 102796 382876 102802 382940
rect 103421 382938 103487 382941
rect 114829 382938 114895 382941
rect 103421 382936 114895 382938
rect 103421 382880 103426 382936
rect 103482 382880 114834 382936
rect 114890 382880 114895 382936
rect 103421 382878 114895 382880
rect 103421 382875 103487 382878
rect 114829 382875 114895 382878
rect 160737 382938 160803 382941
rect 171090 382938 171150 383419
rect 160737 382936 171150 382938
rect 160737 382880 160742 382936
rect 160798 382880 171150 382936
rect 160737 382878 171150 382880
rect 232589 382938 232655 382941
rect 242934 382938 242940 382940
rect 232589 382936 242940 382938
rect 232589 382880 232594 382936
rect 232650 382880 242940 382936
rect 232589 382878 242940 382880
rect 160737 382875 160803 382878
rect 232589 382875 232655 382878
rect 242934 382876 242940 382878
rect 243004 382876 243010 382940
rect 265157 382394 265223 382397
rect 265934 382394 265940 382396
rect 265157 382392 265940 382394
rect 265157 382336 265162 382392
rect 265218 382336 265940 382392
rect 265157 382334 265940 382336
rect 265157 382331 265223 382334
rect 265934 382332 265940 382334
rect 266004 382332 266010 382396
rect 106089 382258 106155 382261
rect 243077 382258 243143 382261
rect 274725 382258 274791 382261
rect 106089 382256 274791 382258
rect 106089 382200 106094 382256
rect 106150 382200 243082 382256
rect 243138 382200 274730 382256
rect 274786 382200 274791 382256
rect 106089 382198 274791 382200
rect 106089 382195 106155 382198
rect 243077 382195 243143 382198
rect 274725 382195 274791 382198
rect 99281 382122 99347 382125
rect 170397 382122 170463 382125
rect 99281 382120 170463 382122
rect 99281 382064 99286 382120
rect 99342 382064 170402 382120
rect 170458 382064 170463 382120
rect 99281 382062 170463 382064
rect 99281 382059 99347 382062
rect 170397 382059 170463 382062
rect 186037 382122 186103 382125
rect 220169 382122 220235 382125
rect 186037 382120 220235 382122
rect 186037 382064 186042 382120
rect 186098 382064 220174 382120
rect 220230 382064 220235 382120
rect 186037 382062 220235 382064
rect 186037 382059 186103 382062
rect 220169 382059 220235 382062
rect 181805 381986 181871 381989
rect 215385 381986 215451 381989
rect 181805 381984 215451 381986
rect 181805 381928 181810 381984
rect 181866 381928 215390 381984
rect 215446 381928 215451 381984
rect 181805 381926 215451 381928
rect 181805 381923 181871 381926
rect 215385 381923 215451 381926
rect 240777 381714 240843 381717
rect 258390 381714 258396 381716
rect 240777 381712 258396 381714
rect 240777 381656 240782 381712
rect 240838 381656 258396 381712
rect 240777 381654 258396 381656
rect 240777 381651 240843 381654
rect 258390 381652 258396 381654
rect 258460 381652 258466 381716
rect 231117 381578 231183 381581
rect 265750 381578 265756 381580
rect 231117 381576 265756 381578
rect 231117 381520 231122 381576
rect 231178 381520 265756 381576
rect 231117 381518 265756 381520
rect 231117 381515 231183 381518
rect 265750 381516 265756 381518
rect 265820 381516 265826 381580
rect 215385 381034 215451 381037
rect 215937 381034 216003 381037
rect 215385 381032 216003 381034
rect 215385 380976 215390 381032
rect 215446 380976 215942 381032
rect 215998 380976 216003 381032
rect 215385 380974 216003 380976
rect 215385 380971 215451 380974
rect 215937 380971 216003 380974
rect 243077 381034 243143 381037
rect 244181 381034 244247 381037
rect 243077 381032 244247 381034
rect 243077 380976 243082 381032
rect 243138 380976 244186 381032
rect 244242 380976 244247 381032
rect 243077 380974 244247 380976
rect 243077 380971 243143 380974
rect 244181 380971 244247 380974
rect 3417 380898 3483 380901
rect 120073 380898 120139 380901
rect 3417 380896 120139 380898
rect 3417 380840 3422 380896
rect 3478 380840 120078 380896
rect 120134 380840 120139 380896
rect 3417 380838 120139 380840
rect 3417 380835 3483 380838
rect 120073 380835 120139 380838
rect 189717 380898 189783 380901
rect 281533 380898 281599 380901
rect 189717 380896 281599 380898
rect 189717 380840 189722 380896
rect 189778 380840 281538 380896
rect 281594 380840 281599 380896
rect 189717 380838 281599 380840
rect 189717 380835 189783 380838
rect 281533 380835 281599 380838
rect 108389 380762 108455 380765
rect 180149 380762 180215 380765
rect 108389 380760 180215 380762
rect 108389 380704 108394 380760
rect 108450 380704 180154 380760
rect 180210 380704 180215 380760
rect 108389 380702 180215 380704
rect 108389 380699 108455 380702
rect 180149 380699 180215 380702
rect 186405 380354 186471 380357
rect 220905 380354 220971 380357
rect 186405 380352 220971 380354
rect 186405 380296 186410 380352
rect 186466 380296 220910 380352
rect 220966 380296 220971 380352
rect 186405 380294 220971 380296
rect 186405 380291 186471 380294
rect 220905 380291 220971 380294
rect 155769 380218 155835 380221
rect 189165 380218 189231 380221
rect 155769 380216 189231 380218
rect 155769 380160 155774 380216
rect 155830 380160 189170 380216
rect 189226 380160 189231 380216
rect 155769 380158 189231 380160
rect 155769 380155 155835 380158
rect 189165 380155 189231 380158
rect 108389 379538 108455 379541
rect 108941 379538 109007 379541
rect 108389 379536 109007 379538
rect 108389 379480 108394 379536
rect 108450 379480 108946 379536
rect 109002 379480 109007 379536
rect 108389 379478 109007 379480
rect 108389 379475 108455 379478
rect 108941 379475 109007 379478
rect 88425 379402 88491 379405
rect 123661 379402 123727 379405
rect 88425 379400 123727 379402
rect 88425 379344 88430 379400
rect 88486 379344 123666 379400
rect 123722 379344 123727 379400
rect 88425 379342 123727 379344
rect 88425 379339 88491 379342
rect 123661 379339 123727 379342
rect 173249 379402 173315 379405
rect 276422 379402 276428 379404
rect 173249 379400 276428 379402
rect 173249 379344 173254 379400
rect 173310 379344 276428 379400
rect 173249 379342 276428 379344
rect 173249 379339 173315 379342
rect 276422 379340 276428 379342
rect 276492 379340 276498 379404
rect 154481 378858 154547 378861
rect 206461 378858 206527 378861
rect 154481 378856 206527 378858
rect 154481 378800 154486 378856
rect 154542 378800 206466 378856
rect 206522 378800 206527 378856
rect 154481 378798 206527 378800
rect 154481 378795 154547 378798
rect 206461 378795 206527 378798
rect 106089 378722 106155 378725
rect 117313 378722 117379 378725
rect 106089 378720 117379 378722
rect 106089 378664 106094 378720
rect 106150 378664 117318 378720
rect 117374 378664 117379 378720
rect 106089 378662 117379 378664
rect 106089 378659 106155 378662
rect 117313 378659 117379 378662
rect 123477 378722 123543 378725
rect 187693 378722 187759 378725
rect 123477 378720 187759 378722
rect 123477 378664 123482 378720
rect 123538 378664 187698 378720
rect 187754 378664 187759 378720
rect 123477 378662 187759 378664
rect 123477 378659 123543 378662
rect 187693 378659 187759 378662
rect 247125 378722 247191 378725
rect 254526 378722 254532 378724
rect 247125 378720 254532 378722
rect 247125 378664 247130 378720
rect 247186 378664 254532 378720
rect 247125 378662 254532 378664
rect 247125 378659 247191 378662
rect 254526 378660 254532 378662
rect 254596 378660 254602 378724
rect 582373 378450 582439 378453
rect 583520 378450 584960 378540
rect 582373 378448 584960 378450
rect 582373 378392 582378 378448
rect 582434 378392 584960 378448
rect 582373 378390 584960 378392
rect 582373 378387 582439 378390
rect 583520 378300 584960 378390
rect 67817 378042 67883 378045
rect 152917 378042 152983 378045
rect 67817 378040 152983 378042
rect 67817 377984 67822 378040
rect 67878 377984 152922 378040
rect 152978 377984 152983 378040
rect 67817 377982 152983 377984
rect 67817 377979 67883 377982
rect 152917 377979 152983 377982
rect 187693 378042 187759 378045
rect 287094 378042 287100 378044
rect 187693 378040 287100 378042
rect 187693 377984 187698 378040
rect 187754 377984 287100 378040
rect 187693 377982 287100 377984
rect 187693 377979 187759 377982
rect 287094 377980 287100 377982
rect 287164 377980 287170 378044
rect 152917 377362 152983 377365
rect 162117 377362 162183 377365
rect 152917 377360 162183 377362
rect 152917 377304 152922 377360
rect 152978 377304 162122 377360
rect 162178 377304 162183 377360
rect 152917 377302 162183 377304
rect 152917 377299 152983 377302
rect 162117 377299 162183 377302
rect 234337 377362 234403 377365
rect 258390 377362 258396 377364
rect 234337 377360 258396 377362
rect 234337 377304 234342 377360
rect 234398 377304 258396 377360
rect 234337 377302 258396 377304
rect 234337 377299 234403 377302
rect 258390 377300 258396 377302
rect 258460 377300 258466 377364
rect 122097 376682 122163 376685
rect 267958 376682 267964 376684
rect 122097 376680 267964 376682
rect 122097 376624 122102 376680
rect 122158 376624 267964 376680
rect 122097 376622 267964 376624
rect 122097 376619 122163 376622
rect 267958 376620 267964 376622
rect 268028 376682 268034 376684
rect 268377 376682 268443 376685
rect 268028 376680 268443 376682
rect 268028 376624 268382 376680
rect 268438 376624 268443 376680
rect 268028 376622 268443 376624
rect 268028 376620 268034 376622
rect 268377 376619 268443 376622
rect 86953 376546 87019 376549
rect 144821 376546 144887 376549
rect 186957 376546 187023 376549
rect 86953 376544 187023 376546
rect 86953 376488 86958 376544
rect 87014 376488 144826 376544
rect 144882 376488 186962 376544
rect 187018 376488 187023 376544
rect 86953 376486 187023 376488
rect 86953 376483 87019 376486
rect 144821 376483 144887 376486
rect 186957 376483 187023 376486
rect 65977 376002 66043 376005
rect 80145 376002 80211 376005
rect 65977 376000 80211 376002
rect 65977 375944 65982 376000
rect 66038 375944 80150 376000
rect 80206 375944 80211 376000
rect 65977 375942 80211 375944
rect 65977 375939 66043 375942
rect 80145 375939 80211 375942
rect 229737 376002 229803 376005
rect 270534 376002 270540 376004
rect 229737 376000 270540 376002
rect 229737 375944 229742 376000
rect 229798 375944 270540 376000
rect 229737 375942 270540 375944
rect 229737 375939 229803 375942
rect 270534 375940 270540 375942
rect 270604 375940 270610 376004
rect 188838 375396 188844 375460
rect 188908 375458 188914 375460
rect 190453 375458 190519 375461
rect 188908 375456 190519 375458
rect 188908 375400 190458 375456
rect 190514 375400 190519 375456
rect 188908 375398 190519 375400
rect 188908 375396 188914 375398
rect 190453 375395 190519 375398
rect 142245 375322 142311 375325
rect 142797 375322 142863 375325
rect 186405 375322 186471 375325
rect 142245 375320 186471 375322
rect 142245 375264 142250 375320
rect 142306 375264 142802 375320
rect 142858 375264 186410 375320
rect 186466 375264 186471 375320
rect 142245 375262 186471 375264
rect 142245 375259 142311 375262
rect 142797 375259 142863 375262
rect 186405 375259 186471 375262
rect 239397 375322 239463 375325
rect 291193 375322 291259 375325
rect 239397 375320 291259 375322
rect 239397 375264 239402 375320
rect 239458 375264 291198 375320
rect 291254 375264 291259 375320
rect 239397 375262 291259 375264
rect 239397 375259 239463 375262
rect 291193 375259 291259 375262
rect 181989 375186 182055 375189
rect 208393 375186 208459 375189
rect 181989 375184 208459 375186
rect 181989 375128 181994 375184
rect 182050 375128 208398 375184
rect 208454 375128 208459 375184
rect 181989 375126 208459 375128
rect 181989 375123 182055 375126
rect 208393 375123 208459 375126
rect 232497 374642 232563 374645
rect 249057 374642 249123 374645
rect 232497 374640 249123 374642
rect 232497 374584 232502 374640
rect 232558 374584 249062 374640
rect 249118 374584 249123 374640
rect 232497 374582 249123 374584
rect 232497 374579 232563 374582
rect 249057 374579 249123 374582
rect 180701 374100 180767 374101
rect 180701 374098 180748 374100
rect 180656 374096 180748 374098
rect 180812 374098 180818 374100
rect 180656 374040 180706 374096
rect 180656 374038 180748 374040
rect 180701 374036 180748 374038
rect 180812 374038 180894 374098
rect 180812 374036 180818 374038
rect 180701 374035 180767 374036
rect 180701 373962 180767 373965
rect 182817 373962 182883 373965
rect 249701 373962 249767 373965
rect 180656 373960 180810 373962
rect 180656 373904 180706 373960
rect 180762 373904 180810 373960
rect 180656 373902 180810 373904
rect 180701 373899 180810 373902
rect 182817 373960 249767 373962
rect 182817 373904 182822 373960
rect 182878 373904 249706 373960
rect 249762 373904 249767 373960
rect 182817 373902 249767 373904
rect 182817 373899 182883 373902
rect 249701 373899 249767 373902
rect 180750 373828 180810 373899
rect 180742 373764 180748 373828
rect 180812 373764 180818 373828
rect 220261 373418 220327 373421
rect 241646 373418 241652 373420
rect 220261 373416 241652 373418
rect 220261 373360 220266 373416
rect 220322 373360 241652 373416
rect 220261 373358 241652 373360
rect 220261 373355 220327 373358
rect 241646 373356 241652 373358
rect 241716 373356 241722 373420
rect 235257 373282 235323 373285
rect 260966 373282 260972 373284
rect 235257 373280 260972 373282
rect 235257 373224 235262 373280
rect 235318 373224 260972 373280
rect 235257 373222 260972 373224
rect 235257 373219 235323 373222
rect 260966 373220 260972 373222
rect 261036 373220 261042 373284
rect 187550 372676 187556 372740
rect 187620 372738 187626 372740
rect 190545 372738 190611 372741
rect 187620 372736 190611 372738
rect 187620 372680 190550 372736
rect 190606 372680 190611 372736
rect 187620 372678 190611 372680
rect 187620 372676 187626 372678
rect 190545 372675 190611 372678
rect 107653 372602 107719 372605
rect 247033 372602 247099 372605
rect 107653 372600 247099 372602
rect 107653 372544 107658 372600
rect 107714 372544 247038 372600
rect 247094 372544 247099 372600
rect 107653 372542 247099 372544
rect 107653 372539 107719 372542
rect 247033 372539 247099 372542
rect 161054 371860 161060 371924
rect 161124 371922 161130 371924
rect 164325 371922 164391 371925
rect 161124 371920 164391 371922
rect 161124 371864 164330 371920
rect 164386 371864 164391 371920
rect 161124 371862 164391 371864
rect 161124 371860 161130 371862
rect 164325 371859 164391 371862
rect 227621 371922 227687 371925
rect 262254 371922 262260 371924
rect 227621 371920 262260 371922
rect 227621 371864 227626 371920
rect 227682 371864 262260 371920
rect 227621 371862 262260 371864
rect 227621 371859 227687 371862
rect 262254 371860 262260 371862
rect 262324 371860 262330 371924
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 99281 370698 99347 370701
rect 111006 370698 111012 370700
rect 99281 370696 111012 370698
rect 99281 370640 99286 370696
rect 99342 370640 111012 370696
rect 99281 370638 111012 370640
rect 99281 370635 99347 370638
rect 111006 370636 111012 370638
rect 111076 370636 111082 370700
rect 238109 370698 238175 370701
rect 262305 370698 262371 370701
rect 238109 370696 262371 370698
rect 238109 370640 238114 370696
rect 238170 370640 262310 370696
rect 262366 370640 262371 370696
rect 238109 370638 262371 370640
rect 238109 370635 238175 370638
rect 262305 370635 262371 370638
rect 84101 370562 84167 370565
rect 92790 370562 92796 370564
rect 84101 370560 92796 370562
rect 84101 370504 84106 370560
rect 84162 370504 92796 370560
rect 84101 370502 92796 370504
rect 84101 370499 84167 370502
rect 92790 370500 92796 370502
rect 92860 370500 92866 370564
rect 104801 370562 104867 370565
rect 187693 370562 187759 370565
rect 104801 370560 187759 370562
rect 104801 370504 104806 370560
rect 104862 370504 187698 370560
rect 187754 370504 187759 370560
rect 104801 370502 187759 370504
rect 104801 370499 104867 370502
rect 187693 370499 187759 370502
rect 221457 370562 221523 370565
rect 248454 370562 248460 370564
rect 221457 370560 248460 370562
rect 221457 370504 221462 370560
rect 221518 370504 248460 370560
rect 221457 370502 248460 370504
rect 221457 370499 221523 370502
rect 248454 370500 248460 370502
rect 248524 370500 248530 370564
rect 150249 369746 150315 369749
rect 280245 369748 280311 369749
rect 280245 369746 280292 369748
rect 150249 369744 280292 369746
rect 280356 369746 280362 369748
rect 150249 369688 150254 369744
rect 150310 369688 280250 369744
rect 150249 369686 280292 369688
rect 150249 369683 150315 369686
rect 280245 369684 280292 369686
rect 280356 369686 280438 369746
rect 280356 369684 280362 369686
rect 280245 369683 280311 369684
rect 70393 369066 70459 369069
rect 70894 369066 70900 369068
rect 70393 369064 70900 369066
rect 70393 369008 70398 369064
rect 70454 369008 70900 369064
rect 70393 369006 70900 369008
rect 70393 369003 70459 369006
rect 70894 369004 70900 369006
rect 70964 369066 70970 369068
rect 71681 369066 71747 369069
rect 70964 369064 71747 369066
rect 70964 369008 71686 369064
rect 71742 369008 71747 369064
rect 70964 369006 71747 369008
rect 70964 369004 70970 369006
rect 71681 369003 71747 369006
rect 214649 369066 214715 369069
rect 248638 369066 248644 369068
rect 214649 369064 248644 369066
rect 214649 369008 214654 369064
rect 214710 369008 248644 369064
rect 214649 369006 248644 369008
rect 214649 369003 214715 369006
rect 248638 369004 248644 369006
rect 248708 369004 248714 369068
rect 157977 368386 158043 368389
rect 250437 368386 250503 368389
rect 157977 368384 250503 368386
rect 157977 368328 157982 368384
rect 158038 368328 250442 368384
rect 250498 368328 250503 368384
rect 157977 368326 250503 368328
rect 157977 368323 158043 368326
rect 250437 368323 250503 368326
rect 137461 367026 137527 367029
rect 137737 367026 137803 367029
rect 176653 367026 176719 367029
rect 177389 367026 177455 367029
rect 137461 367024 177455 367026
rect 137461 366968 137466 367024
rect 137522 366968 137742 367024
rect 137798 366968 176658 367024
rect 176714 366968 177394 367024
rect 177450 366968 177455 367024
rect 137461 366966 177455 366968
rect 137461 366963 137527 366966
rect 137737 366963 137803 366966
rect 176653 366963 176719 366966
rect 177389 366963 177455 366966
rect 184841 367026 184907 367029
rect 292573 367026 292639 367029
rect 184841 367024 292639 367026
rect 184841 366968 184846 367024
rect 184902 366968 292578 367024
rect 292634 366968 292639 367024
rect 184841 366966 292639 366968
rect 184841 366963 184907 366966
rect 292573 366963 292639 366966
rect 174629 366346 174695 366349
rect 184841 366346 184907 366349
rect 174629 366344 184907 366346
rect 174629 366288 174634 366344
rect 174690 366288 184846 366344
rect 184902 366288 184907 366344
rect 174629 366286 184907 366288
rect 174629 366283 174695 366286
rect 184841 366283 184907 366286
rect 199377 366346 199443 366349
rect 247217 366346 247283 366349
rect 199377 366344 247283 366346
rect 199377 366288 199382 366344
rect 199438 366288 247222 366344
rect 247278 366288 247283 366344
rect 199377 366286 247283 366288
rect 199377 366283 199443 366286
rect 247217 366283 247283 366286
rect 137277 365666 137343 365669
rect 253933 365666 253999 365669
rect 137277 365664 253999 365666
rect 137277 365608 137282 365664
rect 137338 365608 253938 365664
rect 253994 365608 253999 365664
rect 137277 365606 253999 365608
rect 137277 365603 137343 365606
rect 253933 365603 253999 365606
rect 582465 365122 582531 365125
rect 583520 365122 584960 365212
rect 582465 365120 584960 365122
rect 582465 365064 582470 365120
rect 582526 365064 584960 365120
rect 582465 365062 584960 365064
rect 582465 365059 582531 365062
rect 583520 364972 584960 365062
rect 180701 364444 180767 364445
rect 180701 364442 180748 364444
rect 180656 364440 180748 364442
rect 180812 364442 180818 364444
rect 180656 364384 180706 364440
rect 180656 364382 180748 364384
rect 180701 364380 180748 364382
rect 180812 364382 180894 364442
rect 180812 364380 180818 364382
rect 180701 364379 180767 364380
rect 180701 364306 180767 364309
rect 180656 364304 180810 364306
rect 180656 364248 180706 364304
rect 180762 364248 180810 364304
rect 180656 364246 180810 364248
rect 180701 364243 180810 364246
rect 180750 364172 180810 364243
rect 180742 364108 180748 364172
rect 180812 364108 180818 364172
rect 202137 363626 202203 363629
rect 256693 363626 256759 363629
rect 202137 363624 256759 363626
rect 202137 363568 202142 363624
rect 202198 363568 256698 363624
rect 256754 363568 256759 363624
rect 202137 363566 256759 363568
rect 202137 363563 202203 363566
rect 256693 363563 256759 363566
rect 209037 362266 209103 362269
rect 263726 362266 263732 362268
rect 209037 362264 263732 362266
rect 209037 362208 209042 362264
rect 209098 362208 263732 362264
rect 209037 362206 263732 362208
rect 209037 362203 209103 362206
rect 263726 362204 263732 362206
rect 263796 362204 263802 362268
rect 266629 361722 266695 361725
rect 266854 361722 266860 361724
rect 266629 361720 266860 361722
rect 266629 361664 266634 361720
rect 266690 361664 266860 361720
rect 266629 361662 266860 361664
rect 266629 361659 266695 361662
rect 266854 361660 266860 361662
rect 266924 361660 266930 361724
rect 109033 361586 109099 361589
rect 249609 361586 249675 361589
rect 109033 361584 249675 361586
rect 109033 361528 109038 361584
rect 109094 361528 249614 361584
rect 249670 361528 249675 361584
rect 109033 361526 249675 361528
rect 109033 361523 109099 361526
rect 249609 361523 249675 361526
rect 224217 360906 224283 360909
rect 273478 360906 273484 360908
rect 224217 360904 273484 360906
rect 224217 360848 224222 360904
rect 224278 360848 273484 360904
rect 224217 360846 273484 360848
rect 224217 360843 224283 360846
rect 273478 360844 273484 360846
rect 273548 360844 273554 360908
rect 109033 360226 109099 360229
rect 109677 360226 109743 360229
rect 109033 360224 109743 360226
rect 109033 360168 109038 360224
rect 109094 360168 109682 360224
rect 109738 360168 109743 360224
rect 109033 360166 109743 360168
rect 109033 360163 109099 360166
rect 109677 360163 109743 360166
rect 270769 360226 270835 360229
rect 271086 360226 271092 360228
rect 270769 360224 271092 360226
rect 270769 360168 270774 360224
rect 270830 360168 271092 360224
rect 270769 360166 271092 360168
rect 270769 360163 270835 360166
rect 271086 360164 271092 360166
rect 271156 360164 271162 360228
rect 216673 360090 216739 360093
rect 217409 360090 217475 360093
rect 252502 360090 252508 360092
rect 216673 360088 252508 360090
rect 216673 360032 216678 360088
rect 216734 360032 217414 360088
rect 217470 360032 252508 360088
rect 216673 360030 252508 360032
rect 216673 360027 216739 360030
rect 217409 360027 217475 360030
rect 252502 360028 252508 360030
rect 252572 360028 252578 360092
rect 200757 359410 200823 359413
rect 273294 359410 273300 359412
rect 200757 359408 273300 359410
rect 200757 359352 200762 359408
rect 200818 359352 273300 359408
rect 200757 359350 273300 359352
rect 200757 359347 200823 359350
rect 273294 359348 273300 359350
rect 273364 359348 273370 359412
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 233877 358050 233943 358053
rect 262213 358050 262279 358053
rect 233877 358048 262279 358050
rect 233877 357992 233882 358048
rect 233938 357992 262218 358048
rect 262274 357992 262279 358048
rect 233877 357990 262279 357992
rect 233877 357987 233943 357990
rect 262213 357987 262279 357990
rect 67633 357370 67699 357373
rect 68870 357370 68876 357372
rect 67633 357368 68876 357370
rect 67633 357312 67638 357368
rect 67694 357312 68876 357368
rect 67633 357310 68876 357312
rect 67633 357307 67699 357310
rect 68870 357308 68876 357310
rect 68940 357370 68946 357372
rect 155217 357370 155283 357373
rect 68940 357368 155283 357370
rect 68940 357312 155222 357368
rect 155278 357312 155283 357368
rect 68940 357310 155283 357312
rect 68940 357308 68946 357310
rect 155217 357307 155283 357310
rect 236637 356690 236703 356693
rect 269062 356690 269068 356692
rect 236637 356688 269068 356690
rect 236637 356632 236642 356688
rect 236698 356632 269068 356688
rect 236637 356630 269068 356632
rect 236637 356627 236703 356630
rect 269062 356628 269068 356630
rect 269132 356628 269138 356692
rect 180701 354924 180767 354925
rect 180701 354922 180748 354924
rect 180656 354920 180748 354922
rect 180812 354922 180818 354924
rect 180656 354864 180706 354920
rect 180656 354862 180748 354864
rect 180701 354860 180748 354862
rect 180812 354862 180894 354922
rect 180812 354860 180818 354862
rect 180701 354859 180767 354860
rect 180609 354650 180675 354653
rect 180742 354650 180748 354652
rect 180609 354648 180748 354650
rect 180609 354592 180614 354648
rect 180670 354592 180748 354648
rect 180609 354590 180748 354592
rect 180609 354587 180675 354590
rect 180742 354588 180748 354590
rect 180812 354588 180818 354652
rect 206553 352610 206619 352613
rect 259494 352610 259500 352612
rect 206553 352608 259500 352610
rect 206553 352552 206558 352608
rect 206614 352552 259500 352608
rect 206553 352550 259500 352552
rect 206553 352547 206619 352550
rect 259494 352548 259500 352550
rect 259564 352548 259570 352612
rect 195237 351930 195303 351933
rect 232497 351930 232563 351933
rect 195237 351928 232563 351930
rect 195237 351872 195242 351928
rect 195298 351872 232502 351928
rect 232558 351872 232563 351928
rect 195237 351870 232563 351872
rect 195237 351867 195303 351870
rect 232497 351867 232563 351870
rect 582557 351930 582623 351933
rect 583520 351930 584960 352020
rect 582557 351928 584960 351930
rect 582557 351872 582562 351928
rect 582618 351872 584960 351928
rect 582557 351870 584960 351872
rect 582557 351867 582623 351870
rect 583520 351780 584960 351870
rect 224309 351114 224375 351117
rect 266302 351114 266308 351116
rect 224309 351112 266308 351114
rect 224309 351056 224314 351112
rect 224370 351056 266308 351112
rect 224309 351054 266308 351056
rect 224309 351051 224375 351054
rect 266302 351052 266308 351054
rect 266372 351052 266378 351116
rect 159766 349828 159772 349892
rect 159836 349890 159842 349892
rect 201677 349890 201743 349893
rect 159836 349888 201743 349890
rect 159836 349832 201682 349888
rect 201738 349832 201743 349888
rect 159836 349830 201743 349832
rect 159836 349828 159842 349830
rect 201677 349827 201743 349830
rect 220169 349890 220235 349893
rect 262254 349890 262260 349892
rect 220169 349888 262260 349890
rect 220169 349832 220174 349888
rect 220230 349832 262260 349888
rect 220169 349830 262260 349832
rect 220169 349827 220235 349830
rect 262254 349828 262260 349830
rect 262324 349828 262330 349892
rect 124806 349692 124812 349756
rect 124876 349754 124882 349756
rect 195237 349754 195303 349757
rect 124876 349752 195303 349754
rect 124876 349696 195242 349752
rect 195298 349696 195303 349752
rect 124876 349694 195303 349696
rect 124876 349692 124882 349694
rect 195237 349691 195303 349694
rect 209773 349754 209839 349757
rect 277526 349754 277532 349756
rect 209773 349752 277532 349754
rect 209773 349696 209778 349752
rect 209834 349696 277532 349752
rect 209773 349694 277532 349696
rect 209773 349691 209839 349694
rect 277526 349692 277532 349694
rect 277596 349692 277602 349756
rect 221549 348530 221615 348533
rect 262438 348530 262444 348532
rect 221549 348528 262444 348530
rect 221549 348472 221554 348528
rect 221610 348472 262444 348528
rect 221549 348470 262444 348472
rect 221549 348467 221615 348470
rect 262438 348468 262444 348470
rect 262508 348468 262514 348532
rect 211889 348394 211955 348397
rect 277393 348394 277459 348397
rect 211889 348392 277459 348394
rect 211889 348336 211894 348392
rect 211950 348336 277398 348392
rect 277454 348336 277459 348392
rect 211889 348334 277459 348336
rect 211889 348331 211955 348334
rect 277393 348331 277459 348334
rect 142797 347714 142863 347717
rect 143257 347714 143323 347717
rect 153837 347714 153903 347717
rect 142797 347712 153903 347714
rect 142797 347656 142802 347712
rect 142858 347656 143262 347712
rect 143318 347656 153842 347712
rect 153898 347656 153903 347712
rect 142797 347654 153903 347656
rect 142797 347651 142863 347654
rect 143257 347651 143323 347654
rect 153837 347651 153903 347654
rect 24853 347034 24919 347037
rect 142797 347034 142863 347037
rect 24853 347032 142863 347034
rect 24853 346976 24858 347032
rect 24914 346976 142802 347032
rect 142858 346976 142863 347032
rect 24853 346974 142863 346976
rect 24853 346971 24919 346974
rect 142797 346971 142863 346974
rect 171041 347034 171107 347037
rect 180609 347034 180675 347037
rect 171041 347032 180675 347034
rect 171041 346976 171046 347032
rect 171102 346976 180614 347032
rect 180670 346976 180675 347032
rect 171041 346974 180675 346976
rect 171041 346971 171107 346974
rect 180609 346971 180675 346974
rect 204897 347034 204963 347037
rect 232589 347034 232655 347037
rect 204897 347032 232655 347034
rect 204897 346976 204902 347032
rect 204958 346976 232594 347032
rect 232650 346976 232655 347032
rect 204897 346974 232655 346976
rect 204897 346971 204963 346974
rect 232589 346971 232655 346974
rect 166758 346428 166764 346492
rect 166828 346490 166834 346492
rect 173249 346490 173315 346493
rect 166828 346488 173315 346490
rect 166828 346432 173254 346488
rect 173310 346432 173315 346488
rect 166828 346430 173315 346432
rect 166828 346428 166834 346430
rect 173249 346427 173315 346430
rect 189165 346490 189231 346493
rect 226241 346490 226307 346493
rect 189165 346488 226307 346490
rect 189165 346432 189170 346488
rect 189226 346432 226246 346488
rect 226302 346432 226307 346488
rect 189165 346430 226307 346432
rect 189165 346427 189231 346430
rect 226198 346427 226307 346430
rect 226198 346354 226258 346427
rect 253054 346354 253060 346356
rect 226198 346294 253060 346354
rect 253054 346292 253060 346294
rect 253124 346292 253130 346356
rect 188889 345674 188955 345677
rect 220261 345674 220327 345677
rect 188889 345672 220327 345674
rect 188889 345616 188894 345672
rect 188950 345616 220266 345672
rect 220322 345616 220327 345672
rect 188889 345614 220327 345616
rect 188889 345611 188955 345614
rect 220261 345611 220327 345614
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 166901 344314 166967 344317
rect 244222 344314 244228 344316
rect 166901 344312 244228 344314
rect 166901 344256 166906 344312
rect 166962 344256 244228 344312
rect 166901 344254 244228 344256
rect 166901 344251 166967 344254
rect 244222 344252 244228 344254
rect 244292 344252 244298 344316
rect 179321 343090 179387 343093
rect 202137 343090 202203 343093
rect 179321 343088 202203 343090
rect 179321 343032 179326 343088
rect 179382 343032 202142 343088
rect 202198 343032 202203 343088
rect 179321 343030 202203 343032
rect 179321 343027 179387 343030
rect 202137 343027 202203 343030
rect 191097 342954 191163 342957
rect 238017 342954 238083 342957
rect 191097 342952 238083 342954
rect 191097 342896 191102 342952
rect 191158 342896 238022 342952
rect 238078 342896 238083 342952
rect 191097 342894 238083 342896
rect 191097 342891 191163 342894
rect 238017 342891 238083 342894
rect 169661 341458 169727 341461
rect 178033 341458 178099 341461
rect 169661 341456 178099 341458
rect 169661 341400 169666 341456
rect 169722 341400 178038 341456
rect 178094 341400 178099 341456
rect 169661 341398 178099 341400
rect 169661 341395 169727 341398
rect 178033 341395 178099 341398
rect 180609 341458 180675 341461
rect 231117 341458 231183 341461
rect 180609 341456 231183 341458
rect 180609 341400 180614 341456
rect 180670 341400 231122 341456
rect 231178 341400 231183 341456
rect 180609 341398 231183 341400
rect 180609 341395 180675 341398
rect 231117 341395 231183 341398
rect 177573 340916 177639 340917
rect 177573 340912 177620 340916
rect 177684 340914 177690 340916
rect 177573 340856 177578 340912
rect 177573 340852 177620 340856
rect 177684 340854 177730 340914
rect 177684 340852 177690 340854
rect 177573 340851 177639 340852
rect 177614 340172 177620 340236
rect 177684 340234 177690 340236
rect 207657 340234 207723 340237
rect 177684 340232 207723 340234
rect 177684 340176 207662 340232
rect 207718 340176 207723 340232
rect 177684 340174 207723 340176
rect 177684 340172 177690 340174
rect 207657 340171 207723 340174
rect 196617 340098 196683 340101
rect 278865 340098 278931 340101
rect 196617 340096 278931 340098
rect 196617 340040 196622 340096
rect 196678 340040 278870 340096
rect 278926 340040 278931 340096
rect 196617 340038 278931 340040
rect 196617 340035 196683 340038
rect 278865 340035 278931 340038
rect 240041 339826 240107 339829
rect 245694 339826 245700 339828
rect 240041 339824 245700 339826
rect 240041 339768 240046 339824
rect 240102 339768 245700 339824
rect 240041 339766 245700 339768
rect 240041 339763 240107 339766
rect 245694 339764 245700 339766
rect 245764 339764 245770 339828
rect 81934 339492 81940 339556
rect 82004 339554 82010 339556
rect 82721 339554 82787 339557
rect 82004 339552 82787 339554
rect 82004 339496 82726 339552
rect 82782 339496 82787 339552
rect 82004 339494 82787 339496
rect 82004 339492 82010 339494
rect 82721 339491 82787 339494
rect 148501 338874 148567 338877
rect 177573 338874 177639 338877
rect 207197 338874 207263 338877
rect 148501 338872 207263 338874
rect 148501 338816 148506 338872
rect 148562 338816 177578 338872
rect 177634 338816 207202 338872
rect 207258 338816 207263 338872
rect 148501 338814 207263 338816
rect 148501 338811 148567 338814
rect 177573 338811 177639 338814
rect 207197 338811 207263 338814
rect 20713 338738 20779 338741
rect 158621 338738 158687 338741
rect 201493 338738 201559 338741
rect 20713 338736 201559 338738
rect 20713 338680 20718 338736
rect 20774 338680 158626 338736
rect 158682 338680 201498 338736
rect 201554 338680 201559 338736
rect 20713 338678 201559 338680
rect 20713 338675 20779 338678
rect 158621 338675 158687 338678
rect 201493 338675 201559 338678
rect 224217 338738 224283 338741
rect 263542 338738 263548 338740
rect 224217 338736 263548 338738
rect 224217 338680 224222 338736
rect 224278 338680 263548 338736
rect 224217 338678 263548 338680
rect 224217 338675 224283 338678
rect 263542 338676 263548 338678
rect 263612 338676 263618 338740
rect 583520 338452 584960 338692
rect 219433 338194 219499 338197
rect 202830 338192 219499 338194
rect 202830 338136 219438 338192
rect 219494 338136 219499 338192
rect 202830 338134 219499 338136
rect 153193 338058 153259 338061
rect 158478 338058 158484 338060
rect 153193 338056 158484 338058
rect 153193 338000 153198 338056
rect 153254 338000 158484 338056
rect 153193 337998 158484 338000
rect 153193 337995 153259 337998
rect 158478 337996 158484 337998
rect 158548 338058 158554 338060
rect 202830 338058 202890 338134
rect 219433 338131 219499 338134
rect 158548 337998 202890 338058
rect 205633 338058 205699 338061
rect 206553 338058 206619 338061
rect 205633 338056 206619 338058
rect 205633 338000 205638 338056
rect 205694 338000 206558 338056
rect 206614 338000 206619 338056
rect 205633 337998 206619 338000
rect 158548 337996 158554 337998
rect 205633 337995 205699 337998
rect 206553 337995 206619 337998
rect 223573 338058 223639 338061
rect 224309 338058 224375 338061
rect 223573 338056 224375 338058
rect 223573 338000 223578 338056
rect 223634 338000 224314 338056
rect 224370 338000 224375 338056
rect 223573 337998 224375 338000
rect 223573 337995 223639 337998
rect 224309 337995 224375 337998
rect 178033 337924 178099 337925
rect 177982 337922 177988 337924
rect 177942 337862 177988 337922
rect 178052 337920 178099 337924
rect 178094 337864 178099 337920
rect 177982 337860 177988 337862
rect 178052 337860 178099 337864
rect 178033 337859 178099 337860
rect 128997 337378 129063 337381
rect 178033 337378 178099 337381
rect 223573 337378 223639 337381
rect 128997 337376 161490 337378
rect 128997 337320 129002 337376
rect 129058 337320 161490 337376
rect 128997 337318 161490 337320
rect 128997 337315 129063 337318
rect 161430 337242 161490 337318
rect 178033 337376 223639 337378
rect 178033 337320 178038 337376
rect 178094 337320 223578 337376
rect 223634 337320 223639 337376
rect 178033 337318 223639 337320
rect 178033 337315 178099 337318
rect 223573 337315 223639 337318
rect 178125 337242 178191 337245
rect 178718 337242 178724 337244
rect 161430 337240 178724 337242
rect 161430 337184 178130 337240
rect 178186 337184 178724 337240
rect 161430 337182 178724 337184
rect 178125 337179 178191 337182
rect 178718 337180 178724 337182
rect 178788 337180 178794 337244
rect 144126 336772 144132 336836
rect 144196 336834 144202 336836
rect 205633 336834 205699 336837
rect 144196 336832 205699 336834
rect 144196 336776 205638 336832
rect 205694 336776 205699 336832
rect 144196 336774 205699 336776
rect 144196 336772 144202 336774
rect 205633 336771 205699 336774
rect 220813 336698 220879 336701
rect 221549 336698 221615 336701
rect 220813 336696 221615 336698
rect 220813 336640 220818 336696
rect 220874 336640 221554 336696
rect 221610 336640 221615 336696
rect 220813 336638 221615 336640
rect 220813 336635 220879 336638
rect 221549 336635 221615 336638
rect 126237 336018 126303 336021
rect 190545 336018 190611 336021
rect 215477 336018 215543 336021
rect 126237 336016 215543 336018
rect 126237 335960 126242 336016
rect 126298 335960 190550 336016
rect 190606 335960 215482 336016
rect 215538 335960 215543 336016
rect 126237 335958 215543 335960
rect 126237 335955 126303 335958
rect 190545 335955 190611 335958
rect 215477 335955 215543 335958
rect 217409 336018 217475 336021
rect 266353 336018 266419 336021
rect 217409 336016 266419 336018
rect 217409 335960 217414 336016
rect 217470 335960 266358 336016
rect 266414 335960 266419 336016
rect 217409 335958 266419 335960
rect 217409 335955 217475 335958
rect 266353 335955 266419 335958
rect 17953 335474 18019 335477
rect 220813 335474 220879 335477
rect 17953 335472 220879 335474
rect 17953 335416 17958 335472
rect 18014 335416 220818 335472
rect 220874 335416 220879 335472
rect 17953 335414 220879 335416
rect 17953 335411 18019 335414
rect 220813 335411 220879 335414
rect 154021 334794 154087 334797
rect 172278 334794 172284 334796
rect 154021 334792 172284 334794
rect 154021 334736 154026 334792
rect 154082 334736 172284 334792
rect 154021 334734 172284 334736
rect 154021 334731 154087 334734
rect 172278 334732 172284 334734
rect 172348 334794 172354 334796
rect 202873 334794 202939 334797
rect 172348 334792 202939 334794
rect 172348 334736 202878 334792
rect 202934 334736 202939 334792
rect 172348 334734 202939 334736
rect 172348 334732 172354 334734
rect 202873 334731 202939 334734
rect 134701 334658 134767 334661
rect 178585 334660 178651 334661
rect 178534 334658 178540 334660
rect 134701 334656 178540 334658
rect 178604 334658 178651 334660
rect 204161 334658 204227 334661
rect 226333 334658 226399 334661
rect 178604 334656 178732 334658
rect 134701 334600 134706 334656
rect 134762 334600 178540 334656
rect 178646 334600 178732 334656
rect 134701 334598 178540 334600
rect 134701 334595 134767 334598
rect 178534 334596 178540 334598
rect 178604 334598 178732 334600
rect 204161 334656 226399 334658
rect 204161 334600 204166 334656
rect 204222 334600 226338 334656
rect 226394 334600 226399 334656
rect 204161 334598 226399 334600
rect 178604 334596 178651 334598
rect 178585 334595 178651 334596
rect 204161 334595 204227 334598
rect 226333 334595 226399 334598
rect 244917 334658 244983 334661
rect 263542 334658 263548 334660
rect 244917 334656 263548 334658
rect 244917 334600 244922 334656
rect 244978 334600 263548 334656
rect 244917 334598 263548 334600
rect 244917 334595 244983 334598
rect 263542 334596 263548 334598
rect 263612 334596 263618 334660
rect 22737 334114 22803 334117
rect 200113 334114 200179 334117
rect 200757 334114 200823 334117
rect 22737 334112 200823 334114
rect 22737 334056 22742 334112
rect 22798 334056 200118 334112
rect 200174 334056 200762 334112
rect 200818 334056 200823 334112
rect 22737 334054 200823 334056
rect 22737 334051 22803 334054
rect 200113 334051 200179 334054
rect 200757 334051 200823 334054
rect 137921 333434 137987 333437
rect 150433 333434 150499 333437
rect 137921 333432 150499 333434
rect 137921 333376 137926 333432
rect 137982 333376 150438 333432
rect 150494 333376 150499 333432
rect 137921 333374 150499 333376
rect 137921 333371 137987 333374
rect 150433 333371 150499 333374
rect 11053 333298 11119 333301
rect 169017 333300 169083 333301
rect 168966 333298 168972 333300
rect 11053 333296 168972 333298
rect 169036 333298 169083 333300
rect 188797 333298 188863 333301
rect 258390 333298 258396 333300
rect 169036 333296 169164 333298
rect 11053 333240 11058 333296
rect 11114 333240 168972 333296
rect 169078 333240 169164 333296
rect 11053 333238 168972 333240
rect 11053 333235 11119 333238
rect 168966 333236 168972 333238
rect 169036 333238 169164 333240
rect 188797 333296 258396 333298
rect 188797 333240 188802 333296
rect 188858 333240 258396 333296
rect 188797 333238 258396 333240
rect 169036 333236 169083 333238
rect 169017 333235 169083 333236
rect 188797 333235 188863 333238
rect 258390 333236 258396 333238
rect 258460 333236 258466 333300
rect 150433 332618 150499 332621
rect 230657 332618 230723 332621
rect 150433 332616 230723 332618
rect 150433 332560 150438 332616
rect 150494 332560 230662 332616
rect 230718 332560 230723 332616
rect 150433 332558 230723 332560
rect 150433 332555 150499 332558
rect 230657 332555 230723 332558
rect -960 332196 480 332436
rect 135897 331938 135963 331941
rect 173750 331938 173756 331940
rect 135897 331936 173756 331938
rect 135897 331880 135902 331936
rect 135958 331880 173756 331936
rect 135897 331878 173756 331880
rect 135897 331875 135963 331878
rect 173750 331876 173756 331878
rect 173820 331938 173826 331940
rect 207105 331938 207171 331941
rect 173820 331936 207171 331938
rect 173820 331880 207110 331936
rect 207166 331880 207171 331936
rect 173820 331878 207171 331880
rect 173820 331876 173826 331878
rect 207105 331875 207171 331878
rect 16573 331802 16639 331805
rect 168097 331802 168163 331805
rect 201585 331802 201651 331805
rect 259678 331802 259684 331804
rect 16573 331800 201651 331802
rect 16573 331744 16578 331800
rect 16634 331744 168102 331800
rect 168158 331744 201590 331800
rect 201646 331744 201651 331800
rect 16573 331742 201651 331744
rect 16573 331739 16639 331742
rect 168097 331739 168163 331742
rect 201585 331739 201651 331742
rect 258030 331742 259684 331802
rect 197445 331258 197511 331261
rect 231853 331258 231919 331261
rect 197445 331256 231919 331258
rect 197445 331200 197450 331256
rect 197506 331200 231858 331256
rect 231914 331200 231919 331256
rect 197445 331198 231919 331200
rect 197445 331195 197511 331198
rect 231853 331195 231919 331198
rect 249885 331258 249951 331261
rect 258030 331258 258090 331742
rect 259678 331740 259684 331742
rect 259748 331802 259754 331804
rect 298277 331802 298343 331805
rect 259748 331800 298343 331802
rect 259748 331744 298282 331800
rect 298338 331744 298343 331800
rect 259748 331742 298343 331744
rect 259748 331740 259754 331742
rect 298277 331739 298343 331742
rect 249885 331256 258090 331258
rect 249885 331200 249890 331256
rect 249946 331200 258090 331256
rect 249885 331198 258090 331200
rect 249885 331195 249951 331198
rect 30373 330442 30439 330445
rect 189073 330442 189139 330445
rect 222285 330442 222351 330445
rect 30373 330440 222351 330442
rect 30373 330384 30378 330440
rect 30434 330384 189078 330440
rect 189134 330384 222290 330440
rect 222346 330384 222351 330440
rect 30373 330382 222351 330384
rect 30373 330379 30439 330382
rect 189073 330379 189139 330382
rect 222285 330379 222351 330382
rect 248321 330442 248387 330445
rect 266302 330442 266308 330444
rect 248321 330440 266308 330442
rect 248321 330384 248326 330440
rect 248382 330384 266308 330440
rect 248321 330382 266308 330384
rect 248321 330379 248387 330382
rect 266302 330380 266308 330382
rect 266372 330380 266378 330444
rect 90357 329898 90423 329901
rect 233877 329898 233943 329901
rect 90357 329896 233943 329898
rect 90357 329840 90362 329896
rect 90418 329840 233882 329896
rect 233938 329840 233943 329896
rect 90357 329838 233943 329840
rect 90357 329835 90423 329838
rect 233877 329835 233943 329838
rect 249057 329218 249123 329221
rect 270534 329218 270540 329220
rect 249057 329216 270540 329218
rect 249057 329160 249062 329216
rect 249118 329160 270540 329216
rect 249057 329158 270540 329160
rect 249057 329155 249123 329158
rect 270534 329156 270540 329158
rect 270604 329156 270610 329220
rect 193029 329082 193095 329085
rect 255262 329082 255268 329084
rect 193029 329080 255268 329082
rect 193029 329024 193034 329080
rect 193090 329024 255268 329080
rect 193029 329022 255268 329024
rect 193029 329019 193095 329022
rect 255262 329020 255268 329022
rect 255332 329020 255338 329084
rect 137277 328674 137343 328677
rect 211337 328674 211403 328677
rect 211889 328674 211955 328677
rect 137277 328672 211955 328674
rect 137277 328616 137282 328672
rect 137338 328616 211342 328672
rect 211398 328616 211894 328672
rect 211950 328616 211955 328672
rect 137277 328614 211955 328616
rect 137277 328611 137343 328614
rect 211337 328611 211403 328614
rect 211889 328611 211955 328614
rect 149789 328538 149855 328541
rect 229277 328538 229343 328541
rect 229737 328538 229803 328541
rect 149789 328536 229803 328538
rect 149789 328480 149794 328536
rect 149850 328480 229282 328536
rect 229338 328480 229742 328536
rect 229798 328480 229803 328536
rect 149789 328478 229803 328480
rect 149789 328475 149855 328478
rect 229277 328475 229343 328478
rect 229737 328475 229803 328478
rect 133137 327858 133203 327861
rect 170990 327858 170996 327860
rect 133137 327856 170996 327858
rect 133137 327800 133142 327856
rect 133198 327800 170996 327856
rect 133137 327798 170996 327800
rect 133137 327795 133203 327798
rect 170990 327796 170996 327798
rect 171060 327858 171066 327860
rect 225137 327858 225203 327861
rect 171060 327856 225203 327858
rect 171060 327800 225142 327856
rect 225198 327800 225203 327856
rect 171060 327798 225203 327800
rect 171060 327796 171066 327798
rect 225137 327795 225203 327798
rect 27613 327722 27679 327725
rect 173566 327722 173572 327724
rect 27613 327720 173572 327722
rect 27613 327664 27618 327720
rect 27674 327664 173572 327720
rect 27613 327662 173572 327664
rect 27613 327659 27679 327662
rect 173566 327660 173572 327662
rect 173636 327722 173642 327724
rect 220905 327722 220971 327725
rect 173636 327720 220971 327722
rect 173636 327664 220910 327720
rect 220966 327664 220971 327720
rect 173636 327662 220971 327664
rect 173636 327660 173642 327662
rect 220905 327659 220971 327662
rect 235257 327722 235323 327725
rect 276238 327722 276244 327724
rect 235257 327720 276244 327722
rect 235257 327664 235262 327720
rect 235318 327664 276244 327720
rect 235257 327662 276244 327664
rect 235257 327659 235323 327662
rect 276238 327660 276244 327662
rect 276308 327660 276314 327724
rect 162117 327178 162183 327181
rect 259494 327178 259500 327180
rect 162117 327176 259500 327178
rect 162117 327120 162122 327176
rect 162178 327120 259500 327176
rect 162117 327118 259500 327120
rect 162117 327115 162183 327118
rect 259494 327116 259500 327118
rect 259564 327116 259570 327180
rect 164049 327042 164115 327045
rect 197445 327042 197511 327045
rect 161430 327040 197511 327042
rect 161430 326984 164054 327040
rect 164110 326984 197450 327040
rect 197506 326984 197511 327040
rect 161430 326982 197511 326984
rect 144177 326498 144243 326501
rect 161430 326498 161490 326982
rect 164049 326979 164115 326982
rect 197445 326979 197511 326982
rect 144177 326496 161490 326498
rect 144177 326440 144182 326496
rect 144238 326440 161490 326496
rect 144177 326438 161490 326440
rect 144177 326435 144243 326438
rect 142889 326362 142955 326365
rect 190453 326362 190519 326365
rect 211429 326362 211495 326365
rect 142889 326360 211495 326362
rect 142889 326304 142894 326360
rect 142950 326304 190458 326360
rect 190514 326304 211434 326360
rect 211490 326304 211495 326360
rect 142889 326302 211495 326304
rect 142889 326299 142955 326302
rect 190453 326299 190519 326302
rect 211429 326299 211495 326302
rect 253381 325818 253447 325821
rect 280286 325818 280292 325820
rect 253381 325816 280292 325818
rect 253381 325760 253386 325816
rect 253442 325760 280292 325816
rect 253381 325758 280292 325760
rect 253381 325755 253447 325758
rect 280286 325756 280292 325758
rect 280356 325818 280362 325820
rect 280521 325818 280587 325821
rect 280356 325816 280587 325818
rect 280356 325760 280526 325816
rect 280582 325760 280587 325816
rect 280356 325758 280587 325760
rect 280356 325756 280362 325758
rect 280521 325755 280587 325758
rect 580901 325274 580967 325277
rect 583520 325274 584960 325364
rect 580901 325272 584960 325274
rect 580901 325216 580906 325272
rect 580962 325216 584960 325272
rect 580901 325214 584960 325216
rect 580901 325211 580967 325214
rect 583520 325124 584960 325214
rect 130377 325002 130443 325005
rect 213913 325002 213979 325005
rect 130377 325000 213979 325002
rect 130377 324944 130382 325000
rect 130438 324944 213918 325000
rect 213974 324944 213979 325000
rect 130377 324942 213979 324944
rect 130377 324939 130443 324942
rect 213913 324939 213979 324942
rect 258717 325002 258783 325005
rect 274582 325002 274588 325004
rect 258717 325000 274588 325002
rect 258717 324944 258722 325000
rect 258778 324944 274588 325000
rect 258717 324942 274588 324944
rect 258717 324939 258783 324942
rect 274582 324940 274588 324942
rect 274652 324940 274658 325004
rect 22093 324458 22159 324461
rect 220997 324458 221063 324461
rect 22093 324456 221063 324458
rect 22093 324400 22098 324456
rect 22154 324400 221002 324456
rect 221058 324400 221063 324456
rect 22093 324398 221063 324400
rect 22093 324395 22159 324398
rect 220997 324395 221063 324398
rect 40033 323642 40099 323645
rect 176009 323642 176075 323645
rect 40033 323640 176075 323642
rect 40033 323584 40038 323640
rect 40094 323584 176014 323640
rect 176070 323584 176075 323640
rect 40033 323582 176075 323584
rect 40033 323579 40099 323582
rect 176009 323579 176075 323582
rect 184790 323580 184796 323644
rect 184860 323642 184866 323644
rect 191097 323642 191163 323645
rect 184860 323640 191163 323642
rect 184860 323584 191102 323640
rect 191158 323584 191163 323640
rect 184860 323582 191163 323584
rect 184860 323580 184866 323582
rect 191097 323579 191163 323582
rect 130469 322962 130535 322965
rect 269205 322962 269271 322965
rect 130469 322960 269271 322962
rect 130469 322904 130474 322960
rect 130530 322904 269210 322960
rect 269266 322904 269271 322960
rect 130469 322902 269271 322904
rect 130469 322899 130535 322902
rect 269205 322899 269271 322902
rect 175089 322282 175155 322285
rect 203057 322282 203123 322285
rect 161430 322280 203123 322282
rect 161430 322224 175094 322280
rect 175150 322224 203062 322280
rect 203118 322224 203123 322280
rect 161430 322222 203123 322224
rect 28993 322146 29059 322149
rect 161430 322146 161490 322222
rect 175089 322219 175155 322222
rect 203057 322219 203123 322222
rect 28993 322144 161490 322146
rect 28993 322088 28998 322144
rect 29054 322088 161490 322144
rect 28993 322086 161490 322088
rect 178769 322146 178835 322149
rect 265249 322146 265315 322149
rect 178769 322144 265315 322146
rect 178769 322088 178774 322144
rect 178830 322088 265254 322144
rect 265310 322088 265315 322144
rect 178769 322086 265315 322088
rect 28993 322083 29059 322086
rect 178769 322083 178835 322086
rect 265249 322083 265315 322086
rect 162526 321540 162532 321604
rect 162596 321602 162602 321604
rect 166390 321602 166396 321604
rect 162596 321542 166396 321602
rect 162596 321540 162602 321542
rect 166390 321540 166396 321542
rect 166460 321540 166466 321604
rect 174537 321602 174603 321605
rect 175181 321602 175247 321605
rect 252461 321602 252527 321605
rect 174537 321600 252527 321602
rect 174537 321544 174542 321600
rect 174598 321544 175186 321600
rect 175242 321544 252466 321600
rect 252522 321544 252527 321600
rect 174537 321542 252527 321544
rect 174537 321539 174603 321542
rect 175181 321539 175247 321542
rect 252461 321539 252527 321542
rect 77201 321466 77267 321469
rect 140589 321466 140655 321469
rect 253381 321466 253447 321469
rect 77201 321464 253447 321466
rect 77201 321408 77206 321464
rect 77262 321408 140594 321464
rect 140650 321408 253386 321464
rect 253442 321408 253447 321464
rect 77201 321406 253447 321408
rect 77201 321403 77267 321406
rect 140589 321403 140655 321406
rect 253381 321403 253447 321406
rect 75913 321058 75979 321061
rect 77201 321058 77267 321061
rect 75913 321056 77267 321058
rect 75913 321000 75918 321056
rect 75974 321000 77206 321056
rect 77262 321000 77267 321056
rect 75913 320998 77267 321000
rect 75913 320995 75979 320998
rect 77201 320995 77267 320998
rect 154021 320786 154087 320789
rect 165521 320786 165587 320789
rect 226977 320786 227043 320789
rect 154021 320784 227043 320786
rect 154021 320728 154026 320784
rect 154082 320728 165526 320784
rect 165582 320728 226982 320784
rect 227038 320728 227043 320784
rect 154021 320726 227043 320728
rect 154021 320723 154087 320726
rect 165521 320723 165587 320726
rect 226977 320723 227043 320726
rect 104934 320588 104940 320652
rect 105004 320650 105010 320652
rect 106038 320650 106044 320652
rect 105004 320590 106044 320650
rect 105004 320588 105010 320590
rect 106038 320588 106044 320590
rect 106108 320650 106114 320652
rect 106181 320650 106247 320653
rect 106108 320648 106247 320650
rect 106108 320592 106186 320648
rect 106242 320592 106247 320648
rect 106108 320590 106247 320592
rect 106108 320588 106114 320590
rect 106181 320587 106247 320590
rect 250989 320242 251055 320245
rect 294045 320242 294111 320245
rect 250989 320240 294111 320242
rect 250989 320184 250994 320240
rect 251050 320184 294050 320240
rect 294106 320184 294111 320240
rect 250989 320182 294111 320184
rect 250989 320179 251055 320182
rect 294045 320179 294111 320182
rect 223665 320106 223731 320109
rect 224217 320106 224283 320109
rect 267825 320108 267891 320109
rect 267774 320106 267780 320108
rect 223665 320104 224283 320106
rect 223665 320048 223670 320104
rect 223726 320048 224222 320104
rect 224278 320048 224283 320104
rect 223665 320046 224283 320048
rect 267734 320046 267780 320106
rect 267844 320104 267891 320108
rect 267886 320048 267891 320104
rect 223665 320043 223731 320046
rect 224217 320043 224283 320046
rect 267774 320044 267780 320046
rect 267844 320044 267891 320048
rect 267825 320043 267891 320044
rect -960 319290 480 319380
rect 78438 319364 78444 319428
rect 78508 319426 78514 319428
rect 178677 319426 178743 319429
rect 78508 319424 178743 319426
rect 78508 319368 178682 319424
rect 178738 319368 178743 319424
rect 78508 319366 178743 319368
rect 78508 319364 78514 319366
rect 178677 319363 178743 319366
rect 196709 319426 196775 319429
rect 266445 319426 266511 319429
rect 196709 319424 266511 319426
rect 196709 319368 196714 319424
rect 196770 319368 266450 319424
rect 266506 319368 266511 319424
rect 196709 319366 266511 319368
rect 196709 319363 196775 319366
rect 266445 319363 266511 319366
rect 267774 319364 267780 319428
rect 267844 319426 267850 319428
rect 267917 319426 267983 319429
rect 267844 319424 267983 319426
rect 267844 319368 267922 319424
rect 267978 319368 267983 319424
rect 267844 319366 267983 319368
rect 267844 319364 267850 319366
rect 267917 319363 267983 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 37273 318882 37339 318885
rect 223665 318882 223731 318885
rect 37273 318880 223731 318882
rect 37273 318824 37278 318880
rect 37334 318824 223670 318880
rect 223726 318824 223731 318880
rect 37273 318822 223731 318824
rect 37273 318819 37339 318822
rect 223665 318819 223731 318822
rect 86718 318004 86724 318068
rect 86788 318066 86794 318068
rect 149697 318066 149763 318069
rect 86788 318064 149763 318066
rect 86788 318008 149702 318064
rect 149758 318008 149763 318064
rect 86788 318006 149763 318008
rect 86788 318004 86794 318006
rect 149697 318003 149763 318006
rect 237465 318066 237531 318069
rect 264973 318066 265039 318069
rect 237465 318064 265039 318066
rect 237465 318008 237470 318064
rect 237526 318008 264978 318064
rect 265034 318008 265039 318064
rect 237465 318006 265039 318008
rect 237465 318003 237531 318006
rect 264973 318003 265039 318006
rect 160686 317596 160692 317660
rect 160756 317658 160762 317660
rect 161238 317658 161244 317660
rect 160756 317598 161244 317658
rect 160756 317596 160762 317598
rect 161238 317596 161244 317598
rect 161308 317658 161314 317660
rect 204345 317658 204411 317661
rect 161308 317656 204411 317658
rect 161308 317600 204350 317656
rect 204406 317600 204411 317656
rect 161308 317598 204411 317600
rect 161308 317596 161314 317598
rect 204345 317595 204411 317598
rect 129181 317522 129247 317525
rect 277393 317522 277459 317525
rect 277761 317522 277827 317525
rect 129181 317520 277827 317522
rect 129181 317464 129186 317520
rect 129242 317464 277398 317520
rect 277454 317464 277766 317520
rect 277822 317464 277827 317520
rect 129181 317462 277827 317464
rect 129181 317459 129247 317462
rect 277393 317459 277459 317462
rect 277761 317459 277827 317462
rect 87597 317386 87663 317389
rect 88241 317386 88307 317389
rect 87597 317384 88307 317386
rect 87597 317328 87602 317384
rect 87658 317328 88246 317384
rect 88302 317328 88307 317384
rect 87597 317326 88307 317328
rect 87597 317323 87663 317326
rect 88241 317323 88307 317326
rect 82721 316706 82787 316709
rect 90214 316706 90220 316708
rect 82721 316704 90220 316706
rect 82721 316648 82726 316704
rect 82782 316648 90220 316704
rect 82721 316646 90220 316648
rect 82721 316643 82787 316646
rect 90214 316644 90220 316646
rect 90284 316644 90290 316708
rect 87597 316162 87663 316165
rect 266445 316162 266511 316165
rect 87597 316160 266511 316162
rect 87597 316104 87602 316160
rect 87658 316104 266450 316160
rect 266506 316104 266511 316160
rect 87597 316102 266511 316104
rect 87597 316099 87663 316102
rect 266445 316099 266511 316102
rect 109534 315284 109540 315348
rect 109604 315346 109610 315348
rect 175917 315346 175983 315349
rect 109604 315344 175983 315346
rect 109604 315288 175922 315344
rect 175978 315288 175983 315344
rect 109604 315286 175983 315288
rect 109604 315284 109610 315286
rect 175917 315283 175983 315286
rect 186221 315346 186287 315349
rect 193305 315346 193371 315349
rect 186221 315344 193371 315346
rect 186221 315288 186226 315344
rect 186282 315288 193310 315344
rect 193366 315288 193371 315344
rect 186221 315286 193371 315288
rect 186221 315283 186287 315286
rect 193305 315283 193371 315286
rect 193397 314938 193463 314941
rect 196014 314938 196020 314940
rect 193397 314936 196020 314938
rect 193397 314880 193402 314936
rect 193458 314880 196020 314936
rect 193397 314878 196020 314880
rect 193397 314875 193463 314878
rect 196014 314876 196020 314878
rect 196084 314876 196090 314940
rect 144269 314802 144335 314805
rect 234705 314802 234771 314805
rect 235257 314802 235323 314805
rect 144269 314800 235323 314802
rect 144269 314744 144274 314800
rect 144330 314744 234710 314800
rect 234766 314744 235262 314800
rect 235318 314744 235323 314800
rect 144269 314742 235323 314744
rect 144269 314739 144335 314742
rect 234705 314739 234771 314742
rect 235257 314739 235323 314742
rect 187550 314060 187556 314124
rect 187620 314122 187626 314124
rect 204897 314122 204963 314125
rect 187620 314120 204963 314122
rect 187620 314064 204902 314120
rect 204958 314064 204963 314120
rect 187620 314062 204963 314064
rect 187620 314060 187626 314062
rect 204897 314059 204963 314062
rect 71037 313986 71103 313989
rect 78254 313986 78260 313988
rect 71037 313984 78260 313986
rect 71037 313928 71042 313984
rect 71098 313928 78260 313984
rect 71037 313926 78260 313928
rect 71037 313923 71103 313926
rect 78254 313924 78260 313926
rect 78324 313924 78330 313988
rect 78581 313986 78647 313989
rect 85798 313986 85804 313988
rect 78581 313984 85804 313986
rect 78581 313928 78586 313984
rect 78642 313928 85804 313984
rect 78581 313926 85804 313928
rect 78581 313923 78647 313926
rect 85798 313924 85804 313926
rect 85868 313924 85874 313988
rect 86861 313986 86927 313989
rect 94446 313986 94452 313988
rect 86861 313984 94452 313986
rect 86861 313928 86866 313984
rect 86922 313928 94452 313984
rect 86861 313926 94452 313928
rect 86861 313923 86927 313926
rect 94446 313924 94452 313926
rect 94516 313924 94522 313988
rect 95141 313986 95207 313989
rect 104934 313986 104940 313988
rect 95141 313984 104940 313986
rect 95141 313928 95146 313984
rect 95202 313928 104940 313984
rect 95141 313926 104940 313928
rect 95141 313923 95207 313926
rect 104934 313924 104940 313926
rect 105004 313924 105010 313988
rect 147213 313986 147279 313989
rect 188337 313986 188403 313989
rect 147213 313984 188403 313986
rect 147213 313928 147218 313984
rect 147274 313928 188342 313984
rect 188398 313928 188403 313984
rect 147213 313926 188403 313928
rect 147213 313923 147279 313926
rect 188337 313923 188403 313926
rect 209313 313986 209379 313989
rect 282913 313986 282979 313989
rect 209313 313984 282979 313986
rect 209313 313928 209318 313984
rect 209374 313928 282918 313984
rect 282974 313928 282979 313984
rect 209313 313926 282979 313928
rect 209313 313923 209379 313926
rect 282913 313923 282979 313926
rect 140037 313306 140103 313309
rect 208393 313306 208459 313309
rect 209313 313306 209379 313309
rect 140037 313304 209379 313306
rect 140037 313248 140042 313304
rect 140098 313248 208398 313304
rect 208454 313248 209318 313304
rect 209374 313248 209379 313304
rect 140037 313246 209379 313248
rect 140037 313243 140103 313246
rect 208393 313243 208459 313246
rect 209313 313243 209379 313246
rect 91001 312490 91067 312493
rect 98494 312490 98500 312492
rect 91001 312488 98500 312490
rect 91001 312432 91006 312488
rect 91062 312432 98500 312488
rect 91001 312430 98500 312432
rect 91001 312427 91067 312430
rect 98494 312428 98500 312430
rect 98564 312428 98570 312492
rect 183461 312490 183527 312493
rect 197997 312490 198063 312493
rect 183461 312488 198063 312490
rect 183461 312432 183466 312488
rect 183522 312432 198002 312488
rect 198058 312432 198063 312488
rect 183461 312430 198063 312432
rect 183461 312427 183527 312430
rect 197997 312427 198063 312430
rect 223481 312490 223547 312493
rect 269481 312490 269547 312493
rect 223481 312488 269547 312490
rect 223481 312432 223486 312488
rect 223542 312432 269486 312488
rect 269542 312432 269547 312488
rect 223481 312430 269547 312432
rect 223481 312427 223547 312430
rect 269481 312427 269547 312430
rect 582649 312082 582715 312085
rect 583520 312082 584960 312172
rect 582649 312080 584960 312082
rect 582649 312024 582654 312080
rect 582710 312024 584960 312080
rect 582649 312022 584960 312024
rect 582649 312019 582715 312022
rect 92473 311946 92539 311949
rect 270769 311946 270835 311949
rect 92473 311944 270835 311946
rect 92473 311888 92478 311944
rect 92534 311888 270774 311944
rect 270830 311888 270835 311944
rect 583520 311932 584960 312022
rect 92473 311886 270835 311888
rect 92473 311883 92539 311886
rect 270769 311883 270835 311886
rect 218697 311810 218763 311813
rect 248689 311810 248755 311813
rect 249609 311810 249675 311813
rect 218697 311808 249675 311810
rect 218697 311752 218702 311808
rect 218758 311752 248694 311808
rect 248750 311752 249614 311808
rect 249670 311752 249675 311808
rect 218697 311750 249675 311752
rect 218697 311747 218763 311750
rect 248689 311747 248755 311750
rect 249609 311747 249675 311750
rect 87454 311204 87460 311268
rect 87524 311266 87530 311268
rect 89713 311266 89779 311269
rect 87524 311264 89779 311266
rect 87524 311208 89718 311264
rect 89774 311208 89779 311264
rect 87524 311206 89779 311208
rect 87524 311204 87530 311206
rect 89713 311203 89779 311206
rect 253197 311266 253263 311269
rect 256734 311266 256740 311268
rect 253197 311264 256740 311266
rect 253197 311208 253202 311264
rect 253258 311208 256740 311264
rect 253197 311206 256740 311208
rect 253197 311203 253263 311206
rect 256734 311204 256740 311206
rect 256804 311204 256810 311268
rect 79961 311130 80027 311133
rect 87086 311130 87092 311132
rect 79961 311128 87092 311130
rect 79961 311072 79966 311128
rect 80022 311072 87092 311128
rect 79961 311070 87092 311072
rect 79961 311067 80027 311070
rect 87086 311068 87092 311070
rect 87156 311068 87162 311132
rect 94497 311130 94563 311133
rect 106406 311130 106412 311132
rect 94497 311128 106412 311130
rect 94497 311072 94502 311128
rect 94558 311072 106412 311128
rect 94497 311070 106412 311072
rect 94497 311067 94563 311070
rect 106406 311068 106412 311070
rect 106476 311068 106482 311132
rect 190269 311130 190335 311133
rect 209129 311130 209195 311133
rect 190269 311128 209195 311130
rect 190269 311072 190274 311128
rect 190330 311072 209134 311128
rect 209190 311072 209195 311128
rect 190269 311070 209195 311072
rect 190269 311067 190335 311070
rect 209129 311067 209195 311070
rect 222837 311130 222903 311133
rect 253381 311130 253447 311133
rect 222837 311128 253447 311130
rect 222837 311072 222842 311128
rect 222898 311072 253386 311128
rect 253442 311072 253447 311128
rect 222837 311070 253447 311072
rect 222837 311067 222903 311070
rect 253381 311067 253447 311070
rect 248597 310994 248663 310997
rect 249701 310994 249767 310997
rect 248597 310992 249767 310994
rect 248597 310936 248602 310992
rect 248658 310936 249706 310992
rect 249762 310936 249767 310992
rect 248597 310934 249767 310936
rect 248597 310931 248663 310934
rect 249701 310931 249767 310934
rect 147029 310722 147095 310725
rect 196617 310722 196683 310725
rect 147029 310720 196683 310722
rect 147029 310664 147034 310720
rect 147090 310664 196622 310720
rect 196678 310664 196683 310720
rect 147029 310662 196683 310664
rect 147029 310659 147095 310662
rect 196617 310659 196683 310662
rect 187693 310586 187759 310589
rect 237465 310586 237531 310589
rect 187693 310584 237531 310586
rect 187693 310528 187698 310584
rect 187754 310528 237470 310584
rect 237526 310528 237531 310584
rect 187693 310526 237531 310528
rect 187693 310523 187759 310526
rect 237465 310523 237531 310526
rect 249701 310586 249767 310589
rect 295425 310586 295491 310589
rect 249701 310584 295491 310586
rect 249701 310528 249706 310584
rect 249762 310528 295430 310584
rect 295486 310528 295491 310584
rect 249701 310526 295491 310528
rect 249701 310523 249767 310526
rect 295425 310523 295491 310526
rect 148174 310388 148180 310452
rect 148244 310450 148250 310452
rect 153837 310450 153903 310453
rect 148244 310448 153903 310450
rect 148244 310392 153842 310448
rect 153898 310392 153903 310448
rect 148244 310390 153903 310392
rect 148244 310388 148250 310390
rect 153837 310387 153903 310390
rect 244365 310450 244431 310453
rect 245009 310450 245075 310453
rect 244365 310448 245075 310450
rect 244365 310392 244370 310448
rect 244426 310392 245014 310448
rect 245070 310392 245075 310448
rect 244365 310390 245075 310392
rect 244365 310387 244431 310390
rect 245009 310387 245075 310390
rect 124949 309770 125015 309773
rect 187693 309770 187759 309773
rect 124949 309768 187759 309770
rect 124949 309712 124954 309768
rect 125010 309712 187698 309768
rect 187754 309712 187759 309768
rect 124949 309710 187759 309712
rect 124949 309707 125015 309710
rect 187693 309707 187759 309710
rect 212441 309770 212507 309773
rect 267825 309770 267891 309773
rect 212441 309768 267891 309770
rect 212441 309712 212446 309768
rect 212502 309712 267830 309768
rect 267886 309712 267891 309768
rect 212441 309710 267891 309712
rect 212441 309707 212507 309710
rect 267825 309707 267891 309710
rect 173014 309300 173020 309364
rect 173084 309362 173090 309364
rect 210233 309362 210299 309365
rect 210417 309362 210483 309365
rect 173084 309360 210483 309362
rect 173084 309304 210238 309360
rect 210294 309304 210422 309360
rect 210478 309304 210483 309360
rect 173084 309302 210483 309304
rect 173084 309300 173090 309302
rect 210233 309299 210299 309302
rect 210417 309299 210483 309302
rect 184197 309226 184263 309229
rect 231117 309226 231183 309229
rect 184197 309224 231183 309226
rect 184197 309168 184202 309224
rect 184258 309168 231122 309224
rect 231178 309168 231183 309224
rect 184197 309166 231183 309168
rect 184197 309163 184263 309166
rect 231117 309163 231183 309166
rect 244365 309226 244431 309229
rect 295333 309226 295399 309229
rect 244365 309224 295399 309226
rect 244365 309168 244370 309224
rect 244426 309168 295338 309224
rect 295394 309168 295399 309224
rect 244365 309166 295399 309168
rect 244365 309163 244431 309166
rect 295333 309163 295399 309166
rect 194542 309028 194548 309092
rect 194612 309090 194618 309092
rect 195053 309090 195119 309093
rect 194612 309088 195119 309090
rect 194612 309032 195058 309088
rect 195114 309032 195119 309088
rect 194612 309030 195119 309032
rect 194612 309028 194618 309030
rect 195053 309027 195119 309030
rect 88241 308546 88307 308549
rect 97942 308546 97948 308548
rect 88241 308544 97948 308546
rect 88241 308488 88246 308544
rect 88302 308488 97948 308544
rect 88241 308486 97948 308488
rect 88241 308483 88307 308486
rect 97942 308484 97948 308486
rect 98012 308484 98018 308548
rect 52269 308410 52335 308413
rect 281574 308410 281580 308412
rect 52269 308408 281580 308410
rect 52269 308352 52274 308408
rect 52330 308352 281580 308408
rect 52269 308350 281580 308352
rect 52269 308347 52335 308350
rect 281574 308348 281580 308350
rect 281644 308348 281650 308412
rect 188337 308002 188403 308005
rect 220169 308002 220235 308005
rect 188337 308000 220235 308002
rect 188337 307944 188342 308000
rect 188398 307944 220174 308000
rect 220230 307944 220235 308000
rect 188337 307942 220235 307944
rect 188337 307939 188403 307942
rect 220169 307939 220235 307942
rect 138657 307866 138723 307869
rect 195053 307866 195119 307869
rect 138657 307864 195119 307866
rect 138657 307808 138662 307864
rect 138718 307808 195058 307864
rect 195114 307808 195119 307864
rect 138657 307806 195119 307808
rect 138657 307803 138723 307806
rect 195053 307803 195119 307806
rect 247677 307866 247743 307869
rect 299657 307866 299723 307869
rect 247677 307864 299723 307866
rect 247677 307808 247682 307864
rect 247738 307808 299662 307864
rect 299718 307808 299723 307864
rect 247677 307806 299723 307808
rect 247677 307803 247743 307806
rect 299657 307803 299723 307806
rect 70301 307730 70367 307733
rect 71078 307730 71084 307732
rect 70301 307728 71084 307730
rect 70301 307672 70306 307728
rect 70362 307672 71084 307728
rect 70301 307670 71084 307672
rect 70301 307667 70367 307670
rect 71078 307668 71084 307670
rect 71148 307668 71154 307732
rect 86534 307668 86540 307732
rect 86604 307730 86610 307732
rect 91369 307730 91435 307733
rect 86604 307728 91435 307730
rect 86604 307672 91374 307728
rect 91430 307672 91435 307728
rect 86604 307670 91435 307672
rect 86604 307668 86610 307670
rect 91369 307667 91435 307670
rect 240133 307730 240199 307733
rect 241237 307730 241303 307733
rect 240133 307728 241303 307730
rect 240133 307672 240138 307728
rect 240194 307672 241242 307728
rect 241298 307672 241303 307728
rect 240133 307670 241303 307672
rect 240133 307667 240199 307670
rect 241237 307667 241303 307670
rect 269614 307668 269620 307732
rect 269684 307730 269690 307732
rect 270493 307730 270559 307733
rect 269684 307728 270559 307730
rect 269684 307672 270498 307728
rect 270554 307672 270559 307728
rect 269684 307670 270559 307672
rect 269684 307668 269690 307670
rect 270493 307667 270559 307670
rect 95325 307050 95391 307053
rect 109534 307050 109540 307052
rect 95325 307048 109540 307050
rect 95325 306992 95330 307048
rect 95386 306992 109540 307048
rect 95325 306990 109540 306992
rect 95325 306987 95391 306990
rect 109534 306988 109540 306990
rect 109604 306988 109610 307052
rect 218053 307050 218119 307053
rect 246205 307050 246271 307053
rect 218053 307048 246271 307050
rect 218053 306992 218058 307048
rect 218114 306992 246210 307048
rect 246266 306992 246271 307048
rect 218053 306990 246271 306992
rect 218053 306987 218119 306990
rect 246205 306987 246271 306990
rect 246389 307050 246455 307053
rect 260966 307050 260972 307052
rect 246389 307048 260972 307050
rect 246389 306992 246394 307048
rect 246450 306992 260972 307048
rect 246389 306990 260972 306992
rect 246389 306987 246455 306990
rect 260966 306988 260972 306990
rect 261036 306988 261042 307052
rect 185342 306716 185348 306780
rect 185412 306778 185418 306780
rect 223389 306778 223455 306781
rect 185412 306776 223455 306778
rect 185412 306720 223394 306776
rect 223450 306720 223455 306776
rect 185412 306718 223455 306720
rect 185412 306716 185418 306718
rect 223389 306715 223455 306718
rect 77293 306642 77359 306645
rect 86166 306642 86172 306644
rect 77293 306640 86172 306642
rect 77293 306584 77298 306640
rect 77354 306584 86172 306640
rect 77293 306582 86172 306584
rect 77293 306579 77359 306582
rect 86166 306580 86172 306582
rect 86236 306580 86242 306644
rect 149697 306642 149763 306645
rect 209037 306642 209103 306645
rect 149697 306640 209103 306642
rect 149697 306584 149702 306640
rect 149758 306584 209042 306640
rect 209098 306584 209103 306640
rect 149697 306582 209103 306584
rect 149697 306579 149763 306582
rect 209037 306579 209103 306582
rect 5533 306506 5599 306509
rect 176745 306506 176811 306509
rect 5533 306504 176811 306506
rect 5533 306448 5538 306504
rect 5594 306448 176750 306504
rect 176806 306448 176811 306504
rect 5533 306446 176811 306448
rect 5533 306443 5599 306446
rect 176745 306443 176811 306446
rect 185577 306506 185643 306509
rect 241237 306506 241303 306509
rect 185577 306504 241303 306506
rect 185577 306448 185582 306504
rect 185638 306448 241242 306504
rect 241298 306448 241303 306504
rect 185577 306446 241303 306448
rect 185577 306443 185643 306446
rect 241237 306443 241303 306446
rect 245561 306506 245627 306509
rect 277577 306506 277643 306509
rect 245561 306504 277643 306506
rect 245561 306448 245566 306504
rect 245622 306448 277582 306504
rect 277638 306448 277643 306504
rect 245561 306446 277643 306448
rect 245561 306443 245627 306446
rect 277577 306443 277643 306446
rect -960 306234 480 306324
rect 156638 306308 156644 306372
rect 156708 306370 156714 306372
rect 188337 306370 188403 306373
rect 156708 306368 188403 306370
rect 156708 306312 188342 306368
rect 188398 306312 188403 306368
rect 156708 306310 188403 306312
rect 156708 306308 156714 306310
rect 188337 306307 188403 306310
rect 199193 306370 199259 306373
rect 199377 306370 199443 306373
rect 199193 306368 199443 306370
rect 199193 306312 199198 306368
rect 199254 306312 199382 306368
rect 199438 306312 199443 306368
rect 199193 306310 199443 306312
rect 199193 306307 199259 306310
rect 199377 306307 199443 306310
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 244457 305826 244523 305829
rect 273294 305826 273300 305828
rect 244457 305824 273300 305826
rect 244457 305768 244462 305824
rect 244518 305768 273300 305824
rect 244457 305766 273300 305768
rect 244457 305763 244523 305766
rect 273294 305764 273300 305766
rect 273364 305764 273370 305828
rect 145649 305690 145715 305693
rect 164141 305690 164207 305693
rect 194409 305690 194475 305693
rect 145649 305688 194475 305690
rect 145649 305632 145654 305688
rect 145710 305632 164146 305688
rect 164202 305632 194414 305688
rect 194470 305632 194475 305688
rect 145649 305630 194475 305632
rect 145649 305627 145715 305630
rect 164141 305627 164207 305630
rect 194409 305627 194475 305630
rect 218697 305690 218763 305693
rect 245694 305690 245700 305692
rect 218697 305688 245700 305690
rect 218697 305632 218702 305688
rect 218758 305632 245700 305688
rect 218697 305630 245700 305632
rect 218697 305627 218763 305630
rect 245694 305628 245700 305630
rect 245764 305628 245770 305692
rect 262438 305690 262444 305692
rect 258030 305630 262444 305690
rect 184657 305282 184723 305285
rect 258030 305282 258090 305630
rect 262438 305628 262444 305630
rect 262508 305690 262514 305692
rect 299565 305690 299631 305693
rect 262508 305688 299631 305690
rect 262508 305632 299570 305688
rect 299626 305632 299631 305688
rect 262508 305630 299631 305632
rect 262508 305628 262514 305630
rect 299565 305627 299631 305630
rect 184657 305280 258090 305282
rect 184657 305224 184662 305280
rect 184718 305224 258090 305280
rect 184657 305222 258090 305224
rect 184657 305219 184723 305222
rect 188337 305146 188403 305149
rect 205817 305146 205883 305149
rect 206277 305146 206343 305149
rect 188337 305144 206343 305146
rect 188337 305088 188342 305144
rect 188398 305088 205822 305144
rect 205878 305088 206282 305144
rect 206338 305088 206343 305144
rect 188337 305086 206343 305088
rect 188337 305083 188403 305086
rect 205817 305083 205883 305086
rect 206277 305083 206343 305086
rect 241789 305010 241855 305013
rect 244457 305010 244523 305013
rect 241789 305008 244523 305010
rect 241789 304952 241794 305008
rect 241850 304952 244462 305008
rect 244518 304952 244523 305008
rect 241789 304950 244523 304952
rect 241789 304947 241855 304950
rect 244457 304947 244523 304950
rect 86769 304330 86835 304333
rect 95182 304330 95188 304332
rect 86769 304328 95188 304330
rect 86769 304272 86774 304328
rect 86830 304272 95188 304328
rect 86769 304270 95188 304272
rect 86769 304267 86835 304270
rect 95182 304268 95188 304270
rect 95252 304268 95258 304332
rect 246941 304330 247007 304333
rect 252553 304330 252619 304333
rect 246941 304328 252619 304330
rect 246941 304272 246946 304328
rect 247002 304272 252558 304328
rect 252614 304272 252619 304328
rect 246941 304270 252619 304272
rect 246941 304267 247007 304270
rect 252553 304267 252619 304270
rect 69197 304194 69263 304197
rect 75862 304194 75868 304196
rect 69197 304192 75868 304194
rect 69197 304136 69202 304192
rect 69258 304136 75868 304192
rect 69197 304134 75868 304136
rect 69197 304131 69263 304134
rect 75862 304132 75868 304134
rect 75932 304132 75938 304196
rect 84009 304194 84075 304197
rect 92974 304194 92980 304196
rect 84009 304192 92980 304194
rect 84009 304136 84014 304192
rect 84070 304136 92980 304192
rect 84009 304134 92980 304136
rect 84009 304131 84075 304134
rect 92974 304132 92980 304134
rect 93044 304132 93050 304196
rect 101397 304194 101463 304197
rect 113214 304194 113220 304196
rect 101397 304192 113220 304194
rect 101397 304136 101402 304192
rect 101458 304136 113220 304192
rect 101397 304134 113220 304136
rect 101397 304131 101463 304134
rect 113214 304132 113220 304134
rect 113284 304132 113290 304196
rect 141417 304194 141483 304197
rect 180558 304194 180564 304196
rect 141417 304192 180564 304194
rect 141417 304136 141422 304192
rect 141478 304136 180564 304192
rect 141417 304134 180564 304136
rect 141417 304131 141483 304134
rect 180558 304132 180564 304134
rect 180628 304194 180634 304196
rect 214833 304194 214899 304197
rect 180628 304192 214899 304194
rect 180628 304136 214838 304192
rect 214894 304136 214899 304192
rect 180628 304134 214899 304136
rect 180628 304132 180634 304134
rect 214833 304131 214899 304134
rect 247217 304194 247283 304197
rect 277158 304194 277164 304196
rect 247217 304192 277164 304194
rect 247217 304136 247222 304192
rect 247278 304136 277164 304192
rect 247217 304134 277164 304136
rect 247217 304131 247283 304134
rect 277158 304132 277164 304134
rect 277228 304194 277234 304196
rect 281809 304194 281875 304197
rect 277228 304192 281875 304194
rect 277228 304136 281814 304192
rect 281870 304136 281875 304192
rect 277228 304134 281875 304136
rect 277228 304132 277234 304134
rect 281809 304131 281875 304134
rect 240041 303922 240107 303925
rect 269113 303922 269179 303925
rect 240041 303920 269179 303922
rect 240041 303864 240046 303920
rect 240102 303864 269118 303920
rect 269174 303864 269179 303920
rect 240041 303862 269179 303864
rect 240041 303859 240107 303862
rect 269113 303859 269179 303862
rect 188470 303724 188476 303788
rect 188540 303786 188546 303788
rect 194593 303786 194659 303789
rect 195605 303786 195671 303789
rect 188540 303784 195671 303786
rect 188540 303728 194598 303784
rect 194654 303728 195610 303784
rect 195666 303728 195671 303784
rect 188540 303726 195671 303728
rect 188540 303724 188546 303726
rect 194593 303723 194659 303726
rect 195605 303723 195671 303726
rect 252553 303786 252619 303789
rect 263726 303786 263732 303788
rect 252553 303784 263732 303786
rect 252553 303728 252558 303784
rect 252614 303728 263732 303784
rect 252553 303726 263732 303728
rect 252553 303723 252619 303726
rect 263726 303724 263732 303726
rect 263796 303724 263802 303788
rect 66110 303588 66116 303652
rect 66180 303650 66186 303652
rect 69657 303650 69723 303653
rect 66180 303648 69723 303650
rect 66180 303592 69662 303648
rect 69718 303592 69723 303648
rect 66180 303590 69723 303592
rect 66180 303588 66186 303590
rect 69657 303587 69723 303590
rect 76557 303650 76623 303653
rect 83038 303650 83044 303652
rect 76557 303648 83044 303650
rect 76557 303592 76562 303648
rect 76618 303592 83044 303648
rect 76557 303590 83044 303592
rect 76557 303587 76623 303590
rect 83038 303588 83044 303590
rect 83108 303588 83114 303652
rect 186814 303588 186820 303652
rect 186884 303650 186890 303652
rect 201677 303650 201743 303653
rect 202781 303650 202847 303653
rect 186884 303648 202847 303650
rect 186884 303592 201682 303648
rect 201738 303592 202786 303648
rect 202842 303592 202847 303648
rect 186884 303590 202847 303592
rect 186884 303588 186890 303590
rect 201677 303587 201743 303590
rect 202781 303587 202847 303590
rect 211061 303650 211127 303653
rect 232221 303650 232287 303653
rect 211061 303648 232287 303650
rect 211061 303592 211066 303648
rect 211122 303592 232226 303648
rect 232282 303592 232287 303648
rect 211061 303590 232287 303592
rect 211061 303587 211127 303590
rect 232221 303587 232287 303590
rect 158529 303514 158595 303517
rect 163681 303514 163747 303517
rect 158529 303512 163747 303514
rect 158529 303456 158534 303512
rect 158590 303456 163686 303512
rect 163742 303456 163747 303512
rect 158529 303454 163747 303456
rect 158529 303451 158595 303454
rect 163681 303451 163747 303454
rect 184054 302500 184060 302564
rect 184124 302562 184130 302564
rect 212441 302562 212507 302565
rect 184124 302560 212507 302562
rect 184124 302504 212446 302560
rect 212502 302504 212507 302560
rect 184124 302502 212507 302504
rect 184124 302500 184130 302502
rect 212441 302499 212507 302502
rect 105537 302426 105603 302429
rect 241421 302426 241487 302429
rect 250161 302426 250227 302429
rect 105537 302424 250227 302426
rect 105537 302368 105542 302424
rect 105598 302368 241426 302424
rect 241482 302368 250166 302424
rect 250222 302368 250227 302424
rect 105537 302366 250227 302368
rect 105537 302363 105603 302366
rect 241421 302363 241487 302366
rect 250161 302363 250227 302366
rect 252001 302426 252067 302429
rect 285765 302426 285831 302429
rect 252001 302424 285831 302426
rect 252001 302368 252006 302424
rect 252062 302368 285770 302424
rect 285826 302368 285831 302424
rect 252001 302366 285831 302368
rect 252001 302363 252067 302366
rect 285765 302363 285831 302366
rect 179321 302292 179387 302293
rect 179270 302290 179276 302292
rect 179230 302230 179276 302290
rect 179340 302288 179387 302292
rect 223481 302290 223547 302293
rect 179382 302232 179387 302288
rect 179270 302228 179276 302230
rect 179340 302228 179387 302232
rect 179321 302227 179387 302228
rect 179462 302288 223547 302290
rect 179462 302232 223486 302288
rect 223542 302232 223547 302288
rect 179462 302230 223547 302232
rect 179321 302154 179387 302157
rect 179462 302154 179522 302230
rect 223481 302227 223547 302230
rect 238845 302290 238911 302293
rect 582373 302290 582439 302293
rect 238845 302288 582439 302290
rect 238845 302232 238850 302288
rect 238906 302232 582378 302288
rect 582434 302232 582439 302288
rect 238845 302230 582439 302232
rect 238845 302227 238911 302230
rect 582373 302227 582439 302230
rect 179321 302152 179522 302154
rect 179321 302096 179326 302152
rect 179382 302096 179522 302152
rect 179321 302094 179522 302096
rect 239397 302154 239463 302157
rect 246297 302154 246363 302157
rect 239397 302152 246363 302154
rect 239397 302096 239402 302152
rect 239458 302096 246302 302152
rect 246358 302096 246363 302152
rect 239397 302094 246363 302096
rect 179321 302091 179387 302094
rect 239397 302091 239463 302094
rect 246297 302091 246363 302094
rect 142797 301746 142863 301749
rect 166257 301748 166323 301749
rect 166206 301746 166212 301748
rect 142797 301744 166212 301746
rect 166276 301744 166323 301748
rect 234521 301746 234587 301749
rect 142797 301688 142802 301744
rect 142858 301688 166212 301744
rect 166318 301688 166323 301744
rect 142797 301686 166212 301688
rect 142797 301683 142863 301686
rect 166206 301684 166212 301686
rect 166276 301684 166323 301688
rect 166257 301683 166323 301684
rect 234478 301744 234587 301746
rect 234478 301688 234526 301744
rect 234582 301688 234587 301744
rect 234478 301683 234587 301688
rect 251817 301746 251883 301749
rect 254577 301746 254643 301749
rect 251817 301744 254643 301746
rect 251817 301688 251822 301744
rect 251878 301688 254582 301744
rect 254638 301688 254643 301744
rect 251817 301686 254643 301688
rect 251817 301683 251883 301686
rect 254577 301683 254643 301686
rect 159766 301548 159772 301612
rect 159836 301610 159842 301612
rect 160001 301610 160067 301613
rect 216857 301610 216923 301613
rect 159836 301608 216923 301610
rect 159836 301552 160006 301608
rect 160062 301552 216862 301608
rect 216918 301552 216923 301608
rect 159836 301550 216923 301552
rect 159836 301548 159842 301550
rect 160001 301547 160067 301550
rect 216857 301547 216923 301550
rect 115933 301474 115999 301477
rect 234478 301474 234538 301683
rect 243077 301610 243143 301613
rect 291193 301610 291259 301613
rect 243077 301608 291259 301610
rect 243077 301552 243082 301608
rect 243138 301552 291198 301608
rect 291254 301552 291259 301608
rect 243077 301550 291259 301552
rect 243077 301547 243143 301550
rect 291193 301547 291259 301550
rect 236729 301474 236795 301477
rect 269614 301474 269620 301476
rect 115933 301472 236795 301474
rect 115933 301416 115938 301472
rect 115994 301416 236734 301472
rect 236790 301416 236795 301472
rect 115933 301414 236795 301416
rect 115933 301411 115999 301414
rect 236729 301411 236795 301414
rect 253430 301414 269620 301474
rect 187693 301202 187759 301205
rect 218145 301202 218211 301205
rect 251725 301202 251791 301205
rect 187693 301200 218211 301202
rect 187693 301144 187698 301200
rect 187754 301144 218150 301200
rect 218206 301144 218211 301200
rect 187693 301142 218211 301144
rect 187693 301139 187759 301142
rect 218145 301139 218211 301142
rect 238710 301200 251791 301202
rect 238710 301144 251730 301200
rect 251786 301144 251791 301200
rect 253430 301172 253490 301414
rect 269614 301412 269620 301414
rect 269684 301412 269690 301476
rect 238710 301142 251791 301144
rect 189809 301066 189875 301069
rect 189809 301064 193690 301066
rect 189809 301008 189814 301064
rect 189870 301008 193690 301064
rect 189809 301006 193690 301008
rect 189809 301003 189875 301006
rect 193630 300900 193690 301006
rect 199009 300930 199075 300933
rect 198782 300928 199075 300930
rect 198782 300872 199014 300928
rect 199070 300872 199075 300928
rect 198782 300870 199075 300872
rect 198782 300794 198842 300870
rect 199009 300867 199075 300870
rect 217869 300930 217935 300933
rect 238710 300930 238770 301142
rect 251725 301139 251791 301142
rect 250989 301066 251055 301069
rect 266629 301066 266695 301069
rect 250989 301064 266695 301066
rect 250989 301008 250994 301064
rect 251050 301008 266634 301064
rect 266690 301008 266695 301064
rect 250989 301006 266695 301008
rect 250989 301003 251055 301006
rect 266629 301003 266695 301006
rect 217869 300928 238770 300930
rect 217869 300872 217874 300928
rect 217930 300872 238770 300928
rect 217869 300870 238770 300872
rect 251633 300930 251699 300933
rect 251766 300930 251772 300932
rect 251633 300928 251772 300930
rect 251633 300872 251638 300928
rect 251694 300872 251772 300928
rect 251633 300870 251772 300872
rect 217869 300867 217935 300870
rect 251633 300867 251699 300870
rect 251766 300868 251772 300870
rect 251836 300868 251842 300932
rect 258758 300794 258764 300796
rect 180750 300734 198842 300794
rect 253460 300734 258764 300794
rect 82629 300250 82695 300253
rect 91502 300250 91508 300252
rect 82629 300248 91508 300250
rect 82629 300192 82634 300248
rect 82690 300192 91508 300248
rect 82629 300190 91508 300192
rect 82629 300187 82695 300190
rect 91502 300188 91508 300190
rect 91572 300188 91578 300252
rect 12433 300114 12499 300117
rect 156638 300114 156644 300116
rect 12433 300112 156644 300114
rect 12433 300056 12438 300112
rect 12494 300056 156644 300112
rect 12433 300054 156644 300056
rect 12433 300051 12499 300054
rect 156638 300052 156644 300054
rect 156708 300052 156714 300116
rect 180057 300114 180123 300117
rect 180750 300114 180810 300734
rect 258758 300732 258764 300734
rect 258828 300732 258834 300796
rect 245694 300596 245700 300660
rect 245764 300658 245770 300660
rect 253933 300658 253999 300661
rect 245764 300656 253999 300658
rect 245764 300600 253938 300656
rect 253994 300600 253999 300656
rect 245764 300598 253999 300600
rect 245764 300596 245770 300598
rect 253933 300595 253999 300598
rect 255313 300386 255379 300389
rect 253460 300384 255379 300386
rect 253460 300328 255318 300384
rect 255374 300328 255379 300384
rect 253460 300326 255379 300328
rect 255313 300323 255379 300326
rect 180057 300112 180810 300114
rect 180057 300056 180062 300112
rect 180118 300056 180810 300112
rect 180057 300054 180810 300056
rect 180057 300051 180123 300054
rect 258533 299978 258599 299981
rect 253460 299976 258599 299978
rect 253460 299920 258538 299976
rect 258594 299920 258599 299976
rect 253460 299918 258599 299920
rect 258533 299915 258599 299918
rect 188286 299780 188292 299844
rect 188356 299842 188362 299844
rect 190913 299842 190979 299845
rect 188356 299840 190979 299842
rect 188356 299784 190918 299840
rect 190974 299784 190979 299840
rect 188356 299782 190979 299784
rect 188356 299780 188362 299782
rect 190913 299779 190979 299782
rect 191097 299842 191163 299845
rect 254209 299842 254275 299845
rect 270585 299842 270651 299845
rect 191097 299840 193660 299842
rect 191097 299784 191102 299840
rect 191158 299784 193660 299840
rect 191097 299782 193660 299784
rect 253890 299840 270651 299842
rect 253890 299784 254214 299840
rect 254270 299784 270590 299840
rect 270646 299784 270651 299840
rect 253890 299782 270651 299784
rect 191097 299779 191163 299782
rect 253890 299570 253950 299782
rect 254209 299779 254275 299782
rect 270585 299779 270651 299782
rect 253460 299510 253950 299570
rect 150525 299434 150591 299437
rect 193673 299434 193739 299437
rect 150525 299432 193739 299434
rect 150525 299376 150530 299432
rect 150586 299376 193678 299432
rect 193734 299376 193739 299432
rect 150525 299374 193739 299376
rect 150525 299371 150591 299374
rect 193673 299371 193739 299374
rect 253062 298893 253122 299132
rect 253013 298888 253122 298893
rect 253013 298832 253018 298888
rect 253074 298832 253122 298888
rect 253013 298830 253122 298832
rect 253013 298827 253079 298830
rect 11145 298754 11211 298757
rect 150525 298754 150591 298757
rect 11145 298752 150591 298754
rect 11145 298696 11150 298752
rect 11206 298696 150530 298752
rect 150586 298696 150591 298752
rect 11145 298694 150591 298696
rect 11145 298691 11211 298694
rect 150525 298691 150591 298694
rect 191741 298754 191807 298757
rect 256734 298754 256740 298756
rect 191741 298752 193660 298754
rect 191741 298696 191746 298752
rect 191802 298696 193660 298752
rect 191741 298694 193660 298696
rect 253890 298694 256740 298754
rect 191741 298691 191807 298694
rect 253890 298618 253950 298694
rect 256734 298692 256740 298694
rect 256804 298754 256810 298756
rect 284937 298754 285003 298757
rect 299473 298754 299539 298757
rect 256804 298752 299539 298754
rect 256804 298696 284942 298752
rect 284998 298696 299478 298752
rect 299534 298696 299539 298752
rect 256804 298694 299539 298696
rect 256804 298692 256810 298694
rect 284937 298691 285003 298694
rect 299473 298691 299539 298694
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 253460 298558 253950 298618
rect 583520 298604 584960 298694
rect 256601 298210 256667 298213
rect 253460 298208 256667 298210
rect 253460 298152 256606 298208
rect 256662 298152 256667 298208
rect 253460 298150 256667 298152
rect 256601 298147 256667 298150
rect 252829 298074 252895 298077
rect 252829 298072 253490 298074
rect 252829 298016 252834 298072
rect 252890 298016 253490 298072
rect 252829 298014 253490 298016
rect 252829 298011 252895 298014
rect 253430 297802 253490 298014
rect 258758 298012 258764 298076
rect 258828 298074 258834 298076
rect 273437 298074 273503 298077
rect 258828 298072 273503 298074
rect 258828 298016 273442 298072
rect 273498 298016 273503 298072
rect 258828 298014 273503 298016
rect 258828 298012 258834 298014
rect 273437 298011 273503 298014
rect 255313 297802 255379 297805
rect 253430 297800 255379 297802
rect 253430 297772 255318 297800
rect 253460 297744 255318 297772
rect 255374 297744 255379 297800
rect 253460 297742 255379 297744
rect 255313 297739 255379 297742
rect 191741 297666 191807 297669
rect 252829 297666 252895 297669
rect 253013 297666 253079 297669
rect 191741 297664 193660 297666
rect 191741 297608 191746 297664
rect 191802 297608 193660 297664
rect 191741 297606 193660 297608
rect 252829 297664 253079 297666
rect 252829 297608 252834 297664
rect 252890 297608 253018 297664
rect 253074 297608 253079 297664
rect 252829 297606 253079 297608
rect 191741 297603 191807 297606
rect 252829 297603 252895 297606
rect 253013 297603 253079 297606
rect 168465 297396 168531 297397
rect 154430 297332 154436 297396
rect 154500 297394 154506 297396
rect 168414 297394 168420 297396
rect 154500 297334 168420 297394
rect 168484 297392 168531 297396
rect 255262 297394 255268 297396
rect 168526 297336 168531 297392
rect 154500 297332 154506 297334
rect 168414 297332 168420 297334
rect 168484 297332 168531 297336
rect 253460 297334 255268 297394
rect 255262 297332 255268 297334
rect 255332 297332 255338 297396
rect 168465 297331 168531 297332
rect 253430 296850 253490 296956
rect 269798 296850 269804 296852
rect 253430 296790 269804 296850
rect 269798 296788 269804 296790
rect 269868 296788 269874 296852
rect 273437 296850 273503 296853
rect 278865 296850 278931 296853
rect 273437 296848 278931 296850
rect 273437 296792 273442 296848
rect 273498 296792 278870 296848
rect 278926 296792 278931 296848
rect 273437 296790 278931 296792
rect 273437 296787 273503 296790
rect 278865 296787 278931 296790
rect 253933 296578 253999 296581
rect 253460 296576 253999 296578
rect 126421 296170 126487 296173
rect 145557 296170 145623 296173
rect 126421 296168 145623 296170
rect 126421 296112 126426 296168
rect 126482 296112 145562 296168
rect 145618 296112 145623 296168
rect 126421 296110 145623 296112
rect 126421 296107 126487 296110
rect 145557 296107 145623 296110
rect 36537 296034 36603 296037
rect 180057 296034 180123 296037
rect 36537 296032 180123 296034
rect 36537 295976 36542 296032
rect 36598 295976 180062 296032
rect 180118 295976 180123 296032
rect 36537 295974 180123 295976
rect 36537 295971 36603 295974
rect 180057 295971 180123 295974
rect 192017 296034 192083 296037
rect 193630 296034 193690 296548
rect 253460 296520 253938 296576
rect 253994 296520 253999 296576
rect 253460 296518 253999 296520
rect 253933 296515 253999 296518
rect 255589 296170 255655 296173
rect 256601 296170 256667 296173
rect 253460 296168 256667 296170
rect 253460 296112 255594 296168
rect 255650 296112 256606 296168
rect 256662 296112 256667 296168
rect 253460 296110 256667 296112
rect 255589 296107 255655 296110
rect 256601 296107 256667 296110
rect 192017 296032 193690 296034
rect 192017 295976 192022 296032
rect 192078 295976 193690 296032
rect 192017 295974 193690 295976
rect 192017 295971 192083 295974
rect 254025 295626 254091 295629
rect 253460 295624 254091 295626
rect 253460 295568 254030 295624
rect 254086 295568 254091 295624
rect 253460 295566 254091 295568
rect 254025 295563 254091 295566
rect 190177 295490 190243 295493
rect 190177 295488 193660 295490
rect 190177 295432 190182 295488
rect 190238 295432 193660 295488
rect 190177 295430 193660 295432
rect 190177 295427 190243 295430
rect 145557 295354 145623 295357
rect 192017 295354 192083 295357
rect 145557 295352 192083 295354
rect 145557 295296 145562 295352
rect 145618 295296 192022 295352
rect 192078 295296 192083 295352
rect 145557 295294 192083 295296
rect 145557 295291 145623 295294
rect 192017 295291 192083 295294
rect 260833 295218 260899 295221
rect 268009 295218 268075 295221
rect 253460 295216 268075 295218
rect 253460 295160 260838 295216
rect 260894 295160 268014 295216
rect 268070 295160 268075 295216
rect 253460 295158 268075 295160
rect 260833 295155 260899 295158
rect 268009 295155 268075 295158
rect 256325 294810 256391 294813
rect 253460 294808 256391 294810
rect 253460 294752 256330 294808
rect 256386 294752 256391 294808
rect 253460 294750 256391 294752
rect 256325 294747 256391 294750
rect 4153 294538 4219 294541
rect 138657 294538 138723 294541
rect 4153 294536 138723 294538
rect 4153 294480 4158 294536
rect 4214 294480 138662 294536
rect 138718 294480 138723 294536
rect 4153 294478 138723 294480
rect 4153 294475 4219 294478
rect 138657 294475 138723 294478
rect 191741 294402 191807 294405
rect 256601 294402 256667 294405
rect 191741 294400 193660 294402
rect 191741 294344 191746 294400
rect 191802 294344 193660 294400
rect 191741 294342 193660 294344
rect 253460 294400 256667 294402
rect 253460 294344 256606 294400
rect 256662 294344 256667 294400
rect 253460 294342 256667 294344
rect 191741 294339 191807 294342
rect 256601 294339 256667 294342
rect 258390 293994 258396 293996
rect 253460 293934 258396 293994
rect 258390 293932 258396 293934
rect 258460 293932 258466 293996
rect 258809 293858 258875 293861
rect 275001 293858 275067 293861
rect 258809 293856 275067 293858
rect 258809 293800 258814 293856
rect 258870 293800 275006 293856
rect 275062 293800 275067 293856
rect 258809 293798 275067 293800
rect 258809 293795 258875 293798
rect 275001 293795 275067 293798
rect 259678 293586 259684 293588
rect 252908 293556 259684 293586
rect 252878 293526 259684 293556
rect 252878 293453 252938 293526
rect 259678 293524 259684 293526
rect 259748 293524 259754 293588
rect 252829 293448 252938 293453
rect 252829 293392 252834 293448
rect 252890 293392 252938 293448
rect 252829 293390 252938 293392
rect 252829 293387 252895 293390
rect 191557 293314 191623 293317
rect 191557 293312 193660 293314
rect -960 293178 480 293268
rect 191557 293256 191562 293312
rect 191618 293256 193660 293312
rect 191557 293254 193660 293256
rect 191557 293251 191623 293254
rect 3509 293178 3575 293181
rect 254117 293178 254183 293181
rect 256141 293178 256207 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect 253460 293176 256207 293178
rect 253460 293120 254122 293176
rect 254178 293120 256146 293176
rect 256202 293120 256207 293176
rect 253460 293118 256207 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 254117 293115 254183 293118
rect 256141 293115 256207 293118
rect 75453 292634 75519 292637
rect 81934 292634 81940 292636
rect 75453 292632 81940 292634
rect 75453 292576 75458 292632
rect 75514 292576 81940 292632
rect 75453 292574 81940 292576
rect 75453 292571 75519 292574
rect 81934 292572 81940 292574
rect 82004 292572 82010 292636
rect 255957 292634 256023 292637
rect 253460 292632 256023 292634
rect 253460 292576 255962 292632
rect 256018 292576 256023 292632
rect 253460 292574 256023 292576
rect 255957 292571 256023 292574
rect 275001 292634 275067 292637
rect 276197 292634 276263 292637
rect 275001 292632 276263 292634
rect 275001 292576 275006 292632
rect 275062 292576 276202 292632
rect 276258 292576 276263 292632
rect 275001 292574 276263 292576
rect 275001 292571 275067 292574
rect 276197 292571 276263 292574
rect 193029 292226 193095 292229
rect 259637 292226 259703 292229
rect 193029 292224 193660 292226
rect 193029 292168 193034 292224
rect 193090 292168 193660 292224
rect 193029 292166 193660 292168
rect 253460 292224 259703 292226
rect 253460 292168 259642 292224
rect 259698 292168 259703 292224
rect 253460 292166 259703 292168
rect 193029 292163 193095 292166
rect 259637 292163 259703 292166
rect 125041 291818 125107 291821
rect 160686 291818 160692 291820
rect 125041 291816 160692 291818
rect 125041 291760 125046 291816
rect 125102 291760 160692 291816
rect 125041 291758 160692 291760
rect 125041 291755 125107 291758
rect 160686 291756 160692 291758
rect 160756 291756 160762 291820
rect 166206 291756 166212 291820
rect 166276 291818 166282 291820
rect 185342 291818 185348 291820
rect 166276 291758 185348 291818
rect 166276 291756 166282 291758
rect 185342 291756 185348 291758
rect 185412 291756 185418 291820
rect 255957 291818 256023 291821
rect 253460 291816 256023 291818
rect 253460 291760 255962 291816
rect 256018 291760 256023 291816
rect 253460 291758 256023 291760
rect 255957 291755 256023 291758
rect 260741 291818 260807 291821
rect 285673 291818 285739 291821
rect 260741 291816 285739 291818
rect 260741 291760 260746 291816
rect 260802 291760 285678 291816
rect 285734 291760 285739 291816
rect 260741 291758 285739 291760
rect 260741 291755 260807 291758
rect 285673 291755 285739 291758
rect 255681 291682 255747 291685
rect 262213 291682 262279 291685
rect 253430 291680 262279 291682
rect 253430 291624 255686 291680
rect 255742 291624 262218 291680
rect 262274 291624 262279 291680
rect 253430 291622 262279 291624
rect 190361 291410 190427 291413
rect 193029 291410 193095 291413
rect 190361 291408 193095 291410
rect 190361 291352 190366 291408
rect 190422 291352 193034 291408
rect 193090 291352 193095 291408
rect 253430 291380 253490 291622
rect 255681 291619 255747 291622
rect 262213 291619 262279 291622
rect 190361 291350 193095 291352
rect 190361 291347 190427 291350
rect 193029 291347 193095 291350
rect 191649 291138 191715 291141
rect 256601 291138 256667 291141
rect 191649 291136 193660 291138
rect 191649 291080 191654 291136
rect 191710 291080 193660 291136
rect 191649 291078 193660 291080
rect 253430 291136 256667 291138
rect 253430 291080 256606 291136
rect 256662 291080 256667 291136
rect 253430 291078 256667 291080
rect 191649 291075 191715 291078
rect 253430 290972 253490 291078
rect 256601 291075 256667 291078
rect 258165 290866 258231 290869
rect 258390 290866 258396 290868
rect 258165 290864 258396 290866
rect 258165 290808 258170 290864
rect 258226 290808 258396 290864
rect 258165 290806 258396 290808
rect 258165 290803 258231 290806
rect 258390 290804 258396 290806
rect 258460 290804 258466 290868
rect 253430 290322 253490 290564
rect 253430 290262 258090 290322
rect 191189 290050 191255 290053
rect 255497 290050 255563 290053
rect 191189 290048 193660 290050
rect 191189 289992 191194 290048
rect 191250 289992 193660 290048
rect 191189 289990 193660 289992
rect 253460 290048 255563 290050
rect 253460 289992 255502 290048
rect 255558 289992 255563 290048
rect 253460 289990 255563 289992
rect 191189 289987 191255 289990
rect 255497 289987 255563 289990
rect 80881 289914 80947 289917
rect 81014 289914 81020 289916
rect 80881 289912 81020 289914
rect 80881 289856 80886 289912
rect 80942 289856 81020 289912
rect 80881 289854 81020 289856
rect 80881 289851 80947 289854
rect 81014 289852 81020 289854
rect 81084 289914 81090 289916
rect 100017 289914 100083 289917
rect 81084 289912 100083 289914
rect 81084 289856 100022 289912
rect 100078 289856 100083 289912
rect 81084 289854 100083 289856
rect 258030 289914 258090 290262
rect 582557 289914 582623 289917
rect 258030 289912 582623 289914
rect 258030 289856 582562 289912
rect 582618 289856 582623 289912
rect 258030 289854 582623 289856
rect 81084 289852 81090 289854
rect 100017 289851 100083 289854
rect 582557 289851 582623 289854
rect 175273 289778 175339 289781
rect 176101 289778 176167 289781
rect 259678 289778 259684 289780
rect 175273 289776 176167 289778
rect 175273 289720 175278 289776
rect 175334 289720 176106 289776
rect 176162 289720 176167 289776
rect 175273 289718 176167 289720
rect 175273 289715 175339 289718
rect 176101 289715 176167 289718
rect 253430 289718 259684 289778
rect 253430 289612 253490 289718
rect 259678 289716 259684 289718
rect 259748 289778 259754 289780
rect 260741 289778 260807 289781
rect 259748 289776 260807 289778
rect 259748 289720 260746 289776
rect 260802 289720 260807 289776
rect 259748 289718 260807 289720
rect 259748 289716 259754 289718
rect 260741 289715 260807 289718
rect 255497 289234 255563 289237
rect 253460 289232 255563 289234
rect 253460 289176 255502 289232
rect 255558 289176 255563 289232
rect 253460 289174 255563 289176
rect 255497 289171 255563 289174
rect 50889 289098 50955 289101
rect 175273 289098 175339 289101
rect 50889 289096 175339 289098
rect 50889 289040 50894 289096
rect 50950 289040 175278 289096
rect 175334 289040 175339 289096
rect 50889 289038 175339 289040
rect 50889 289035 50955 289038
rect 175273 289035 175339 289038
rect 191741 288962 191807 288965
rect 191741 288960 193660 288962
rect 191741 288904 191746 288960
rect 191802 288904 193660 288960
rect 191741 288902 193660 288904
rect 191741 288899 191807 288902
rect 259494 288826 259500 288828
rect 253460 288766 259500 288826
rect 259494 288764 259500 288766
rect 259564 288764 259570 288828
rect 91502 288492 91508 288556
rect 91572 288554 91578 288556
rect 95233 288554 95299 288557
rect 91572 288552 95299 288554
rect 91572 288496 95238 288552
rect 95294 288496 95299 288552
rect 91572 288494 95299 288496
rect 91572 288492 91578 288494
rect 95233 288491 95299 288494
rect 268101 288418 268167 288421
rect 269205 288418 269271 288421
rect 253460 288416 269271 288418
rect 253460 288360 268106 288416
rect 268162 288360 269210 288416
rect 269266 288360 269271 288416
rect 253460 288358 269271 288360
rect 268101 288355 268167 288358
rect 269205 288355 269271 288358
rect 255497 288010 255563 288013
rect 253460 288008 255563 288010
rect 253460 287952 255502 288008
rect 255558 287952 255563 288008
rect 253460 287950 255563 287952
rect 255497 287947 255563 287950
rect 88977 287738 89043 287741
rect 99966 287738 99972 287740
rect 88977 287736 99972 287738
rect 88977 287680 88982 287736
rect 89038 287680 99972 287736
rect 88977 287678 99972 287680
rect 88977 287675 89043 287678
rect 99966 287676 99972 287678
rect 100036 287676 100042 287740
rect 107561 287738 107627 287741
rect 166809 287738 166875 287741
rect 179321 287738 179387 287741
rect 107561 287736 180810 287738
rect 107561 287680 107566 287736
rect 107622 287680 166814 287736
rect 166870 287680 179326 287736
rect 179382 287680 180810 287736
rect 107561 287678 180810 287680
rect 107561 287675 107627 287678
rect 166809 287675 166875 287678
rect 179321 287675 179387 287678
rect 85849 287194 85915 287197
rect 86769 287194 86835 287197
rect 102133 287194 102199 287197
rect 85849 287192 102199 287194
rect 85849 287136 85854 287192
rect 85910 287136 86774 287192
rect 86830 287136 102138 287192
rect 102194 287136 102199 287192
rect 85849 287134 102199 287136
rect 180750 287194 180810 287678
rect 193630 287194 193690 287844
rect 255313 287602 255379 287605
rect 253460 287600 255379 287602
rect 253460 287544 255318 287600
rect 255374 287544 255379 287600
rect 253460 287542 255379 287544
rect 255313 287539 255379 287542
rect 180750 287134 193690 287194
rect 85849 287131 85915 287134
rect 86769 287131 86835 287134
rect 102133 287131 102199 287134
rect 79174 286996 79180 287060
rect 79244 287058 79250 287060
rect 79317 287058 79383 287061
rect 257429 287058 257495 287061
rect 79244 287056 79383 287058
rect 79244 287000 79322 287056
rect 79378 287000 79383 287056
rect 79244 286998 79383 287000
rect 253460 287056 257495 287058
rect 253460 287000 257434 287056
rect 257490 287000 257495 287056
rect 253460 286998 257495 287000
rect 79244 286996 79250 286998
rect 79317 286995 79383 286998
rect 257429 286995 257495 286998
rect 191741 286786 191807 286789
rect 191741 286784 193660 286786
rect 191741 286728 191746 286784
rect 191802 286728 193660 286784
rect 191741 286726 193660 286728
rect 191741 286723 191807 286726
rect 255405 286650 255471 286653
rect 253460 286648 255471 286650
rect 253460 286592 255410 286648
rect 255466 286592 255471 286648
rect 253460 286590 255471 286592
rect 255405 286587 255471 286590
rect 257429 286514 257495 286517
rect 267733 286514 267799 286517
rect 257429 286512 267799 286514
rect 257429 286456 257434 286512
rect 257490 286456 267738 286512
rect 267794 286456 267799 286512
rect 257429 286454 267799 286456
rect 257429 286451 257495 286454
rect 267733 286451 267799 286454
rect 281625 286378 281691 286381
rect 258030 286376 281691 286378
rect 258030 286320 281630 286376
rect 281686 286320 281691 286376
rect 258030 286318 281691 286320
rect 255497 286242 255563 286245
rect 253460 286240 255563 286242
rect 253460 286184 255502 286240
rect 255558 286184 255563 286240
rect 253460 286182 255563 286184
rect 255497 286179 255563 286182
rect 90265 286106 90331 286109
rect 91001 286106 91067 286109
rect 256693 286106 256759 286109
rect 258030 286106 258090 286318
rect 281625 286315 281691 286318
rect 90265 286104 91067 286106
rect 90265 286048 90270 286104
rect 90326 286048 91006 286104
rect 91062 286048 91067 286104
rect 90265 286046 91067 286048
rect 90265 286043 90331 286046
rect 91001 286043 91067 286046
rect 253430 286104 258090 286106
rect 253430 286048 256698 286104
rect 256754 286048 258090 286104
rect 253430 286046 258090 286048
rect 68461 285970 68527 285973
rect 79317 285970 79383 285973
rect 68461 285968 79383 285970
rect 68461 285912 68466 285968
rect 68522 285912 79322 285968
rect 79378 285912 79383 285968
rect 68461 285910 79383 285912
rect 68461 285907 68527 285910
rect 79317 285907 79383 285910
rect 83089 285970 83155 285973
rect 84101 285970 84167 285973
rect 83089 285968 89730 285970
rect 83089 285912 83094 285968
rect 83150 285912 84106 285968
rect 84162 285912 89730 285968
rect 83089 285910 89730 285912
rect 83089 285907 83155 285910
rect 84101 285907 84167 285910
rect 73286 285772 73292 285836
rect 73356 285834 73362 285836
rect 80421 285834 80487 285837
rect 73356 285832 80487 285834
rect 73356 285776 80426 285832
rect 80482 285776 80487 285832
rect 73356 285774 80487 285776
rect 73356 285772 73362 285774
rect 80421 285771 80487 285774
rect 82629 285834 82695 285837
rect 87086 285834 87092 285836
rect 82629 285832 87092 285834
rect 82629 285776 82634 285832
rect 82690 285776 87092 285832
rect 82629 285774 87092 285776
rect 82629 285771 82695 285774
rect 87086 285772 87092 285774
rect 87156 285772 87162 285836
rect 89670 285834 89730 285910
rect 104433 285834 104499 285837
rect 89670 285832 104499 285834
rect 89670 285776 104438 285832
rect 104494 285776 104499 285832
rect 253430 285804 253490 286046
rect 256693 286043 256759 286046
rect 89670 285774 104499 285776
rect 104433 285771 104499 285774
rect 93945 285698 94011 285701
rect 152641 285698 152707 285701
rect 93945 285696 152707 285698
rect 93945 285640 93950 285696
rect 94006 285640 152646 285696
rect 152702 285640 152707 285696
rect 93945 285638 152707 285640
rect 93945 285635 94011 285638
rect 152641 285635 152707 285638
rect 189717 285698 189783 285701
rect 189717 285696 193660 285698
rect 189717 285640 189722 285696
rect 189778 285640 193660 285696
rect 189717 285638 193660 285640
rect 189717 285635 189783 285638
rect 74625 285562 74691 285565
rect 75453 285562 75519 285565
rect 74625 285560 75519 285562
rect 74625 285504 74630 285560
rect 74686 285504 75458 285560
rect 75514 285504 75519 285560
rect 74625 285502 75519 285504
rect 74625 285499 74691 285502
rect 75453 285499 75519 285502
rect 84653 285564 84719 285565
rect 84653 285560 84700 285564
rect 84764 285562 84770 285564
rect 84653 285504 84658 285560
rect 84653 285500 84700 285504
rect 84764 285502 84810 285562
rect 84764 285500 84770 285502
rect 91134 285500 91140 285564
rect 91204 285562 91210 285564
rect 91277 285562 91343 285565
rect 91204 285560 91343 285562
rect 91204 285504 91282 285560
rect 91338 285504 91343 285560
rect 91204 285502 91343 285504
rect 91204 285500 91210 285502
rect 84653 285499 84719 285500
rect 91277 285499 91343 285502
rect 255405 285426 255471 285429
rect 253460 285424 255471 285426
rect 253460 285368 255410 285424
rect 255466 285368 255471 285424
rect 253460 285366 255471 285368
rect 255405 285363 255471 285366
rect 583520 285276 584960 285516
rect 262397 285018 262463 285021
rect 253460 285016 262463 285018
rect 253460 284960 262402 285016
rect 262458 284960 262463 285016
rect 253460 284958 262463 284960
rect 262397 284955 262463 284958
rect 97901 284882 97967 284885
rect 162117 284882 162183 284885
rect 266537 284882 266603 284885
rect 97901 284880 162183 284882
rect 97901 284824 97906 284880
rect 97962 284824 162122 284880
rect 162178 284824 162183 284880
rect 97901 284822 162183 284824
rect 97901 284819 97967 284822
rect 162117 284819 162183 284822
rect 253430 284880 266603 284882
rect 253430 284824 266542 284880
rect 266598 284824 266603 284880
rect 253430 284822 266603 284824
rect 59169 284610 59235 284613
rect 99097 284610 99163 284613
rect 59169 284608 99163 284610
rect 59169 284552 59174 284608
rect 59230 284552 99102 284608
rect 99158 284552 99163 284608
rect 59169 284550 99163 284552
rect 59169 284547 59235 284550
rect 99097 284547 99163 284550
rect 191741 284610 191807 284613
rect 191741 284608 193660 284610
rect 191741 284552 191746 284608
rect 191802 284552 193660 284608
rect 253430 284580 253490 284822
rect 266537 284819 266603 284822
rect 191741 284550 193660 284552
rect 191741 284547 191807 284550
rect 75269 284474 75335 284477
rect 70166 284472 75335 284474
rect 70166 284416 75274 284472
rect 75330 284416 75335 284472
rect 70166 284414 75335 284416
rect 70166 284204 70226 284414
rect 75269 284411 75335 284414
rect 78213 284474 78279 284477
rect 98085 284474 98151 284477
rect 78213 284472 98151 284474
rect 78213 284416 78218 284472
rect 78274 284416 98090 284472
rect 98146 284416 98151 284472
rect 78213 284414 98151 284416
rect 78213 284411 78279 284414
rect 98085 284411 98151 284414
rect 72918 284276 72924 284340
rect 72988 284338 72994 284340
rect 74625 284338 74691 284341
rect 72988 284336 74691 284338
rect 72988 284280 74630 284336
rect 74686 284280 74691 284336
rect 72988 284278 74691 284280
rect 72988 284276 72994 284278
rect 74625 284275 74691 284278
rect 262397 284338 262463 284341
rect 263961 284338 264027 284341
rect 262397 284336 264027 284338
rect 262397 284280 262402 284336
rect 262458 284280 263966 284336
rect 264022 284280 264027 284336
rect 262397 284278 264027 284280
rect 262397 284275 262463 284278
rect 263961 284275 264027 284278
rect 67398 284140 67404 284204
rect 67468 284202 67474 284204
rect 69238 284202 69244 284204
rect 67468 284142 69244 284202
rect 67468 284140 67474 284142
rect 69238 284140 69244 284142
rect 69308 284140 69314 284204
rect 70158 284140 70164 284204
rect 70228 284140 70234 284204
rect 255405 284066 255471 284069
rect 253460 284064 255471 284066
rect 253460 284008 255410 284064
rect 255466 284008 255471 284064
rect 253460 284006 255471 284008
rect 255405 284003 255471 284006
rect 69197 283794 69263 283797
rect 70071 283794 70137 283797
rect 69197 283792 70137 283794
rect 69197 283736 69202 283792
rect 69258 283736 70076 283792
rect 70132 283736 70137 283792
rect 69197 283734 70137 283736
rect 69197 283731 69263 283734
rect 70071 283731 70137 283734
rect 71630 283732 71636 283796
rect 71700 283794 71706 283796
rect 71957 283794 72023 283797
rect 72831 283794 72897 283797
rect 71700 283792 72897 283794
rect 71700 283736 71962 283792
rect 72018 283736 72836 283792
rect 72892 283736 72897 283792
rect 71700 283734 72897 283736
rect 71700 283732 71706 283734
rect 71957 283731 72023 283734
rect 72831 283731 72897 283734
rect 86718 283596 86724 283660
rect 86788 283658 86794 283660
rect 86861 283658 86927 283661
rect 86788 283656 86927 283658
rect 86788 283600 86866 283656
rect 86922 283600 86927 283656
rect 86788 283598 86927 283600
rect 86788 283596 86794 283598
rect 86861 283595 86927 283598
rect 70209 283522 70275 283525
rect 89805 283524 89871 283525
rect 70209 283520 80070 283522
rect 70209 283464 70214 283520
rect 70270 283464 80070 283520
rect 70209 283462 80070 283464
rect 70209 283459 70275 283462
rect 80010 283386 80070 283462
rect 89805 283520 89852 283524
rect 89916 283522 89922 283524
rect 89805 283464 89810 283520
rect 89805 283460 89852 283464
rect 89916 283462 89962 283522
rect 89916 283460 89922 283462
rect 93710 283460 93716 283524
rect 93780 283522 93786 283524
rect 94037 283522 94103 283525
rect 93780 283520 94103 283522
rect 93780 283464 94042 283520
rect 94098 283464 94103 283520
rect 93780 283462 94103 283464
rect 93780 283460 93786 283462
rect 89805 283459 89871 283460
rect 94037 283459 94103 283462
rect 94262 283460 94268 283524
rect 94332 283522 94338 283524
rect 94681 283522 94747 283525
rect 94332 283520 94747 283522
rect 94332 283464 94686 283520
rect 94742 283464 94747 283520
rect 94332 283462 94747 283464
rect 94332 283460 94338 283462
rect 94681 283459 94747 283462
rect 191741 283522 191807 283525
rect 253430 283522 253490 283628
rect 264973 283522 265039 283525
rect 191741 283520 193660 283522
rect 191741 283464 191746 283520
rect 191802 283464 193660 283520
rect 191741 283462 193660 283464
rect 253430 283520 265039 283522
rect 253430 283464 264978 283520
rect 265034 283464 265039 283520
rect 253430 283462 265039 283464
rect 191741 283459 191807 283462
rect 264973 283459 265039 283462
rect 269798 283460 269804 283524
rect 269868 283522 269874 283524
rect 281533 283522 281599 283525
rect 269868 283520 281599 283522
rect 269868 283464 281538 283520
rect 281594 283464 281599 283520
rect 269868 283462 281599 283464
rect 269868 283460 269874 283462
rect 281533 283459 281599 283462
rect 98913 283386 98979 283389
rect 65934 283326 75194 283386
rect 80010 283384 98979 283386
rect 80010 283328 98918 283384
rect 98974 283328 98979 283384
rect 80010 283326 98979 283328
rect 65934 283253 65994 283326
rect 59261 283250 59327 283253
rect 65885 283250 65994 283253
rect 59261 283248 65994 283250
rect 59261 283192 59266 283248
rect 59322 283192 65890 283248
rect 65946 283192 65994 283248
rect 59261 283190 65994 283192
rect 59261 283187 59327 283190
rect 65885 283187 65951 283190
rect 68686 283188 68692 283252
rect 68756 283250 68762 283252
rect 70945 283250 71011 283253
rect 68756 283248 71011 283250
rect 68756 283192 70950 283248
rect 71006 283192 71011 283248
rect 68756 283190 71011 283192
rect 68756 283188 68762 283190
rect 70945 283187 71011 283190
rect 71814 283188 71820 283252
rect 71884 283250 71890 283252
rect 71957 283250 72023 283253
rect 71884 283248 72023 283250
rect 71884 283192 71962 283248
rect 72018 283192 72023 283248
rect 71884 283190 72023 283192
rect 71884 283188 71890 283190
rect 71957 283187 72023 283190
rect 73102 283188 73108 283252
rect 73172 283250 73178 283252
rect 73245 283250 73311 283253
rect 73172 283248 73311 283250
rect 73172 283192 73250 283248
rect 73306 283192 73311 283248
rect 73172 283190 73311 283192
rect 75134 283250 75194 283326
rect 98913 283323 98979 283326
rect 98862 283250 98868 283252
rect 75134 283190 98868 283250
rect 73172 283188 73178 283190
rect 73245 283187 73311 283190
rect 98862 283188 98868 283190
rect 98932 283188 98938 283252
rect 255497 283250 255563 283253
rect 253460 283248 255563 283250
rect 253460 283192 255502 283248
rect 255558 283192 255563 283248
rect 253460 283190 255563 283192
rect 255497 283187 255563 283190
rect 83457 283116 83523 283117
rect 83406 283114 83412 283116
rect 83366 283054 83412 283114
rect 83476 283112 83523 283116
rect 83518 283056 83523 283112
rect 83406 283052 83412 283054
rect 83476 283052 83523 283056
rect 83457 283051 83523 283052
rect 88609 283114 88675 283117
rect 88742 283114 88748 283116
rect 88609 283112 88748 283114
rect 88609 283056 88614 283112
rect 88670 283056 88748 283112
rect 88609 283054 88748 283056
rect 88609 283051 88675 283054
rect 88742 283052 88748 283054
rect 88812 283052 88818 283116
rect 92381 283114 92447 283117
rect 100201 283114 100267 283117
rect 92381 283112 100267 283114
rect 92381 283056 92386 283112
rect 92442 283056 100206 283112
rect 100262 283056 100267 283112
rect 92381 283054 100267 283056
rect 92381 283051 92447 283054
rect 100201 283051 100267 283054
rect 66253 282978 66319 282981
rect 95325 282980 95391 282981
rect 66253 282976 68908 282978
rect 66253 282920 66258 282976
rect 66314 282920 68908 282976
rect 66253 282918 68908 282920
rect 95325 282976 95372 282980
rect 95436 282978 95442 282980
rect 95325 282920 95330 282976
rect 66253 282915 66319 282918
rect 95325 282916 95372 282920
rect 95436 282918 95482 282978
rect 95436 282916 95442 282918
rect 159766 282916 159772 282980
rect 159836 282978 159842 282980
rect 160277 282978 160343 282981
rect 159836 282976 160343 282978
rect 159836 282920 160282 282976
rect 160338 282920 160343 282976
rect 159836 282918 160343 282920
rect 159836 282916 159842 282918
rect 95325 282915 95391 282916
rect 160277 282915 160343 282918
rect 98913 282842 98979 282845
rect 143441 282842 143507 282845
rect 98913 282840 143507 282842
rect 98913 282784 98918 282840
rect 98974 282784 143446 282840
rect 143502 282784 143507 282840
rect 98913 282782 143507 282784
rect 98913 282779 98979 282782
rect 143441 282779 143507 282782
rect 69013 282706 69079 282709
rect 101489 282706 101555 282709
rect 69013 282704 69122 282706
rect 69013 282648 69018 282704
rect 69074 282648 69122 282704
rect 69013 282643 69122 282648
rect 98716 282704 101555 282706
rect 98716 282648 101494 282704
rect 101550 282648 101555 282704
rect 98716 282646 101555 282648
rect 253430 282706 253490 282812
rect 266445 282706 266511 282709
rect 253430 282704 266511 282706
rect 253430 282648 266450 282704
rect 266506 282648 266511 282704
rect 253430 282646 266511 282648
rect 101489 282643 101555 282646
rect 266445 282643 266511 282646
rect 61929 282162 61995 282165
rect 68553 282162 68619 282165
rect 61929 282160 68619 282162
rect 61929 282104 61934 282160
rect 61990 282104 68558 282160
rect 68614 282104 68619 282160
rect 69062 282132 69122 282643
rect 191741 282434 191807 282437
rect 255405 282434 255471 282437
rect 191741 282432 193660 282434
rect 191741 282376 191746 282432
rect 191802 282376 193660 282432
rect 191741 282374 193660 282376
rect 253460 282432 255471 282434
rect 253460 282376 255410 282432
rect 255466 282376 255471 282432
rect 253460 282374 255471 282376
rect 191741 282371 191807 282374
rect 255405 282371 255471 282374
rect 143441 282162 143507 282165
rect 168373 282162 168439 282165
rect 143441 282160 168439 282162
rect 61929 282102 68619 282104
rect 61929 282099 61995 282102
rect 68553 282099 68619 282102
rect 143441 282104 143446 282160
rect 143502 282104 168378 282160
rect 168434 282104 168439 282160
rect 143441 282102 168439 282104
rect 143441 282099 143507 282102
rect 168373 282099 168439 282102
rect 255497 282026 255563 282029
rect 253460 282024 255563 282026
rect 253460 281968 255502 282024
rect 255558 281968 255563 282024
rect 253460 281966 255563 281968
rect 255497 281963 255563 281966
rect 100753 281890 100819 281893
rect 98716 281888 100819 281890
rect 98716 281832 100758 281888
rect 100814 281832 100819 281888
rect 98716 281830 100819 281832
rect 100753 281827 100819 281830
rect 259361 281618 259427 281621
rect 273437 281618 273503 281621
rect 259361 281616 273503 281618
rect 259361 281560 259366 281616
rect 259422 281560 273442 281616
rect 273498 281560 273503 281616
rect 259361 281558 273503 281560
rect 259361 281555 259427 281558
rect 273437 281555 273503 281558
rect 160093 281482 160159 281485
rect 189717 281482 189783 281485
rect 255405 281482 255471 281485
rect 160093 281480 189783 281482
rect 160093 281424 160098 281480
rect 160154 281424 189722 281480
rect 189778 281424 189783 281480
rect 160093 281422 189783 281424
rect 253460 281480 255471 281482
rect 253460 281424 255410 281480
rect 255466 281424 255471 281480
rect 253460 281422 255471 281424
rect 160093 281419 160159 281422
rect 189717 281419 189783 281422
rect 255405 281419 255471 281422
rect 191741 281346 191807 281349
rect 191741 281344 193660 281346
rect 68878 281213 68938 281316
rect 191741 281288 191746 281344
rect 191802 281288 193660 281344
rect 191741 281286 193660 281288
rect 191741 281283 191807 281286
rect 68878 281208 68987 281213
rect 68878 281152 68926 281208
rect 68982 281152 68987 281208
rect 68878 281150 68987 281152
rect 68921 281147 68987 281150
rect 259269 281074 259335 281077
rect 253460 281072 259335 281074
rect 67909 280530 67975 280533
rect 98686 280530 98746 281044
rect 253460 281016 259274 281072
rect 259330 281016 259335 281072
rect 253460 281014 259335 281016
rect 259269 281011 259335 281014
rect 112621 280802 112687 280805
rect 160093 280802 160159 280805
rect 265065 280802 265131 280805
rect 112621 280800 160159 280802
rect 112621 280744 112626 280800
rect 112682 280744 160098 280800
rect 160154 280744 160159 280800
rect 112621 280742 160159 280744
rect 112621 280739 112687 280742
rect 160093 280739 160159 280742
rect 253430 280800 265131 280802
rect 253430 280744 265070 280800
rect 265126 280744 265131 280800
rect 253430 280742 265131 280744
rect 253430 280636 253490 280742
rect 265065 280739 265131 280742
rect 142981 280530 143047 280533
rect 67909 280528 68908 280530
rect 67909 280472 67914 280528
rect 67970 280472 68908 280528
rect 67909 280470 68908 280472
rect 98686 280528 143047 280530
rect 98686 280472 142986 280528
rect 143042 280472 143047 280528
rect 98686 280470 143047 280472
rect 67909 280467 67975 280470
rect 142981 280467 143047 280470
rect 99966 280258 99972 280260
rect -960 279972 480 280212
rect 98716 280198 99972 280258
rect 99966 280196 99972 280198
rect 100036 280258 100042 280260
rect 100845 280258 100911 280261
rect 100036 280256 100911 280258
rect 100036 280200 100850 280256
rect 100906 280200 100911 280256
rect 100036 280198 100911 280200
rect 100036 280196 100042 280198
rect 100845 280195 100911 280198
rect 192017 280258 192083 280261
rect 255497 280258 255563 280261
rect 192017 280256 193660 280258
rect 192017 280200 192022 280256
rect 192078 280200 193660 280256
rect 192017 280198 193660 280200
rect 253460 280256 255563 280258
rect 253460 280200 255502 280256
rect 255558 280200 255563 280256
rect 253460 280198 255563 280200
rect 192017 280195 192083 280198
rect 255497 280195 255563 280198
rect 166809 280122 166875 280125
rect 167085 280122 167151 280125
rect 166809 280120 167151 280122
rect 166809 280064 166814 280120
rect 166870 280064 167090 280120
rect 167146 280064 167151 280120
rect 166809 280062 167151 280064
rect 166809 280059 166875 280062
rect 167085 280059 167151 280062
rect 259821 279850 259887 279853
rect 253460 279848 267750 279850
rect 253460 279792 259826 279848
rect 259882 279792 267750 279848
rect 253460 279790 267750 279792
rect 259821 279787 259887 279790
rect 67541 279714 67607 279717
rect 67541 279712 68908 279714
rect 67541 279656 67546 279712
rect 67602 279656 68908 279712
rect 67541 279654 68908 279656
rect 67541 279651 67607 279654
rect 99097 279578 99163 279581
rect 99097 279576 103530 279578
rect 99097 279520 99102 279576
rect 99158 279520 103530 279576
rect 99097 279518 103530 279520
rect 99097 279515 99163 279518
rect 100753 279442 100819 279445
rect 98716 279440 100819 279442
rect 98716 279384 100758 279440
rect 100814 279384 100819 279440
rect 98716 279382 100819 279384
rect 103470 279442 103530 279518
rect 166809 279442 166875 279445
rect 259453 279442 259519 279445
rect 264973 279442 265039 279445
rect 103470 279440 166875 279442
rect 103470 279384 166814 279440
rect 166870 279384 166875 279440
rect 103470 279382 166875 279384
rect 253460 279440 265039 279442
rect 253460 279384 259458 279440
rect 259514 279384 264978 279440
rect 265034 279384 265039 279440
rect 253460 279382 265039 279384
rect 267690 279442 267750 279790
rect 283189 279442 283255 279445
rect 267690 279440 283255 279442
rect 267690 279384 283194 279440
rect 283250 279384 283255 279440
rect 267690 279382 283255 279384
rect 100753 279379 100819 279382
rect 166809 279379 166875 279382
rect 259453 279379 259519 279382
rect 264973 279379 265039 279382
rect 283189 279379 283255 279382
rect 191741 279170 191807 279173
rect 191741 279168 193660 279170
rect 191741 279112 191746 279168
rect 191802 279112 193660 279168
rect 191741 279110 193660 279112
rect 191741 279107 191807 279110
rect 255497 279034 255563 279037
rect 253460 279032 255563 279034
rect 253460 278976 255502 279032
rect 255558 278976 255563 279032
rect 253460 278974 255563 278976
rect 255497 278971 255563 278974
rect 66805 278898 66871 278901
rect 264329 278898 264395 278901
rect 267774 278898 267780 278900
rect 66805 278896 68908 278898
rect 66805 278840 66810 278896
rect 66866 278840 68908 278896
rect 66805 278838 68908 278840
rect 264329 278896 267780 278898
rect 264329 278840 264334 278896
rect 264390 278840 267780 278896
rect 264329 278838 267780 278840
rect 66805 278835 66871 278838
rect 264329 278835 264395 278838
rect 267774 278836 267780 278838
rect 267844 278836 267850 278900
rect 100702 278700 100708 278764
rect 100772 278762 100778 278764
rect 105997 278762 106063 278765
rect 137461 278762 137527 278765
rect 100772 278760 137527 278762
rect 100772 278704 106002 278760
rect 106058 278704 137466 278760
rect 137522 278704 137527 278760
rect 100772 278702 137527 278704
rect 100772 278700 100778 278702
rect 105997 278699 106063 278702
rect 137461 278699 137527 278702
rect 101397 278626 101463 278629
rect 98716 278624 101463 278626
rect 98716 278568 101402 278624
rect 101458 278568 101463 278624
rect 98716 278566 101463 278568
rect 101397 278563 101463 278566
rect 255497 278490 255563 278493
rect 253460 278488 255563 278490
rect 253460 278432 255502 278488
rect 255558 278432 255563 278488
rect 253460 278430 255563 278432
rect 255497 278427 255563 278430
rect 258441 278218 258507 278221
rect 260966 278218 260972 278220
rect 253430 278216 260972 278218
rect 253430 278160 258446 278216
rect 258502 278160 260972 278216
rect 253430 278158 260972 278160
rect 67541 278082 67607 278085
rect 153929 278082 153995 278085
rect 184054 278082 184060 278084
rect 67541 278080 68908 278082
rect 67541 278024 67546 278080
rect 67602 278024 68908 278080
rect 67541 278022 68908 278024
rect 153929 278080 184060 278082
rect 153929 278024 153934 278080
rect 153990 278024 184060 278080
rect 153929 278022 184060 278024
rect 67541 278019 67607 278022
rect 153929 278019 153995 278022
rect 184054 278020 184060 278022
rect 184124 278020 184130 278084
rect 191557 278082 191623 278085
rect 191557 278080 193660 278082
rect 191557 278024 191562 278080
rect 191618 278024 193660 278080
rect 253430 278052 253490 278158
rect 258441 278155 258507 278158
rect 260966 278156 260972 278158
rect 261036 278156 261042 278220
rect 259453 278082 259519 278085
rect 292665 278082 292731 278085
rect 259453 278080 292731 278082
rect 191557 278022 193660 278024
rect 259453 278024 259458 278080
rect 259514 278024 292670 278080
rect 292726 278024 292731 278080
rect 259453 278022 292731 278024
rect 191557 278019 191623 278022
rect 259453 278019 259519 278022
rect 292665 278019 292731 278022
rect 100702 277810 100708 277812
rect 98716 277750 100708 277810
rect 100702 277748 100708 277750
rect 100772 277748 100778 277812
rect 255405 277674 255471 277677
rect 253460 277672 255471 277674
rect 253460 277616 255410 277672
rect 255466 277616 255471 277672
rect 253460 277614 255471 277616
rect 255405 277611 255471 277614
rect 255497 277402 255563 277405
rect 262438 277402 262444 277404
rect 255497 277400 262444 277402
rect 255497 277344 255502 277400
rect 255558 277344 262444 277400
rect 255497 277342 262444 277344
rect 255497 277339 255563 277342
rect 262438 277340 262444 277342
rect 262508 277340 262514 277404
rect 67398 277204 67404 277268
rect 67468 277266 67474 277268
rect 67468 277206 68908 277266
rect 67468 277204 67474 277206
rect 253430 277130 253490 277236
rect 253430 277070 258090 277130
rect 101949 276994 102015 276997
rect 106365 276994 106431 276997
rect 98716 276992 106431 276994
rect 98716 276936 101954 276992
rect 102010 276936 106370 276992
rect 106426 276936 106431 276992
rect 98716 276934 106431 276936
rect 101949 276931 102015 276934
rect 106365 276931 106431 276934
rect 191741 276994 191807 276997
rect 191741 276992 193660 276994
rect 191741 276936 191746 276992
rect 191802 276936 193660 276992
rect 191741 276934 193660 276936
rect 191741 276931 191807 276934
rect 255497 276858 255563 276861
rect 253460 276856 255563 276858
rect 253460 276800 255502 276856
rect 255558 276800 255563 276856
rect 253460 276798 255563 276800
rect 255497 276795 255563 276798
rect 130469 276722 130535 276725
rect 154021 276722 154087 276725
rect 130469 276720 154087 276722
rect 130469 276664 130474 276720
rect 130530 276664 154026 276720
rect 154082 276664 154087 276720
rect 130469 276662 154087 276664
rect 130469 276659 130535 276662
rect 154021 276659 154087 276662
rect 160686 276660 160692 276724
rect 160756 276722 160762 276724
rect 166206 276722 166212 276724
rect 160756 276662 166212 276722
rect 160756 276660 160762 276662
rect 166206 276660 166212 276662
rect 166276 276660 166282 276724
rect 258030 276722 258090 277070
rect 273529 276722 273595 276725
rect 277393 276722 277459 276725
rect 258030 276720 277459 276722
rect 258030 276664 273534 276720
rect 273590 276664 277398 276720
rect 277454 276664 277459 276720
rect 258030 276662 277459 276664
rect 273529 276659 273595 276662
rect 277393 276659 277459 276662
rect 66897 276450 66963 276453
rect 255589 276450 255655 276453
rect 66897 276448 68908 276450
rect 66897 276392 66902 276448
rect 66958 276392 68908 276448
rect 66897 276390 68908 276392
rect 253460 276448 255655 276450
rect 253460 276392 255594 276448
rect 255650 276392 255655 276448
rect 253460 276390 255655 276392
rect 66897 276387 66963 276390
rect 255589 276387 255655 276390
rect 100753 276178 100819 276181
rect 98716 276176 100819 276178
rect 98716 276120 100758 276176
rect 100814 276120 100819 276176
rect 98716 276118 100819 276120
rect 100753 276115 100819 276118
rect 65885 276042 65951 276045
rect 67398 276042 67404 276044
rect 65885 276040 67404 276042
rect 65885 275984 65890 276040
rect 65946 275984 67404 276040
rect 65885 275982 67404 275984
rect 65885 275979 65951 275982
rect 67398 275980 67404 275982
rect 67468 275980 67474 276044
rect 255405 276042 255471 276045
rect 253460 276040 255471 276042
rect 253460 275984 255410 276040
rect 255466 275984 255471 276040
rect 253460 275982 255471 275984
rect 255405 275979 255471 275982
rect 191741 275906 191807 275909
rect 191741 275904 193660 275906
rect 191741 275848 191746 275904
rect 191802 275848 193660 275904
rect 191741 275846 193660 275848
rect 191741 275843 191807 275846
rect 66897 275634 66963 275637
rect 66897 275632 68908 275634
rect 66897 275576 66902 275632
rect 66958 275576 68908 275632
rect 66897 275574 68908 275576
rect 66897 275571 66963 275574
rect 258257 275498 258323 275501
rect 253460 275496 258323 275498
rect 253460 275440 258262 275496
rect 258318 275440 258323 275496
rect 253460 275438 258323 275440
rect 258257 275435 258323 275438
rect 100753 275362 100819 275365
rect 98716 275360 100819 275362
rect 98716 275304 100758 275360
rect 100814 275304 100819 275360
rect 98716 275302 100819 275304
rect 100753 275299 100819 275302
rect 193806 275300 193812 275364
rect 193876 275300 193882 275364
rect 57789 275226 57855 275229
rect 66294 275226 66300 275228
rect 57789 275224 66300 275226
rect 57789 275168 57794 275224
rect 57850 275168 66300 275224
rect 57789 275166 66300 275168
rect 57789 275163 57855 275166
rect 66294 275164 66300 275166
rect 66364 275226 66370 275228
rect 66364 275166 68938 275226
rect 66364 275164 66370 275166
rect 68878 274788 68938 275166
rect 157977 274818 158043 274821
rect 193814 274818 193874 275300
rect 255497 275090 255563 275093
rect 253460 275088 255563 275090
rect 253460 275032 255502 275088
rect 255558 275032 255563 275088
rect 253460 275030 255563 275032
rect 255497 275027 255563 275030
rect 157977 274816 193874 274818
rect 157977 274760 157982 274816
rect 158038 274788 193874 274816
rect 158038 274760 193844 274788
rect 157977 274758 193844 274760
rect 157977 274755 158043 274758
rect 189993 274682 190059 274685
rect 190269 274682 190335 274685
rect 191741 274682 191807 274685
rect 255405 274682 255471 274685
rect 189993 274680 191807 274682
rect 189993 274624 189998 274680
rect 190054 274624 190274 274680
rect 190330 274624 191746 274680
rect 191802 274624 191807 274680
rect 189993 274622 191807 274624
rect 253460 274680 255471 274682
rect 253460 274624 255410 274680
rect 255466 274624 255471 274680
rect 253460 274622 255471 274624
rect 189993 274619 190059 274622
rect 190269 274619 190335 274622
rect 191741 274619 191807 274622
rect 255405 274619 255471 274622
rect 100937 274546 101003 274549
rect 98716 274544 101003 274546
rect 98716 274488 100942 274544
rect 100998 274488 101003 274544
rect 98716 274486 101003 274488
rect 100937 274483 101003 274486
rect 255405 274274 255471 274277
rect 253460 274272 255471 274274
rect 253460 274216 255410 274272
rect 255466 274216 255471 274272
rect 253460 274214 255471 274216
rect 255405 274211 255471 274214
rect 66897 274002 66963 274005
rect 66897 274000 68908 274002
rect 66897 273944 66902 274000
rect 66958 273944 68908 274000
rect 66897 273942 68908 273944
rect 66897 273939 66963 273942
rect 255497 273866 255563 273869
rect 253460 273864 255563 273866
rect 253460 273808 255502 273864
rect 255558 273808 255563 273864
rect 253460 273806 255563 273808
rect 255497 273803 255563 273806
rect 100845 273730 100911 273733
rect 98716 273728 100911 273730
rect 98716 273672 100850 273728
rect 100906 273672 100911 273728
rect 98716 273670 100911 273672
rect 100845 273667 100911 273670
rect 191741 273730 191807 273733
rect 191741 273728 193660 273730
rect 191741 273672 191746 273728
rect 191802 273672 193660 273728
rect 191741 273670 193660 273672
rect 191741 273667 191807 273670
rect 270493 273594 270559 273597
rect 270953 273594 271019 273597
rect 253430 273592 271019 273594
rect 253430 273536 270498 273592
rect 270554 273536 270958 273592
rect 271014 273536 271019 273592
rect 253430 273534 271019 273536
rect 253430 273428 253490 273534
rect 270493 273531 270559 273534
rect 270953 273531 271019 273534
rect 66161 272642 66227 272645
rect 68878 272642 68938 273156
rect 100753 272914 100819 272917
rect 98716 272912 100819 272914
rect 98716 272856 100758 272912
rect 100814 272856 100819 272912
rect 98716 272854 100819 272856
rect 100753 272851 100819 272854
rect 253430 272778 253490 272884
rect 262254 272778 262260 272780
rect 253430 272718 262260 272778
rect 262254 272716 262260 272718
rect 262324 272716 262330 272780
rect 64830 272640 68938 272642
rect 64830 272584 66166 272640
rect 66222 272584 68938 272640
rect 64830 272582 68938 272584
rect 191281 272642 191347 272645
rect 191281 272640 193660 272642
rect 191281 272584 191286 272640
rect 191342 272584 193660 272640
rect 191281 272582 193660 272584
rect 63309 272098 63375 272101
rect 64830 272098 64890 272582
rect 66161 272579 66227 272582
rect 191281 272579 191347 272582
rect 101489 272506 101555 272509
rect 188429 272506 188495 272509
rect 255405 272506 255471 272509
rect 101489 272504 188495 272506
rect 101489 272448 101494 272504
rect 101550 272448 188434 272504
rect 188490 272448 188495 272504
rect 101489 272446 188495 272448
rect 253460 272504 255471 272506
rect 253460 272448 255410 272504
rect 255466 272448 255471 272504
rect 253460 272446 255471 272448
rect 101489 272443 101555 272446
rect 188429 272443 188495 272446
rect 255405 272443 255471 272446
rect 259310 272444 259316 272508
rect 259380 272506 259386 272508
rect 291285 272506 291351 272509
rect 259380 272504 291351 272506
rect 259380 272448 291290 272504
rect 291346 272448 291351 272504
rect 259380 272446 291351 272448
rect 259380 272444 259386 272446
rect 291285 272443 291351 272446
rect 66897 272370 66963 272373
rect 66897 272368 68908 272370
rect 66897 272312 66902 272368
rect 66958 272312 68908 272368
rect 66897 272310 68908 272312
rect 66897 272307 66963 272310
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 100845 272098 100911 272101
rect 255405 272098 255471 272101
rect 63309 272096 64890 272098
rect 63309 272040 63314 272096
rect 63370 272040 64890 272096
rect 63309 272038 64890 272040
rect 98716 272096 100911 272098
rect 98716 272040 100850 272096
rect 100906 272040 100911 272096
rect 98716 272038 100911 272040
rect 253460 272096 255471 272098
rect 253460 272040 255410 272096
rect 255466 272040 255471 272096
rect 583520 272084 584960 272174
rect 253460 272038 255471 272040
rect 63309 272035 63375 272038
rect 100845 272035 100911 272038
rect 255405 272035 255471 272038
rect 191741 271554 191807 271557
rect 253430 271554 253490 271660
rect 262397 271554 262463 271557
rect 191741 271552 193660 271554
rect 68878 271010 68938 271524
rect 191741 271496 191746 271552
rect 191802 271496 193660 271552
rect 191741 271494 193660 271496
rect 253430 271552 262463 271554
rect 253430 271496 262402 271552
rect 262458 271496 262463 271552
rect 253430 271494 262463 271496
rect 191741 271491 191807 271494
rect 262397 271491 262463 271494
rect 101213 271282 101279 271285
rect 98716 271280 101279 271282
rect 98716 271224 101218 271280
rect 101274 271224 101279 271280
rect 98716 271222 101279 271224
rect 101213 271219 101279 271222
rect 145557 271282 145623 271285
rect 178953 271282 179019 271285
rect 255497 271282 255563 271285
rect 145557 271280 179019 271282
rect 145557 271224 145562 271280
rect 145618 271224 178958 271280
rect 179014 271224 179019 271280
rect 145557 271222 179019 271224
rect 253460 271280 255563 271282
rect 253460 271224 255502 271280
rect 255558 271224 255563 271280
rect 253460 271222 255563 271224
rect 145557 271219 145623 271222
rect 178953 271219 179019 271222
rect 255497 271219 255563 271222
rect 114461 271146 114527 271149
rect 149789 271146 149855 271149
rect 114461 271144 149855 271146
rect 114461 271088 114466 271144
rect 114522 271088 149794 271144
rect 149850 271088 149855 271144
rect 114461 271086 149855 271088
rect 114461 271083 114527 271086
rect 149789 271083 149855 271086
rect 262397 271146 262463 271149
rect 273345 271146 273411 271149
rect 262397 271144 273411 271146
rect 262397 271088 262402 271144
rect 262458 271088 273350 271144
rect 273406 271088 273411 271144
rect 262397 271086 273411 271088
rect 262397 271083 262463 271086
rect 273345 271083 273411 271086
rect 64830 270950 68938 271010
rect 53465 270738 53531 270741
rect 64830 270738 64890 270950
rect 258390 270874 258396 270876
rect 253460 270814 258396 270874
rect 258390 270812 258396 270814
rect 258460 270874 258466 270876
rect 259126 270874 259132 270876
rect 258460 270814 259132 270874
rect 258460 270812 258466 270814
rect 259126 270812 259132 270814
rect 259196 270812 259202 270876
rect 53465 270736 64890 270738
rect 53465 270680 53470 270736
rect 53526 270680 64890 270736
rect 53465 270678 64890 270680
rect 66897 270738 66963 270741
rect 66897 270736 68908 270738
rect 66897 270680 66902 270736
rect 66958 270680 68908 270736
rect 66897 270678 68908 270680
rect 53465 270675 53531 270678
rect 66897 270675 66963 270678
rect 99465 270466 99531 270469
rect 100753 270466 100819 270469
rect 98716 270464 100819 270466
rect 98716 270408 99470 270464
rect 99526 270408 100758 270464
rect 100814 270408 100819 270464
rect 98716 270406 100819 270408
rect 99465 270403 99531 270406
rect 100753 270403 100819 270406
rect 191189 270466 191255 270469
rect 191189 270464 193660 270466
rect 191189 270408 191194 270464
rect 191250 270408 193660 270464
rect 191189 270406 193660 270408
rect 191189 270403 191255 270406
rect 253430 270194 253490 270436
rect 266486 270194 266492 270196
rect 253430 270134 266492 270194
rect 266486 270132 266492 270134
rect 266556 270132 266562 270196
rect 66897 269922 66963 269925
rect 255405 269922 255471 269925
rect 66897 269920 68908 269922
rect 66897 269864 66902 269920
rect 66958 269864 68908 269920
rect 66897 269862 68908 269864
rect 253460 269920 255471 269922
rect 253460 269864 255410 269920
rect 255466 269864 255471 269920
rect 253460 269862 255471 269864
rect 66897 269859 66963 269862
rect 255405 269859 255471 269862
rect 98686 269378 98746 269620
rect 255405 269514 255471 269517
rect 253460 269512 255471 269514
rect 253460 269456 255410 269512
rect 255466 269456 255471 269512
rect 253460 269454 255471 269456
rect 255405 269451 255471 269454
rect 108297 269378 108363 269381
rect 98686 269376 108363 269378
rect 98686 269320 108302 269376
rect 108358 269320 108363 269376
rect 98686 269318 108363 269320
rect 108297 269315 108363 269318
rect 193397 269378 193463 269381
rect 193397 269376 193660 269378
rect 193397 269320 193402 269376
rect 193458 269320 193660 269376
rect 193397 269318 193660 269320
rect 193397 269315 193463 269318
rect 266486 269180 266492 269244
rect 266556 269242 266562 269244
rect 269297 269242 269363 269245
rect 266556 269240 269363 269242
rect 266556 269184 269302 269240
rect 269358 269184 269363 269240
rect 266556 269182 269363 269184
rect 266556 269180 266562 269182
rect 269297 269179 269363 269182
rect 68878 268562 68938 269076
rect 162710 269044 162716 269108
rect 162780 269106 162786 269108
rect 169201 269106 169267 269109
rect 256785 269106 256851 269109
rect 271137 269108 271203 269109
rect 271086 269106 271092 269108
rect 162780 269104 169267 269106
rect 162780 269048 169206 269104
rect 169262 269048 169267 269104
rect 162780 269046 169267 269048
rect 253460 269104 256851 269106
rect 253460 269048 256790 269104
rect 256846 269048 256851 269104
rect 253460 269046 256851 269048
rect 271046 269046 271092 269106
rect 271156 269104 271203 269108
rect 271198 269048 271203 269104
rect 162780 269044 162786 269046
rect 169201 269043 169267 269046
rect 256785 269043 256851 269046
rect 271086 269044 271092 269046
rect 271156 269044 271203 269048
rect 271137 269043 271203 269044
rect 100753 268834 100819 268837
rect 98716 268832 100819 268834
rect 98716 268776 100758 268832
rect 100814 268776 100819 268832
rect 98716 268774 100819 268776
rect 100753 268771 100819 268774
rect 259361 268698 259427 268701
rect 253460 268696 259427 268698
rect 253460 268640 259366 268696
rect 259422 268640 259427 268696
rect 253460 268638 259427 268640
rect 259361 268635 259427 268638
rect 64830 268502 68938 268562
rect 50797 268018 50863 268021
rect 64830 268018 64890 268502
rect 98862 268364 98868 268428
rect 98932 268426 98938 268428
rect 154021 268426 154087 268429
rect 98932 268424 154087 268426
rect 98932 268368 154026 268424
rect 154082 268368 154087 268424
rect 98932 268366 154087 268368
rect 98932 268364 98938 268366
rect 154021 268363 154087 268366
rect 269614 268364 269620 268428
rect 269684 268426 269690 268428
rect 287145 268426 287211 268429
rect 269684 268424 287211 268426
rect 269684 268368 287150 268424
rect 287206 268368 287211 268424
rect 269684 268366 287211 268368
rect 269684 268364 269690 268366
rect 287145 268363 287211 268366
rect 66713 268290 66779 268293
rect 191189 268290 191255 268293
rect 255405 268290 255471 268293
rect 66713 268288 68908 268290
rect 66713 268232 66718 268288
rect 66774 268232 68908 268288
rect 66713 268230 68908 268232
rect 191189 268288 193660 268290
rect 191189 268232 191194 268288
rect 191250 268232 193660 268288
rect 191189 268230 193660 268232
rect 253460 268288 255471 268290
rect 253460 268232 255410 268288
rect 255466 268232 255471 268288
rect 253460 268230 255471 268232
rect 66713 268227 66779 268230
rect 191189 268227 191255 268230
rect 255405 268227 255471 268230
rect 99005 268018 99071 268021
rect 50797 268016 64890 268018
rect 50797 267960 50802 268016
rect 50858 267960 64890 268016
rect 98164 268016 99071 268018
rect 98164 267988 99010 268016
rect 50797 267958 64890 267960
rect 98134 267960 99010 267988
rect 99066 267960 99071 268016
rect 98134 267958 99071 267960
rect 50797 267955 50863 267958
rect 98134 267885 98194 267958
rect 99005 267955 99071 267958
rect 98085 267880 98194 267885
rect 255405 267882 255471 267885
rect 98085 267824 98090 267880
rect 98146 267824 98194 267880
rect 98085 267822 98194 267824
rect 253460 267880 255471 267882
rect 253460 267824 255410 267880
rect 255466 267824 255471 267880
rect 253460 267822 255471 267824
rect 98085 267819 98151 267822
rect 255405 267819 255471 267822
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 68878 266930 68938 267444
rect 100753 267202 100819 267205
rect 98716 267200 100819 267202
rect 98716 267144 100758 267200
rect 100814 267144 100819 267200
rect 253430 267202 253490 267444
rect 265249 267202 265315 267205
rect 253430 267200 265315 267202
rect 98716 267142 100819 267144
rect 100753 267139 100819 267142
rect 151077 267066 151143 267069
rect 159950 267066 159956 267068
rect 151077 267064 159956 267066
rect 151077 267008 151082 267064
rect 151138 267008 159956 267064
rect 151077 267006 159956 267008
rect 151077 267003 151143 267006
rect 159950 267004 159956 267006
rect 160020 267004 160026 267068
rect 176101 267066 176167 267069
rect 185761 267066 185827 267069
rect 176101 267064 185827 267066
rect 176101 267008 176106 267064
rect 176162 267008 185766 267064
rect 185822 267008 185827 267064
rect 176101 267006 185827 267008
rect 176101 267003 176167 267006
rect 185761 267003 185827 267006
rect 64830 266870 68938 266930
rect 60733 266522 60799 266525
rect 61694 266522 61700 266524
rect 60733 266520 61700 266522
rect 60733 266464 60738 266520
rect 60794 266464 61700 266520
rect 60733 266462 61700 266464
rect 60733 266459 60799 266462
rect 61694 266460 61700 266462
rect 61764 266522 61770 266524
rect 64830 266522 64890 266870
rect 66897 266658 66963 266661
rect 66897 266656 68908 266658
rect 66897 266600 66902 266656
rect 66958 266600 68908 266656
rect 66897 266598 68908 266600
rect 66897 266595 66963 266598
rect 61764 266462 64890 266522
rect 61764 266460 61770 266462
rect 100753 266386 100819 266389
rect 98716 266384 100819 266386
rect 98716 266328 100758 266384
rect 100814 266328 100819 266384
rect 98716 266326 100819 266328
rect 100753 266323 100819 266326
rect 106089 266386 106155 266389
rect 112437 266386 112503 266389
rect 106089 266384 112503 266386
rect 106089 266328 106094 266384
rect 106150 266328 112442 266384
rect 112498 266328 112503 266384
rect 106089 266326 112503 266328
rect 106089 266323 106155 266326
rect 112437 266323 112503 266326
rect 159950 266324 159956 266388
rect 160020 266386 160026 266388
rect 193630 266386 193690 267172
rect 253430 267144 265254 267200
rect 265310 267144 265315 267200
rect 253430 267142 265315 267144
rect 265249 267139 265315 267142
rect 275277 267202 275343 267205
rect 287094 267202 287100 267204
rect 275277 267200 287100 267202
rect 275277 267144 275282 267200
rect 275338 267144 287100 267200
rect 275277 267142 287100 267144
rect 275277 267139 275343 267142
rect 287094 267140 287100 267142
rect 287164 267140 287170 267204
rect 263358 267004 263364 267068
rect 263428 267066 263434 267068
rect 288525 267066 288591 267069
rect 263428 267064 288591 267066
rect 263428 267008 288530 267064
rect 288586 267008 288591 267064
rect 263428 267006 288591 267008
rect 263428 267004 263434 267006
rect 288525 267003 288591 267006
rect 255405 266930 255471 266933
rect 253460 266928 255471 266930
rect 253460 266872 255410 266928
rect 255466 266872 255471 266928
rect 253460 266870 255471 266872
rect 255405 266867 255471 266870
rect 260925 266522 260991 266525
rect 253460 266520 260991 266522
rect 253460 266464 260930 266520
rect 260986 266464 260991 266520
rect 253460 266462 260991 266464
rect 260925 266459 260991 266462
rect 160020 266326 193690 266386
rect 160020 266324 160026 266326
rect 191557 266114 191623 266117
rect 255313 266114 255379 266117
rect 191557 266112 193660 266114
rect 191557 266056 191562 266112
rect 191618 266056 193660 266112
rect 191557 266054 193660 266056
rect 253460 266112 255379 266114
rect 253460 266056 255318 266112
rect 255374 266056 255379 266112
rect 253460 266054 255379 266056
rect 191557 266051 191623 266054
rect 255313 266051 255379 266054
rect 68878 265298 68938 265812
rect 265249 265706 265315 265709
rect 265617 265706 265683 265709
rect 253460 265704 265683 265706
rect 253460 265648 265254 265704
rect 265310 265648 265622 265704
rect 265678 265648 265683 265704
rect 253460 265646 265683 265648
rect 265249 265643 265315 265646
rect 265617 265643 265683 265646
rect 147121 265570 147187 265573
rect 168414 265570 168420 265572
rect 147121 265568 168420 265570
rect 64830 265238 68938 265298
rect 48129 265026 48195 265029
rect 50705 265026 50771 265029
rect 64830 265026 64890 265238
rect 48129 265024 64890 265026
rect 48129 264968 48134 265024
rect 48190 264968 50710 265024
rect 50766 264968 64890 265024
rect 48129 264966 64890 264968
rect 66253 265026 66319 265029
rect 98686 265026 98746 265540
rect 147121 265512 147126 265568
rect 147182 265512 168420 265568
rect 147121 265510 168420 265512
rect 147121 265507 147187 265510
rect 168414 265508 168420 265510
rect 168484 265508 168490 265572
rect 252829 265570 252895 265573
rect 252829 265568 253490 265570
rect 252829 265512 252834 265568
rect 252890 265512 253490 265568
rect 252829 265510 253490 265512
rect 252829 265507 252895 265510
rect 253430 265298 253490 265510
rect 259126 265508 259132 265572
rect 259196 265570 259202 265572
rect 269389 265570 269455 265573
rect 259196 265568 269455 265570
rect 259196 265512 269394 265568
rect 269450 265512 269455 265568
rect 259196 265510 269455 265512
rect 259196 265508 259202 265510
rect 269389 265507 269455 265510
rect 253841 265298 253907 265301
rect 253430 265296 253907 265298
rect 253430 265268 253846 265296
rect 253460 265240 253846 265268
rect 253902 265240 253907 265296
rect 253460 265238 253907 265240
rect 253841 265235 253907 265238
rect 133137 265026 133203 265029
rect 66253 265024 68908 265026
rect 66253 264968 66258 265024
rect 66314 264968 68908 265024
rect 66253 264966 68908 264968
rect 98686 265024 133203 265026
rect 98686 264968 133142 265024
rect 133198 264968 133203 265024
rect 98686 264966 133203 264968
rect 48129 264963 48195 264966
rect 50705 264963 50771 264966
rect 66253 264963 66319 264966
rect 133137 264963 133203 264966
rect 191741 265026 191807 265029
rect 191741 265024 193660 265026
rect 191741 264968 191746 265024
rect 191802 264968 193660 265024
rect 191741 264966 193660 264968
rect 191741 264963 191807 264966
rect 166390 264828 166396 264892
rect 166460 264890 166466 264892
rect 169753 264890 169819 264893
rect 170305 264890 170371 264893
rect 166460 264888 170371 264890
rect 166460 264832 169758 264888
rect 169814 264832 170310 264888
rect 170366 264832 170371 264888
rect 166460 264830 170371 264832
rect 166460 264828 166466 264830
rect 169753 264827 169819 264830
rect 170305 264827 170371 264830
rect 100937 264754 101003 264757
rect 98716 264752 101003 264754
rect 98716 264696 100942 264752
rect 100998 264696 101003 264752
rect 98716 264694 101003 264696
rect 100937 264691 101003 264694
rect 253430 264618 253490 264860
rect 253430 264558 258090 264618
rect 255497 264346 255563 264349
rect 253460 264344 255563 264346
rect 253460 264288 255502 264344
rect 255558 264288 255563 264344
rect 253460 264286 255563 264288
rect 255497 264283 255563 264286
rect 66253 264210 66319 264213
rect 66253 264208 68908 264210
rect 66253 264152 66258 264208
rect 66314 264152 68908 264208
rect 66253 264150 68908 264152
rect 66253 264147 66319 264150
rect 141366 264148 141372 264212
rect 141436 264210 141442 264212
rect 151169 264210 151235 264213
rect 141436 264208 151235 264210
rect 141436 264152 151174 264208
rect 151230 264152 151235 264208
rect 141436 264150 151235 264152
rect 141436 264148 141442 264150
rect 151169 264147 151235 264150
rect 175774 264148 175780 264212
rect 175844 264210 175850 264212
rect 184749 264210 184815 264213
rect 175844 264208 184815 264210
rect 175844 264152 184754 264208
rect 184810 264152 184815 264208
rect 175844 264150 184815 264152
rect 258030 264210 258090 264558
rect 276289 264346 276355 264349
rect 285949 264346 286015 264349
rect 276289 264344 286015 264346
rect 276289 264288 276294 264344
rect 276350 264288 285954 264344
rect 286010 264288 286015 264344
rect 276289 264286 286015 264288
rect 276289 264283 276355 264286
rect 285949 264283 286015 264286
rect 288433 264210 288499 264213
rect 258030 264208 288499 264210
rect 258030 264152 288438 264208
rect 288494 264152 288499 264208
rect 258030 264150 288499 264152
rect 175844 264148 175850 264150
rect 184749 264147 184815 264150
rect 288433 264147 288499 264150
rect 100753 263938 100819 263941
rect 98716 263936 100819 263938
rect 98716 263880 100758 263936
rect 100814 263880 100819 263936
rect 98716 263878 100819 263880
rect 100753 263875 100819 263878
rect 191741 263938 191807 263941
rect 255405 263938 255471 263941
rect 191741 263936 193660 263938
rect 191741 263880 191746 263936
rect 191802 263880 193660 263936
rect 191741 263878 193660 263880
rect 253460 263936 255471 263938
rect 253460 263880 255410 263936
rect 255466 263880 255471 263936
rect 253460 263878 255471 263880
rect 191741 263875 191807 263878
rect 255405 263875 255471 263878
rect 259126 263604 259132 263668
rect 259196 263666 259202 263668
rect 276289 263666 276355 263669
rect 259196 263664 276355 263666
rect 259196 263608 276294 263664
rect 276350 263608 276355 263664
rect 259196 263606 276355 263608
rect 259196 263604 259202 263606
rect 276289 263603 276355 263606
rect 255497 263530 255563 263533
rect 253460 263528 255563 263530
rect 253460 263472 255502 263528
rect 255558 263472 255563 263528
rect 253460 263470 255563 263472
rect 255497 263467 255563 263470
rect 255681 263530 255747 263533
rect 265934 263530 265940 263532
rect 255681 263528 265940 263530
rect 255681 263472 255686 263528
rect 255742 263472 265940 263528
rect 255681 263470 265940 263472
rect 255681 263467 255747 263470
rect 265934 263468 265940 263470
rect 266004 263468 266010 263532
rect 66253 263394 66319 263397
rect 67449 263394 67515 263397
rect 66253 263392 68908 263394
rect 66253 263336 66258 263392
rect 66314 263336 67454 263392
rect 67510 263336 68908 263392
rect 66253 263334 68908 263336
rect 66253 263331 66319 263334
rect 67449 263331 67515 263334
rect 55029 262850 55095 262853
rect 66345 262850 66411 262853
rect 55029 262848 66411 262850
rect 55029 262792 55034 262848
rect 55090 262792 66350 262848
rect 66406 262792 66411 262848
rect 55029 262790 66411 262792
rect 55029 262787 55095 262790
rect 66345 262787 66411 262790
rect 66253 262578 66319 262581
rect 98686 262578 98746 263092
rect 253430 262986 253490 263092
rect 265934 263060 265940 263124
rect 266004 263122 266010 263124
rect 266537 263122 266603 263125
rect 266004 263120 266603 263122
rect 266004 263064 266542 263120
rect 266598 263064 266603 263120
rect 266004 263062 266603 263064
rect 266004 263060 266010 263062
rect 266537 263059 266603 263062
rect 263685 262986 263751 262989
rect 266302 262986 266308 262988
rect 253430 262984 266308 262986
rect 253430 262928 263690 262984
rect 263746 262928 266308 262984
rect 253430 262926 266308 262928
rect 263685 262923 263751 262926
rect 266302 262924 266308 262926
rect 266372 262924 266378 262988
rect 140129 262850 140195 262853
rect 177982 262850 177988 262852
rect 140129 262848 177988 262850
rect 140129 262792 140134 262848
rect 140190 262792 177988 262848
rect 140129 262790 177988 262792
rect 140129 262787 140195 262790
rect 177982 262788 177988 262790
rect 178052 262788 178058 262852
rect 191741 262850 191807 262853
rect 191741 262848 193660 262850
rect 191741 262792 191746 262848
rect 191802 262792 193660 262848
rect 191741 262790 193660 262792
rect 191741 262787 191807 262790
rect 255681 262714 255747 262717
rect 253460 262712 255747 262714
rect 253460 262656 255686 262712
rect 255742 262656 255747 262712
rect 253460 262654 255747 262656
rect 255681 262651 255747 262654
rect 141601 262578 141667 262581
rect 66253 262576 68908 262578
rect 66253 262520 66258 262576
rect 66314 262520 68908 262576
rect 66253 262518 68908 262520
rect 98686 262576 141667 262578
rect 98686 262520 141606 262576
rect 141662 262520 141667 262576
rect 98686 262518 141667 262520
rect 66253 262515 66319 262518
rect 141601 262515 141667 262518
rect 100661 262306 100727 262309
rect 255405 262306 255471 262309
rect 98716 262304 100727 262306
rect 98716 262248 100666 262304
rect 100722 262248 100727 262304
rect 98716 262246 100727 262248
rect 253460 262304 255471 262306
rect 253460 262248 255410 262304
rect 255466 262248 255471 262304
rect 253460 262246 255471 262248
rect 100661 262243 100727 262246
rect 255405 262243 255471 262246
rect 278313 262170 278379 262173
rect 281574 262170 281580 262172
rect 278313 262168 281580 262170
rect 278313 262112 278318 262168
rect 278374 262112 281580 262168
rect 278313 262110 281580 262112
rect 278313 262107 278379 262110
rect 281574 262108 281580 262110
rect 281644 262108 281650 262172
rect 66253 261762 66319 261765
rect 191557 261762 191623 261765
rect 66253 261760 68908 261762
rect 66253 261704 66258 261760
rect 66314 261704 68908 261760
rect 66253 261702 68908 261704
rect 191557 261760 193660 261762
rect 191557 261704 191562 261760
rect 191618 261704 193660 261760
rect 191557 261702 193660 261704
rect 66253 261699 66319 261702
rect 191557 261699 191623 261702
rect 253430 261626 253490 261868
rect 253430 261566 258090 261626
rect 99281 261490 99347 261493
rect 98716 261488 99347 261490
rect 98716 261460 99286 261488
rect 98686 261432 99286 261460
rect 99342 261432 99347 261488
rect 98686 261430 99347 261432
rect 66345 260948 66411 260949
rect 66294 260946 66300 260948
rect 66218 260886 66300 260946
rect 66364 260946 66411 260948
rect 98085 260946 98151 260949
rect 98686 260946 98746 261430
rect 99281 261427 99347 261430
rect 105486 261428 105492 261492
rect 105556 261490 105562 261492
rect 140221 261490 140287 261493
rect 105556 261488 140287 261490
rect 105556 261432 140226 261488
rect 140282 261432 140287 261488
rect 105556 261430 140287 261432
rect 105556 261428 105562 261430
rect 140221 261427 140287 261430
rect 155217 261490 155283 261493
rect 164325 261490 164391 261493
rect 165521 261490 165587 261493
rect 155217 261488 165587 261490
rect 155217 261432 155222 261488
rect 155278 261432 164330 261488
rect 164386 261432 165526 261488
rect 165582 261432 165587 261488
rect 155217 261430 165587 261432
rect 155217 261427 155283 261430
rect 164325 261427 164391 261430
rect 165521 261427 165587 261430
rect 255497 261354 255563 261357
rect 253460 261352 255563 261354
rect 253460 261296 255502 261352
rect 255558 261296 255563 261352
rect 253460 261294 255563 261296
rect 255497 261291 255563 261294
rect 258030 261218 258090 261566
rect 288617 261490 288683 261493
rect 277350 261488 288683 261490
rect 277350 261432 288622 261488
rect 288678 261432 288683 261488
rect 277350 261430 288683 261432
rect 269062 261218 269068 261220
rect 258030 261158 269068 261218
rect 269062 261156 269068 261158
rect 269132 261156 269138 261220
rect 258574 261020 258580 261084
rect 258644 261082 258650 261084
rect 274725 261082 274791 261085
rect 277350 261082 277410 261430
rect 288617 261427 288683 261430
rect 277894 261292 277900 261356
rect 277964 261354 277970 261356
rect 278313 261354 278379 261357
rect 277964 261352 278379 261354
rect 277964 261296 278318 261352
rect 278374 261296 278379 261352
rect 277964 261294 278379 261296
rect 277964 261292 277970 261294
rect 278313 261291 278379 261294
rect 258644 261080 277410 261082
rect 258644 261024 274730 261080
rect 274786 261024 277410 261080
rect 258644 261022 277410 261024
rect 258644 261020 258650 261022
rect 274725 261019 274791 261022
rect 259126 260946 259132 260948
rect 66364 260944 68908 260946
rect 66406 260888 68908 260944
rect 66294 260884 66300 260886
rect 66364 260886 68908 260888
rect 98085 260944 98746 260946
rect 98085 260888 98090 260944
rect 98146 260888 98746 260944
rect 98085 260886 98746 260888
rect 253460 260886 259132 260946
rect 66364 260884 66411 260886
rect 66345 260883 66411 260884
rect 98085 260883 98151 260886
rect 259126 260884 259132 260886
rect 259196 260884 259202 260948
rect 168189 260812 168255 260813
rect 168189 260808 168236 260812
rect 168300 260810 168306 260812
rect 168189 260752 168194 260808
rect 168189 260748 168236 260752
rect 168300 260750 168346 260810
rect 168300 260748 168306 260750
rect 168189 260747 168255 260748
rect 100845 260674 100911 260677
rect 98716 260672 100911 260674
rect 98716 260616 100850 260672
rect 100906 260616 100911 260672
rect 98716 260614 100911 260616
rect 100845 260611 100911 260614
rect 39941 260130 40007 260133
rect 66294 260130 66300 260132
rect 39941 260128 66300 260130
rect 39941 260072 39946 260128
rect 40002 260072 66300 260128
rect 39941 260070 66300 260072
rect 39941 260067 40007 260070
rect 66294 260068 66300 260070
rect 66364 260068 66370 260132
rect 66989 260130 67055 260133
rect 67265 260130 67331 260133
rect 100937 260130 101003 260133
rect 155401 260130 155467 260133
rect 66989 260128 68908 260130
rect 66989 260072 66994 260128
rect 67050 260072 67270 260128
rect 67326 260072 68908 260128
rect 66989 260070 68908 260072
rect 100937 260128 155467 260130
rect 100937 260072 100942 260128
rect 100998 260072 155406 260128
rect 155462 260072 155467 260128
rect 100937 260070 155467 260072
rect 66989 260067 67055 260070
rect 67265 260067 67331 260070
rect 100937 260067 101003 260070
rect 155401 260067 155467 260070
rect 100753 259858 100819 259861
rect 98716 259856 100819 259858
rect 98716 259800 100758 259856
rect 100814 259800 100819 259856
rect 98716 259798 100819 259800
rect 100753 259795 100819 259798
rect 168230 259796 168236 259860
rect 168300 259858 168306 259860
rect 193630 259858 193690 260644
rect 255405 260538 255471 260541
rect 253460 260536 255471 260538
rect 253460 260480 255410 260536
rect 255466 260480 255471 260536
rect 253460 260478 255471 260480
rect 255405 260475 255471 260478
rect 256417 260130 256483 260133
rect 253460 260128 256483 260130
rect 253460 260072 256422 260128
rect 256478 260072 256483 260128
rect 253460 260070 256483 260072
rect 256417 260067 256483 260070
rect 263593 260130 263659 260133
rect 284334 260130 284340 260132
rect 263593 260128 284340 260130
rect 263593 260072 263598 260128
rect 263654 260072 284340 260128
rect 263593 260070 284340 260072
rect 263593 260067 263659 260070
rect 284334 260068 284340 260070
rect 284404 260068 284410 260132
rect 168300 259798 193690 259858
rect 168300 259796 168306 259798
rect 255405 259722 255471 259725
rect 253460 259720 255471 259722
rect 253460 259664 255410 259720
rect 255466 259664 255471 259720
rect 253460 259662 255471 259664
rect 255405 259659 255471 259662
rect 266445 259724 266511 259725
rect 266445 259720 266492 259724
rect 266556 259722 266562 259724
rect 266445 259664 266450 259720
rect 266445 259660 266492 259664
rect 266556 259662 266602 259722
rect 266556 259660 266562 259662
rect 266445 259659 266511 259660
rect 191741 259586 191807 259589
rect 191741 259584 193660 259586
rect 191741 259528 191746 259584
rect 191802 259528 193660 259584
rect 191741 259526 193660 259528
rect 191741 259523 191807 259526
rect 255497 259314 255563 259317
rect 253460 259312 255563 259314
rect 68185 258770 68251 258773
rect 68878 258770 68938 259284
rect 253460 259256 255502 259312
rect 255558 259256 255563 259312
rect 253460 259254 255563 259256
rect 255497 259251 255563 259254
rect 263542 259178 263548 259180
rect 253430 259118 263548 259178
rect 100753 259042 100819 259045
rect 98716 259040 100819 259042
rect 98716 259012 100758 259040
rect 68185 258768 68938 258770
rect 68185 258712 68190 258768
rect 68246 258712 68938 258768
rect 68185 258710 68938 258712
rect 98686 258984 100758 259012
rect 100814 258984 100819 259040
rect 98686 258982 100819 258984
rect 68185 258707 68251 258710
rect 98686 258501 98746 258982
rect 100753 258979 100819 258982
rect 171777 258906 171843 258909
rect 187550 258906 187556 258908
rect 171777 258904 187556 258906
rect 171777 258848 171782 258904
rect 171838 258848 187556 258904
rect 171777 258846 187556 258848
rect 171777 258843 171843 258846
rect 187550 258844 187556 258846
rect 187620 258844 187626 258908
rect 151169 258770 151235 258773
rect 173014 258770 173020 258772
rect 151169 258768 173020 258770
rect 151169 258712 151174 258768
rect 151230 258712 173020 258768
rect 151169 258710 173020 258712
rect 151169 258707 151235 258710
rect 173014 258708 173020 258710
rect 173084 258708 173090 258772
rect 252829 258770 252895 258773
rect 253430 258770 253490 259118
rect 263542 259116 263548 259118
rect 263612 259116 263618 259180
rect 580717 258906 580783 258909
rect 583520 258906 584960 258996
rect 580717 258904 584960 258906
rect 580717 258848 580722 258904
rect 580778 258848 584960 258904
rect 580717 258846 584960 258848
rect 580717 258843 580783 258846
rect 252829 258768 253490 258770
rect 252829 258712 252834 258768
rect 252890 258712 253490 258768
rect 583520 258756 584960 258846
rect 252829 258710 253490 258712
rect 252829 258707 252895 258710
rect 66621 258498 66687 258501
rect 66621 258496 68908 258498
rect 66621 258440 66626 258496
rect 66682 258440 68908 258496
rect 66621 258438 68908 258440
rect 98637 258496 98746 258501
rect 98637 258440 98642 258496
rect 98698 258440 98746 258496
rect 98637 258438 98746 258440
rect 66621 258435 66687 258438
rect 98637 258435 98703 258438
rect 101673 258226 101739 258229
rect 98716 258224 101739 258226
rect 98716 258168 101678 258224
rect 101734 258168 101739 258224
rect 98716 258166 101739 258168
rect 100526 258093 100586 258166
rect 101673 258163 101739 258166
rect 100526 258088 100635 258093
rect 100526 258032 100574 258088
rect 100630 258032 100635 258088
rect 100526 258030 100635 258032
rect 100569 258027 100635 258030
rect 187550 258028 187556 258092
rect 187620 258028 187626 258092
rect 187558 257954 187618 258028
rect 193630 257954 193690 258468
rect 255589 258362 255655 258365
rect 253460 258360 255655 258362
rect 253460 258304 255594 258360
rect 255650 258304 255655 258360
rect 253460 258302 255655 258304
rect 255589 258299 255655 258302
rect 266445 258090 266511 258093
rect 266445 258088 266554 258090
rect 266445 258032 266450 258088
rect 266506 258032 266554 258088
rect 266445 258027 266554 258032
rect 276422 258028 276428 258092
rect 276492 258028 276498 258092
rect 255405 257954 255471 257957
rect 187558 257894 193690 257954
rect 253460 257952 255471 257954
rect 253460 257896 255410 257952
rect 255466 257896 255471 257952
rect 253460 257894 255471 257896
rect 266494 257954 266554 258027
rect 270718 257954 270724 257956
rect 266494 257894 270724 257954
rect 255405 257891 255471 257894
rect 270718 257892 270724 257894
rect 270788 257954 270794 257956
rect 276430 257954 276490 258028
rect 270788 257894 276490 257954
rect 270788 257892 270794 257894
rect 66253 257682 66319 257685
rect 66253 257680 68908 257682
rect 66253 257624 66258 257680
rect 66314 257624 68908 257680
rect 66253 257622 68908 257624
rect 66253 257619 66319 257622
rect 256877 257546 256943 257549
rect 253460 257544 256943 257546
rect 253460 257488 256882 257544
rect 256938 257488 256943 257544
rect 253460 257486 256943 257488
rect 256877 257483 256943 257486
rect 102041 257410 102107 257413
rect 98716 257408 102107 257410
rect 98716 257352 102046 257408
rect 102102 257352 102107 257408
rect 98716 257350 102107 257352
rect 102041 257347 102107 257350
rect 177297 257410 177363 257413
rect 184790 257410 184796 257412
rect 177297 257408 184796 257410
rect 177297 257352 177302 257408
rect 177358 257352 184796 257408
rect 177297 257350 184796 257352
rect 177297 257347 177363 257350
rect 184790 257348 184796 257350
rect 184860 257348 184866 257412
rect 177798 257212 177804 257276
rect 177868 257274 177874 257276
rect 187049 257274 187115 257277
rect 177868 257272 187115 257274
rect 177868 257216 187054 257272
rect 187110 257216 187115 257272
rect 177868 257214 187115 257216
rect 177868 257212 177874 257214
rect 187049 257211 187115 257214
rect 66662 256804 66668 256868
rect 66732 256866 66738 256868
rect 67357 256866 67423 256869
rect 66732 256864 68908 256866
rect 66732 256808 67362 256864
rect 67418 256808 68908 256864
rect 66732 256806 68908 256808
rect 66732 256804 66738 256806
rect 67357 256803 67423 256806
rect 184790 256668 184796 256732
rect 184860 256730 184866 256732
rect 193630 256730 193690 257380
rect 258574 257138 258580 257140
rect 253460 257078 258580 257138
rect 258574 257076 258580 257078
rect 258644 257076 258650 257140
rect 262765 257138 262831 257141
rect 267958 257138 267964 257140
rect 262765 257136 267964 257138
rect 262765 257080 262770 257136
rect 262826 257080 267964 257136
rect 262765 257078 267964 257080
rect 262765 257075 262831 257078
rect 267958 257076 267964 257078
rect 268028 257076 268034 257140
rect 267958 257002 267964 257004
rect 184860 256670 193690 256730
rect 253430 256942 267964 257002
rect 253430 256700 253490 256942
rect 267958 256940 267964 256942
rect 268028 257002 268034 257004
rect 275277 257002 275343 257005
rect 268028 257000 275343 257002
rect 268028 256944 275282 257000
rect 275338 256944 275343 257000
rect 268028 256942 275343 256944
rect 268028 256940 268034 256942
rect 275277 256939 275343 256942
rect 280337 256730 280403 256733
rect 285622 256730 285628 256732
rect 258030 256728 285628 256730
rect 258030 256672 280342 256728
rect 280398 256672 285628 256728
rect 258030 256670 285628 256672
rect 184860 256668 184866 256670
rect 100753 256594 100819 256597
rect 98716 256592 100819 256594
rect 98716 256536 100758 256592
rect 100814 256536 100819 256592
rect 98716 256534 100819 256536
rect 100753 256531 100819 256534
rect 190637 256322 190703 256325
rect 255405 256322 255471 256325
rect 190637 256320 193660 256322
rect 190637 256264 190642 256320
rect 190698 256264 193660 256320
rect 190637 256262 193660 256264
rect 253460 256320 255471 256322
rect 253460 256264 255410 256320
rect 255466 256264 255471 256320
rect 253460 256262 255471 256264
rect 190637 256259 190703 256262
rect 255405 256259 255471 256262
rect 258030 256186 258090 256670
rect 280337 256667 280403 256670
rect 285622 256668 285628 256670
rect 285692 256668 285698 256732
rect 253430 256126 258090 256186
rect 66897 256050 66963 256053
rect 66897 256048 68908 256050
rect 66897 255992 66902 256048
rect 66958 255992 68908 256048
rect 66897 255990 68908 255992
rect 66897 255987 66963 255990
rect 39849 255914 39915 255917
rect 46841 255914 46907 255917
rect 39849 255912 46907 255914
rect 39849 255856 39854 255912
rect 39910 255856 46846 255912
rect 46902 255856 46907 255912
rect 39849 255854 46907 255856
rect 39849 255851 39915 255854
rect 46841 255851 46907 255854
rect 100845 255778 100911 255781
rect 98716 255776 100911 255778
rect 98716 255720 100850 255776
rect 100906 255720 100911 255776
rect 253430 255748 253490 256126
rect 266302 255852 266308 255916
rect 266372 255914 266378 255916
rect 280286 255914 280292 255916
rect 266372 255854 280292 255914
rect 266372 255852 266378 255854
rect 280286 255852 280292 255854
rect 280356 255852 280362 255916
rect 98716 255718 100911 255720
rect 100845 255715 100911 255718
rect 255313 255370 255379 255373
rect 253460 255368 255379 255370
rect 253460 255312 255318 255368
rect 255374 255312 255379 255368
rect 253460 255310 255379 255312
rect 255313 255307 255379 255310
rect 66713 255234 66779 255237
rect 66713 255232 68908 255234
rect 66713 255176 66718 255232
rect 66774 255176 68908 255232
rect 66713 255174 68908 255176
rect 66713 255171 66779 255174
rect 66897 254418 66963 254421
rect 98686 254418 98746 254932
rect 108389 254418 108455 254421
rect 193630 254418 193690 255204
rect 255497 254962 255563 254965
rect 253460 254960 255563 254962
rect 253460 254904 255502 254960
rect 255558 254904 255563 254960
rect 253460 254902 255563 254904
rect 255497 254899 255563 254902
rect 255405 254554 255471 254557
rect 253460 254552 255471 254554
rect 253460 254496 255410 254552
rect 255466 254496 255471 254552
rect 253460 254494 255471 254496
rect 255405 254491 255471 254494
rect 66897 254416 68908 254418
rect 66897 254360 66902 254416
rect 66958 254360 68908 254416
rect 66897 254358 68908 254360
rect 98686 254416 108455 254418
rect 98686 254360 108394 254416
rect 108450 254360 108455 254416
rect 98686 254358 108455 254360
rect 66897 254355 66963 254358
rect 108389 254355 108455 254358
rect 180750 254358 193690 254418
rect 170765 254284 170831 254285
rect 170765 254280 170812 254284
rect 170876 254282 170882 254284
rect -960 254146 480 254236
rect 170765 254224 170770 254280
rect 170765 254220 170812 254224
rect 170876 254222 170922 254282
rect 170876 254220 170882 254222
rect 170765 254219 170831 254220
rect 3417 254146 3483 254149
rect 100753 254146 100819 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect 98716 254144 100819 254146
rect 98716 254088 100758 254144
rect 100814 254088 100819 254144
rect 98716 254086 100819 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 100753 254083 100819 254086
rect 180057 254010 180123 254013
rect 180609 254010 180675 254013
rect 180750 254010 180810 254358
rect 263501 254282 263567 254285
rect 253430 254280 263567 254282
rect 253430 254224 263506 254280
rect 263562 254224 263567 254280
rect 253430 254222 263567 254224
rect 190637 254146 190703 254149
rect 190637 254144 193660 254146
rect 190637 254088 190642 254144
rect 190698 254088 193660 254144
rect 253430 254116 253490 254222
rect 263501 254219 263567 254222
rect 190637 254086 193660 254088
rect 190637 254083 190703 254086
rect 263593 254012 263659 254013
rect 263542 254010 263548 254012
rect 180057 254008 180810 254010
rect 180057 253952 180062 254008
rect 180118 253952 180614 254008
rect 180670 253952 180810 254008
rect 180057 253950 180810 253952
rect 263502 253950 263548 254010
rect 263612 254008 263659 254012
rect 263654 253952 263659 254008
rect 180057 253947 180123 253950
rect 180609 253947 180675 253950
rect 263542 253948 263548 253950
rect 263612 253948 263659 253952
rect 263593 253947 263659 253948
rect 177614 253812 177620 253876
rect 177684 253874 177690 253876
rect 177684 253814 194058 253874
rect 177684 253812 177690 253814
rect 66897 253602 66963 253605
rect 66897 253600 68908 253602
rect 66897 253544 66902 253600
rect 66958 253544 68908 253600
rect 66897 253542 68908 253544
rect 66897 253539 66963 253542
rect 104249 253330 104315 253333
rect 98716 253328 104315 253330
rect 98716 253272 104254 253328
rect 104310 253272 104315 253328
rect 98716 253270 104315 253272
rect 104249 253267 104315 253270
rect 66161 252786 66227 252789
rect 66621 252786 66687 252789
rect 66161 252784 68908 252786
rect 66161 252728 66166 252784
rect 66222 252728 66626 252784
rect 66682 252728 68908 252784
rect 66161 252726 68908 252728
rect 66161 252723 66227 252726
rect 66621 252723 66687 252726
rect 191649 252650 191715 252653
rect 193998 252652 194058 253814
rect 254025 253738 254091 253741
rect 253460 253736 254091 253738
rect 253460 253680 254030 253736
rect 254086 253680 254091 253736
rect 253460 253678 254091 253680
rect 254025 253675 254091 253678
rect 255405 253330 255471 253333
rect 253460 253328 255471 253330
rect 253460 253272 255410 253328
rect 255466 253272 255471 253328
rect 253460 253270 255471 253272
rect 255405 253267 255471 253270
rect 262254 253268 262260 253332
rect 262324 253330 262330 253332
rect 262489 253330 262555 253333
rect 263358 253330 263364 253332
rect 262324 253328 263364 253330
rect 262324 253272 262494 253328
rect 262550 253272 263364 253328
rect 262324 253270 263364 253272
rect 262324 253268 262330 253270
rect 262489 253267 262555 253270
rect 263358 253268 263364 253270
rect 263428 253268 263434 253332
rect 256417 253194 256483 253197
rect 262438 253194 262444 253196
rect 256417 253192 262444 253194
rect 256417 253136 256422 253192
rect 256478 253136 262444 253192
rect 256417 253134 262444 253136
rect 256417 253131 256483 253134
rect 262438 253132 262444 253134
rect 262508 253194 262514 253196
rect 296805 253194 296871 253197
rect 262508 253192 296871 253194
rect 262508 253136 296810 253192
rect 296866 253136 296871 253192
rect 262508 253134 296871 253136
rect 262508 253132 262514 253134
rect 296805 253131 296871 253134
rect 258390 252786 258396 252788
rect 253460 252726 258396 252786
rect 258390 252724 258396 252726
rect 258460 252724 258466 252788
rect 191782 252650 191788 252652
rect 191649 252648 191788 252650
rect 191649 252592 191654 252648
rect 191710 252592 191788 252648
rect 191649 252590 191788 252592
rect 191649 252587 191715 252590
rect 191782 252588 191788 252590
rect 191852 252588 191858 252652
rect 193990 252588 193996 252652
rect 194060 252588 194066 252652
rect 100937 252514 101003 252517
rect 253933 252514 253999 252517
rect 582465 252514 582531 252517
rect 98716 252512 101003 252514
rect 98716 252456 100942 252512
rect 100998 252456 101003 252512
rect 98716 252454 101003 252456
rect 100937 252451 101003 252454
rect 253430 252512 582531 252514
rect 253430 252456 253938 252512
rect 253994 252456 582470 252512
rect 582526 252456 582531 252512
rect 253430 252454 582531 252456
rect 253430 252348 253490 252454
rect 253933 252451 253999 252454
rect 582465 252451 582531 252454
rect 66621 251970 66687 251973
rect 156597 251970 156663 251973
rect 163446 251970 163452 251972
rect 66621 251968 68908 251970
rect 66621 251912 66626 251968
rect 66682 251912 68908 251968
rect 66621 251910 68908 251912
rect 156597 251968 163452 251970
rect 156597 251912 156602 251968
rect 156658 251912 163452 251968
rect 156597 251910 163452 251912
rect 66621 251907 66687 251910
rect 156597 251907 156663 251910
rect 163446 251908 163452 251910
rect 163516 251970 163522 251972
rect 164141 251970 164207 251973
rect 163516 251968 164207 251970
rect 163516 251912 164146 251968
rect 164202 251912 164207 251968
rect 163516 251910 164207 251912
rect 163516 251908 163522 251910
rect 164141 251907 164207 251910
rect 191741 251970 191807 251973
rect 255405 251970 255471 251973
rect 191741 251968 193660 251970
rect 191741 251912 191746 251968
rect 191802 251912 193660 251968
rect 191741 251910 193660 251912
rect 253460 251968 255471 251970
rect 253460 251912 255410 251968
rect 255466 251912 255471 251968
rect 253460 251910 255471 251912
rect 191741 251907 191807 251910
rect 255405 251907 255471 251910
rect 266302 251908 266308 251972
rect 266372 251970 266378 251972
rect 266445 251970 266511 251973
rect 266372 251968 266511 251970
rect 266372 251912 266450 251968
rect 266506 251912 266511 251968
rect 266372 251910 266511 251912
rect 266372 251908 266378 251910
rect 266445 251907 266511 251910
rect 179270 251772 179276 251836
rect 179340 251834 179346 251836
rect 188337 251834 188403 251837
rect 179340 251832 188403 251834
rect 179340 251776 188342 251832
rect 188398 251776 188403 251832
rect 179340 251774 188403 251776
rect 179340 251772 179346 251774
rect 188337 251771 188403 251774
rect 98318 251292 98378 251668
rect 255497 251562 255563 251565
rect 253460 251560 255563 251562
rect 253460 251504 255502 251560
rect 255558 251504 255563 251560
rect 253460 251502 255563 251504
rect 255497 251499 255563 251502
rect 98310 251228 98316 251292
rect 98380 251228 98386 251292
rect 66253 251154 66319 251157
rect 100937 251154 101003 251157
rect 101254 251154 101260 251156
rect 66253 251152 68908 251154
rect 66253 251096 66258 251152
rect 66314 251096 68908 251152
rect 66253 251094 68908 251096
rect 100937 251152 101260 251154
rect 100937 251096 100942 251152
rect 100998 251096 101260 251152
rect 100937 251094 101260 251096
rect 66253 251091 66319 251094
rect 100937 251091 101003 251094
rect 101254 251092 101260 251094
rect 101324 251154 101330 251156
rect 122097 251154 122163 251157
rect 101324 251152 122163 251154
rect 101324 251096 122102 251152
rect 122158 251096 122163 251152
rect 101324 251094 122163 251096
rect 101324 251092 101330 251094
rect 122097 251091 122163 251094
rect 168414 251092 168420 251156
rect 168484 251154 168490 251156
rect 169201 251154 169267 251157
rect 169569 251154 169635 251157
rect 255497 251154 255563 251157
rect 168484 251152 169635 251154
rect 168484 251096 169206 251152
rect 169262 251096 169574 251152
rect 169630 251096 169635 251152
rect 168484 251094 169635 251096
rect 253460 251152 255563 251154
rect 253460 251096 255502 251152
rect 255558 251096 255563 251152
rect 253460 251094 255563 251096
rect 168484 251092 168490 251094
rect 169201 251091 169267 251094
rect 169569 251091 169635 251094
rect 255497 251091 255563 251094
rect 100753 250882 100819 250885
rect 98716 250880 100819 250882
rect 98716 250824 100758 250880
rect 100814 250824 100819 250880
rect 98716 250822 100819 250824
rect 100753 250819 100819 250822
rect 191557 250882 191623 250885
rect 191557 250880 193660 250882
rect 191557 250824 191562 250880
rect 191618 250824 193660 250880
rect 191557 250822 193660 250824
rect 191557 250819 191623 250822
rect 255405 250746 255471 250749
rect 253460 250744 255471 250746
rect 253460 250688 255410 250744
rect 255466 250688 255471 250744
rect 253460 250686 255471 250688
rect 255405 250683 255471 250686
rect 155718 250412 155724 250476
rect 155788 250474 155794 250476
rect 168465 250474 168531 250477
rect 288525 250474 288591 250477
rect 304257 250474 304323 250477
rect 155788 250472 168531 250474
rect 155788 250416 168470 250472
rect 168526 250416 168531 250472
rect 155788 250414 168531 250416
rect 155788 250412 155794 250414
rect 168465 250411 168531 250414
rect 277350 250472 304323 250474
rect 277350 250416 288530 250472
rect 288586 250416 304262 250472
rect 304318 250416 304323 250472
rect 277350 250414 304323 250416
rect 59169 250066 59235 250069
rect 68878 250066 68938 250308
rect 101489 250066 101555 250069
rect 59169 250064 68938 250066
rect 59169 250008 59174 250064
rect 59230 250008 68938 250064
rect 59169 250006 68938 250008
rect 98716 250064 101555 250066
rect 98716 250008 101494 250064
rect 101550 250008 101555 250064
rect 98716 250006 101555 250008
rect 253430 250066 253490 250308
rect 258390 250066 258396 250068
rect 253430 250006 258396 250066
rect 59169 250003 59235 250006
rect 101489 250003 101555 250006
rect 258390 250004 258396 250006
rect 258460 250066 258466 250068
rect 259310 250066 259316 250068
rect 258460 250006 259316 250066
rect 258460 250004 258466 250006
rect 259310 250004 259316 250006
rect 259380 250004 259386 250068
rect 255405 249930 255471 249933
rect 277350 249930 277410 250414
rect 288525 250411 288591 250414
rect 304257 250411 304323 250414
rect 255405 249928 277410 249930
rect 255405 249872 255410 249928
rect 255466 249872 277410 249928
rect 255405 249870 277410 249872
rect 255405 249867 255471 249870
rect 191649 249794 191715 249797
rect 255589 249794 255655 249797
rect 191649 249792 193660 249794
rect 191649 249736 191654 249792
rect 191710 249736 193660 249792
rect 191649 249734 193660 249736
rect 253460 249792 255655 249794
rect 253460 249736 255594 249792
rect 255650 249736 255655 249792
rect 253460 249734 255655 249736
rect 191649 249731 191715 249734
rect 255589 249731 255655 249734
rect 67817 249522 67883 249525
rect 67817 249520 68908 249522
rect 67817 249464 67822 249520
rect 67878 249464 68908 249520
rect 67817 249462 68908 249464
rect 67817 249459 67883 249462
rect 255497 249386 255563 249389
rect 253460 249384 255563 249386
rect 253460 249328 255502 249384
rect 255558 249328 255563 249384
rect 253460 249326 255563 249328
rect 255497 249323 255563 249326
rect 99373 249250 99439 249253
rect 98716 249248 99439 249250
rect 98716 249192 99378 249248
rect 99434 249192 99439 249248
rect 98716 249190 99439 249192
rect 99373 249187 99439 249190
rect 166809 249114 166875 249117
rect 193438 249114 193444 249116
rect 166809 249112 193444 249114
rect 166809 249056 166814 249112
rect 166870 249056 193444 249112
rect 166809 249054 193444 249056
rect 166809 249051 166875 249054
rect 193438 249052 193444 249054
rect 193508 249052 193514 249116
rect 255405 248978 255471 248981
rect 253460 248976 255471 248978
rect 253460 248920 255410 248976
rect 255466 248920 255471 248976
rect 253460 248918 255471 248920
rect 255405 248915 255471 248918
rect 66897 248706 66963 248709
rect 66897 248704 68908 248706
rect 66897 248648 66902 248704
rect 66958 248648 68908 248704
rect 66897 248646 68908 248648
rect 66897 248643 66963 248646
rect 100845 248434 100911 248437
rect 98716 248432 100911 248434
rect 98716 248376 100850 248432
rect 100906 248376 100911 248432
rect 98716 248374 100911 248376
rect 100845 248371 100911 248374
rect 166758 248372 166764 248436
rect 166828 248434 166834 248436
rect 193630 248434 193690 248676
rect 166828 248374 193690 248434
rect 253430 248434 253490 248540
rect 255405 248434 255471 248437
rect 253430 248432 255471 248434
rect 253430 248376 255410 248432
rect 255466 248376 255471 248432
rect 253430 248374 255471 248376
rect 166828 248372 166834 248374
rect 255405 248371 255471 248374
rect 255497 248162 255563 248165
rect 253460 248160 255563 248162
rect 253460 248104 255502 248160
rect 255558 248104 255563 248160
rect 253460 248102 255563 248104
rect 255497 248099 255563 248102
rect 66621 247890 66687 247893
rect 66621 247888 68908 247890
rect 66621 247832 66626 247888
rect 66682 247832 68908 247888
rect 66621 247830 68908 247832
rect 66621 247827 66687 247830
rect 181989 247754 182055 247757
rect 192334 247754 192340 247756
rect 181989 247752 192340 247754
rect 181989 247696 181994 247752
rect 182050 247696 192340 247752
rect 181989 247694 192340 247696
rect 181989 247691 182055 247694
rect 192334 247692 192340 247694
rect 192404 247692 192410 247756
rect 113909 247618 113975 247621
rect 179413 247618 179479 247621
rect 191741 247618 191807 247621
rect 113909 247616 180810 247618
rect 98134 247212 98194 247588
rect 113909 247560 113914 247616
rect 113970 247560 179418 247616
rect 179474 247560 180810 247616
rect 113909 247558 180810 247560
rect 113909 247555 113975 247558
rect 179413 247555 179479 247558
rect 180750 247482 180810 247558
rect 191741 247616 193660 247618
rect 191741 247560 191746 247616
rect 191802 247560 193660 247616
rect 191741 247558 193660 247560
rect 191741 247555 191807 247558
rect 191782 247482 191788 247484
rect 180750 247422 191788 247482
rect 191782 247420 191788 247422
rect 191852 247420 191858 247484
rect 253430 247482 253490 247724
rect 272517 247482 272583 247485
rect 253430 247480 272583 247482
rect 253430 247424 272522 247480
rect 272578 247424 272583 247480
rect 253430 247422 272583 247424
rect 272517 247419 272583 247422
rect 98126 247148 98132 247212
rect 98196 247148 98202 247212
rect 255497 247210 255563 247213
rect 253460 247208 255563 247210
rect 253460 247152 255502 247208
rect 255558 247152 255563 247208
rect 253460 247150 255563 247152
rect 255497 247147 255563 247150
rect 67357 247074 67423 247077
rect 272517 247074 272583 247077
rect 274582 247074 274588 247076
rect 67357 247072 68908 247074
rect 67357 247016 67362 247072
rect 67418 247016 68908 247072
rect 67357 247014 68908 247016
rect 272517 247072 274588 247074
rect 272517 247016 272522 247072
rect 272578 247016 274588 247072
rect 272517 247014 274588 247016
rect 67357 247011 67423 247014
rect 272517 247011 272583 247014
rect 274582 247012 274588 247014
rect 274652 247012 274658 247076
rect 101581 246802 101647 246805
rect 255681 246802 255747 246805
rect 98716 246800 101647 246802
rect 98716 246744 101586 246800
rect 101642 246744 101647 246800
rect 98716 246742 101647 246744
rect 253460 246800 255747 246802
rect 253460 246744 255686 246800
rect 255742 246744 255747 246800
rect 253460 246742 255747 246744
rect 101581 246739 101647 246742
rect 255681 246739 255747 246742
rect 67449 246258 67515 246261
rect 159357 246258 159423 246261
rect 171041 246258 171107 246261
rect 67449 246256 68908 246258
rect 67449 246200 67454 246256
rect 67510 246200 68908 246256
rect 67449 246198 68908 246200
rect 159357 246256 171150 246258
rect 159357 246200 159362 246256
rect 159418 246200 171046 246256
rect 171102 246200 171150 246256
rect 159357 246198 171150 246200
rect 67449 246195 67515 246198
rect 159357 246195 159423 246198
rect 171041 246195 171150 246198
rect 101029 245986 101095 245989
rect 98716 245984 101095 245986
rect 98716 245928 101034 245984
rect 101090 245928 101095 245984
rect 98716 245926 101095 245928
rect 101029 245923 101095 245926
rect 171090 245714 171150 246195
rect 193630 245714 193690 246500
rect 257286 246394 257292 246396
rect 253460 246334 257292 246394
rect 257286 246332 257292 246334
rect 257356 246332 257362 246396
rect 257521 246394 257587 246397
rect 263593 246394 263659 246397
rect 257521 246392 263659 246394
rect 257521 246336 257526 246392
rect 257582 246336 263598 246392
rect 263654 246336 263659 246392
rect 257521 246334 263659 246336
rect 257521 246331 257587 246334
rect 263593 246331 263659 246334
rect 255497 246258 255563 246261
rect 263869 246258 263935 246261
rect 272149 246258 272215 246261
rect 255497 246256 272215 246258
rect 255497 246200 255502 246256
rect 255558 246200 263874 246256
rect 263930 246200 272154 246256
rect 272210 246200 272215 246256
rect 255497 246198 272215 246200
rect 255497 246195 255563 246198
rect 263869 246195 263935 246198
rect 272149 246195 272215 246198
rect 255589 245986 255655 245989
rect 253460 245984 255655 245986
rect 253460 245928 255594 245984
rect 255650 245928 255655 245984
rect 253460 245926 255655 245928
rect 255589 245923 255655 245926
rect 171090 245654 193690 245714
rect 255497 245578 255563 245581
rect 253460 245576 255563 245578
rect 253460 245520 255502 245576
rect 255558 245520 255563 245576
rect 253460 245518 255563 245520
rect 255497 245515 255563 245518
rect 582465 245578 582531 245581
rect 583520 245578 584960 245668
rect 582465 245576 584960 245578
rect 582465 245520 582470 245576
rect 582526 245520 584960 245576
rect 582465 245518 584960 245520
rect 582465 245515 582531 245518
rect 65926 245380 65932 245444
rect 65996 245442 66002 245444
rect 65996 245382 68908 245442
rect 583520 245428 584960 245518
rect 65996 245380 66002 245382
rect 100845 245170 100911 245173
rect 98716 245168 100911 245170
rect 98716 245112 100850 245168
rect 100906 245112 100911 245168
rect 98716 245110 100911 245112
rect 100845 245107 100911 245110
rect 113817 244898 113883 244901
rect 187693 244898 187759 244901
rect 113817 244896 187759 244898
rect 113817 244840 113822 244896
rect 113878 244840 187698 244896
rect 187754 244840 187759 244896
rect 113817 244838 187759 244840
rect 113817 244835 113883 244838
rect 187693 244835 187759 244838
rect 187049 244626 187115 244629
rect 193630 244626 193690 245412
rect 255681 245170 255747 245173
rect 253460 245168 255747 245170
rect 253460 245112 255686 245168
rect 255742 245112 255747 245168
rect 253460 245110 255747 245112
rect 255681 245107 255747 245110
rect 255589 244762 255655 244765
rect 253460 244760 255655 244762
rect 253460 244704 255594 244760
rect 255650 244704 255655 244760
rect 253460 244702 255655 244704
rect 255589 244699 255655 244702
rect 187049 244624 193690 244626
rect 69062 244357 69122 244596
rect 187049 244568 187054 244624
rect 187110 244568 193690 244624
rect 187049 244566 193690 244568
rect 187049 244563 187115 244566
rect 188337 244490 188403 244493
rect 188337 244488 193690 244490
rect 188337 244432 188342 244488
rect 188398 244432 193690 244488
rect 188337 244430 193690 244432
rect 188337 244427 188403 244430
rect 69013 244352 69122 244357
rect 100937 244354 101003 244357
rect 69013 244296 69018 244352
rect 69074 244296 69122 244352
rect 69013 244294 69122 244296
rect 98716 244352 101003 244354
rect 98716 244296 100942 244352
rect 100998 244296 101003 244352
rect 193630 244324 193690 244430
rect 98716 244294 101003 244296
rect 69013 244291 69079 244294
rect 100937 244291 101003 244294
rect 255497 244218 255563 244221
rect 253460 244216 255563 244218
rect 253460 244160 255502 244216
rect 255558 244160 255563 244216
rect 253460 244158 255563 244160
rect 255497 244155 255563 244158
rect 66529 243810 66595 243813
rect 66529 243808 68908 243810
rect 66529 243752 66534 243808
rect 66590 243752 68908 243808
rect 66529 243750 68908 243752
rect 66529 243747 66595 243750
rect 253430 243674 253490 243780
rect 255773 243674 255839 243677
rect 277485 243676 277551 243677
rect 270534 243674 270540 243676
rect 253430 243672 270540 243674
rect 253430 243616 255778 243672
rect 255834 243616 270540 243672
rect 253430 243614 270540 243616
rect 255773 243611 255839 243614
rect 270534 243612 270540 243614
rect 270604 243612 270610 243676
rect 277485 243672 277532 243676
rect 277596 243674 277602 243676
rect 277485 243616 277490 243672
rect 277485 243612 277532 243616
rect 277596 243614 277642 243674
rect 277596 243612 277602 243614
rect 277485 243611 277551 243612
rect 100845 243538 100911 243541
rect 98716 243536 100911 243538
rect 98716 243480 100850 243536
rect 100906 243480 100911 243536
rect 98716 243478 100911 243480
rect 100845 243475 100911 243478
rect 255589 243538 255655 243541
rect 271965 243538 272031 243541
rect 255589 243536 272031 243538
rect 255589 243480 255594 243536
rect 255650 243480 271970 243536
rect 272026 243480 272031 243536
rect 255589 243478 272031 243480
rect 255589 243475 255655 243478
rect 271965 243475 272031 243478
rect 191741 243266 191807 243269
rect 252878 243268 252938 243372
rect 191741 243264 193660 243266
rect 191741 243208 191746 243264
rect 191802 243208 193660 243264
rect 191741 243206 193660 243208
rect 191741 243203 191807 243206
rect 252870 243204 252876 243268
rect 252940 243266 252946 243268
rect 252940 243206 253858 243266
rect 252940 243204 252946 243206
rect 66897 242994 66963 242997
rect 66897 242992 68908 242994
rect 66897 242936 66902 242992
rect 66958 242936 68908 242992
rect 66897 242934 68908 242936
rect 66897 242931 66963 242934
rect 252878 242861 252938 242964
rect 183277 242858 183343 242861
rect 193673 242858 193739 242861
rect 183277 242856 193739 242858
rect 183277 242800 183282 242856
rect 183338 242800 193678 242856
rect 193734 242800 193739 242856
rect 183277 242798 193739 242800
rect 183277 242795 183343 242798
rect 193673 242795 193739 242798
rect 252829 242856 252938 242861
rect 252829 242800 252834 242856
rect 252890 242800 252938 242856
rect 252829 242798 252938 242800
rect 253798 242858 253858 243206
rect 287053 242858 287119 242861
rect 253798 242856 287119 242858
rect 253798 242800 287058 242856
rect 287114 242800 287119 242856
rect 253798 242798 287119 242800
rect 252829 242795 252895 242798
rect 287053 242795 287119 242798
rect 100845 242722 100911 242725
rect 98716 242720 100911 242722
rect 98716 242664 100850 242720
rect 100906 242664 100911 242720
rect 98716 242662 100911 242664
rect 100845 242659 100911 242662
rect 184197 242722 184263 242725
rect 184933 242722 184999 242725
rect 184197 242720 184999 242722
rect 184197 242664 184202 242720
rect 184258 242664 184938 242720
rect 184994 242664 184999 242720
rect 184197 242662 184999 242664
rect 184197 242659 184263 242662
rect 184933 242659 184999 242662
rect 98177 242586 98243 242589
rect 98177 242584 142170 242586
rect 98177 242528 98182 242584
rect 98238 242528 142170 242584
rect 98177 242526 142170 242528
rect 98177 242523 98243 242526
rect 66897 242178 66963 242181
rect 142110 242178 142170 242526
rect 252878 242453 252938 242556
rect 252878 242448 252987 242453
rect 252878 242392 252926 242448
rect 252982 242392 252987 242448
rect 252878 242390 252987 242392
rect 252921 242387 252987 242390
rect 156045 242178 156111 242181
rect 172053 242178 172119 242181
rect 255589 242178 255655 242181
rect 66897 242176 68908 242178
rect 66897 242120 66902 242176
rect 66958 242120 68908 242176
rect 66897 242118 68908 242120
rect 142110 242176 172119 242178
rect 142110 242120 156050 242176
rect 156106 242120 172058 242176
rect 172114 242120 172119 242176
rect 253460 242176 255655 242178
rect 142110 242118 172119 242120
rect 66897 242115 66963 242118
rect 156045 242115 156111 242118
rect 172053 242115 172119 242118
rect 105629 241906 105695 241909
rect 98716 241904 105695 241906
rect 98716 241848 105634 241904
rect 105690 241848 105695 241904
rect 98716 241846 105695 241848
rect 105629 241843 105695 241846
rect 68686 241708 68692 241772
rect 68756 241770 68762 241772
rect 69841 241770 69907 241773
rect 70945 241772 71011 241773
rect 68756 241768 69907 241770
rect 68756 241712 69846 241768
rect 69902 241712 69907 241768
rect 68756 241710 69907 241712
rect 68756 241708 68762 241710
rect 69841 241707 69907 241710
rect 70894 241708 70900 241772
rect 70964 241770 71011 241772
rect 90357 241770 90423 241773
rect 91502 241770 91508 241772
rect 70964 241768 71056 241770
rect 71006 241712 71056 241768
rect 70964 241710 71056 241712
rect 90357 241768 91508 241770
rect 90357 241712 90362 241768
rect 90418 241712 91508 241768
rect 90357 241710 91508 241712
rect 70964 241708 71011 241710
rect 70945 241707 71011 241708
rect 90357 241707 90423 241710
rect 91502 241708 91508 241710
rect 91572 241708 91578 241772
rect 82721 241634 82787 241637
rect 84694 241634 84700 241636
rect 82721 241632 84700 241634
rect 82721 241576 82726 241632
rect 82782 241576 84700 241632
rect 82721 241574 84700 241576
rect 82721 241571 82787 241574
rect 84694 241572 84700 241574
rect 84764 241572 84770 241636
rect 184197 241634 184263 241637
rect 193630 241634 193690 242148
rect 253460 242120 255594 242176
rect 255650 242120 255655 242176
rect 253460 242118 255655 242120
rect 255589 242115 255655 242118
rect 197854 241980 197860 242044
rect 197924 242042 197930 242044
rect 198089 242042 198155 242045
rect 242985 242044 243051 242045
rect 242934 242042 242940 242044
rect 197924 242040 198155 242042
rect 197924 241984 198094 242040
rect 198150 241984 198155 242040
rect 197924 241982 198155 241984
rect 242894 241982 242940 242042
rect 243004 242040 243051 242044
rect 243046 241984 243051 242040
rect 197924 241980 197930 241982
rect 198089 241979 198155 241982
rect 242934 241980 242940 241982
rect 243004 241980 243051 241984
rect 242985 241979 243051 241980
rect 250161 242042 250227 242045
rect 251030 242042 251036 242044
rect 250161 242040 251036 242042
rect 250161 241984 250166 242040
rect 250222 241984 251036 242040
rect 250161 241982 251036 241984
rect 250161 241979 250227 241982
rect 251030 241980 251036 241982
rect 251100 241980 251106 242044
rect 255497 241770 255563 241773
rect 253460 241768 255563 241770
rect 253460 241712 255502 241768
rect 255558 241712 255563 241768
rect 253460 241710 255563 241712
rect 255497 241707 255563 241710
rect 184197 241632 193690 241634
rect 184197 241576 184202 241632
rect 184258 241576 193690 241632
rect 184197 241574 193690 241576
rect 184197 241571 184263 241574
rect 68829 241500 68895 241501
rect 68829 241498 68876 241500
rect 68784 241496 68876 241498
rect 68784 241440 68834 241496
rect 68784 241438 68876 241440
rect 68829 241436 68876 241438
rect 68940 241436 68946 241500
rect 71313 241498 71379 241501
rect 102869 241498 102935 241501
rect 71313 241496 102935 241498
rect 71313 241440 71318 241496
rect 71374 241440 102874 241496
rect 102930 241440 102935 241496
rect 71313 241438 102935 241440
rect 68829 241435 68895 241436
rect 71313 241435 71379 241438
rect 102869 241435 102935 241438
rect 254577 241498 254643 241501
rect 255773 241498 255839 241501
rect 254577 241496 255839 241498
rect 254577 241440 254582 241496
rect 254638 241440 255778 241496
rect 255834 241440 255839 241496
rect 254577 241438 255839 241440
rect 254577 241435 254643 241438
rect 255773 241435 255839 241438
rect 60457 241362 60523 241365
rect 81801 241362 81867 241365
rect 84326 241362 84332 241364
rect 60457 241360 64890 241362
rect 60457 241304 60462 241360
rect 60518 241304 64890 241360
rect 60457 241302 64890 241304
rect 60457 241299 60523 241302
rect 64830 241226 64890 241302
rect 81801 241360 84332 241362
rect 81801 241304 81806 241360
rect 81862 241304 84332 241360
rect 81801 241302 84332 241304
rect 81801 241299 81867 241302
rect 84326 241300 84332 241302
rect 84396 241300 84402 241364
rect 74625 241226 74691 241229
rect 64830 241224 74691 241226
rect -960 241090 480 241180
rect 64830 241168 74630 241224
rect 74686 241168 74691 241224
rect 64830 241166 74691 241168
rect 74625 241163 74691 241166
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 187693 241090 187759 241093
rect 207657 241090 207723 241093
rect 187693 241088 207723 241090
rect 187693 241032 187698 241088
rect 187754 241032 207662 241088
rect 207718 241032 207723 241088
rect 187693 241030 207723 241032
rect 187693 241027 187759 241030
rect 207657 241027 207723 241030
rect 244917 241090 244983 241093
rect 252870 241090 252876 241092
rect 244917 241088 252876 241090
rect 244917 241032 244922 241088
rect 244978 241032 252876 241088
rect 244917 241030 252876 241032
rect 244917 241027 244983 241030
rect 252870 241028 252876 241030
rect 252940 241028 252946 241092
rect 188521 240954 188587 240957
rect 212441 240954 212507 240957
rect 258390 240954 258396 240956
rect 188521 240952 258396 240954
rect 188521 240896 188526 240952
rect 188582 240896 212446 240952
rect 212502 240896 258396 240952
rect 188521 240894 258396 240896
rect 188521 240891 188587 240894
rect 212441 240891 212507 240894
rect 258390 240892 258396 240894
rect 258460 240892 258466 240956
rect 92381 240818 92447 240821
rect 254577 240818 254643 240821
rect 92381 240816 254643 240818
rect 92381 240760 92386 240816
rect 92442 240760 254582 240816
rect 254638 240760 254643 240816
rect 92381 240758 254643 240760
rect 92381 240755 92447 240758
rect 254577 240755 254643 240758
rect 267774 240484 267780 240548
rect 267844 240546 267850 240548
rect 268101 240546 268167 240549
rect 267844 240544 268167 240546
rect 267844 240488 268106 240544
rect 268162 240488 268167 240544
rect 267844 240486 268167 240488
rect 267844 240484 267850 240486
rect 268101 240483 268167 240486
rect 67633 240138 67699 240141
rect 68829 240138 68895 240141
rect 67633 240136 68895 240138
rect 67633 240080 67638 240136
rect 67694 240080 68834 240136
rect 68890 240080 68895 240136
rect 67633 240078 68895 240080
rect 67633 240075 67699 240078
rect 68829 240075 68895 240078
rect 86534 240076 86540 240140
rect 86604 240138 86610 240140
rect 86677 240138 86743 240141
rect 86604 240136 86743 240138
rect 86604 240080 86682 240136
rect 86738 240080 86743 240136
rect 86604 240078 86743 240080
rect 86604 240076 86610 240078
rect 86677 240075 86743 240078
rect 93485 240140 93551 240141
rect 93485 240136 93532 240140
rect 93596 240138 93602 240140
rect 97073 240138 97139 240141
rect 97758 240138 97764 240140
rect 93485 240080 93490 240136
rect 93485 240076 93532 240080
rect 93596 240078 93642 240138
rect 97073 240136 97764 240138
rect 97073 240080 97078 240136
rect 97134 240080 97764 240136
rect 97073 240078 97764 240080
rect 93596 240076 93602 240078
rect 93485 240075 93551 240076
rect 97073 240075 97139 240078
rect 97758 240076 97764 240078
rect 97828 240076 97834 240140
rect 191782 240076 191788 240140
rect 191852 240138 191858 240140
rect 192017 240138 192083 240141
rect 191852 240136 192083 240138
rect 191852 240080 192022 240136
rect 192078 240080 192083 240136
rect 191852 240078 192083 240080
rect 191852 240076 191858 240078
rect 192017 240075 192083 240078
rect 193305 240138 193371 240141
rect 193990 240138 193996 240140
rect 193305 240136 193996 240138
rect 193305 240080 193310 240136
rect 193366 240080 193996 240136
rect 193305 240078 193996 240080
rect 193305 240075 193371 240078
rect 193990 240076 193996 240078
rect 194060 240076 194066 240140
rect 66110 239940 66116 240004
rect 66180 240002 66186 240004
rect 68870 240002 68876 240004
rect 66180 239942 68876 240002
rect 66180 239940 66186 239942
rect 68870 239940 68876 239942
rect 68940 240002 68946 240004
rect 69381 240002 69447 240005
rect 68940 240000 69447 240002
rect 68940 239944 69386 240000
rect 69442 239944 69447 240000
rect 68940 239942 69447 239944
rect 68940 239940 68946 239942
rect 69381 239939 69447 239942
rect 73102 239940 73108 240004
rect 73172 240002 73178 240004
rect 73797 240002 73863 240005
rect 73172 240000 73863 240002
rect 73172 239944 73802 240000
rect 73858 239944 73863 240000
rect 73172 239942 73863 239944
rect 73172 239940 73178 239942
rect 73797 239939 73863 239942
rect 85573 240002 85639 240005
rect 87454 240002 87460 240004
rect 85573 240000 87460 240002
rect 85573 239944 85578 240000
rect 85634 239944 87460 240000
rect 85573 239942 87460 239944
rect 85573 239939 85639 239942
rect 87454 239940 87460 239942
rect 87524 239940 87530 240004
rect 95693 240002 95759 240005
rect 95877 240002 95943 240005
rect 105537 240002 105603 240005
rect 95693 240000 105603 240002
rect 95693 239944 95698 240000
rect 95754 239944 95882 240000
rect 95938 239944 105542 240000
rect 105598 239944 105603 240000
rect 95693 239942 105603 239944
rect 95693 239939 95759 239942
rect 95877 239939 95943 239942
rect 105537 239939 105603 239942
rect 242249 240002 242315 240005
rect 242709 240002 242775 240005
rect 273478 240002 273484 240004
rect 242249 240000 273484 240002
rect 242249 239944 242254 240000
rect 242310 239944 242714 240000
rect 242770 239944 273484 240000
rect 242249 239942 273484 239944
rect 242249 239939 242315 239942
rect 242709 239939 242775 239942
rect 273478 239940 273484 239942
rect 273548 239940 273554 240004
rect 72601 239866 72667 239869
rect 188429 239866 188495 239869
rect 251817 239866 251883 239869
rect 72601 239864 161490 239866
rect 72601 239808 72606 239864
rect 72662 239808 161490 239864
rect 72601 239806 161490 239808
rect 72601 239803 72667 239806
rect 88425 239458 88491 239461
rect 89621 239458 89687 239461
rect 112621 239458 112687 239461
rect 88425 239456 112687 239458
rect 88425 239400 88430 239456
rect 88486 239400 89626 239456
rect 89682 239400 112626 239456
rect 112682 239400 112687 239456
rect 88425 239398 112687 239400
rect 161430 239458 161490 239806
rect 188429 239864 251883 239866
rect 188429 239808 188434 239864
rect 188490 239808 251822 239864
rect 251878 239808 251883 239864
rect 188429 239806 251883 239808
rect 188429 239803 188495 239806
rect 251817 239803 251883 239806
rect 172513 239458 172579 239461
rect 201534 239458 201540 239460
rect 161430 239456 201540 239458
rect 161430 239400 172518 239456
rect 172574 239400 201540 239456
rect 161430 239398 201540 239400
rect 88425 239395 88491 239398
rect 89621 239395 89687 239398
rect 112621 239395 112687 239398
rect 172513 239395 172579 239398
rect 201534 239396 201540 239398
rect 201604 239458 201610 239460
rect 247493 239458 247559 239461
rect 201604 239456 247559 239458
rect 201604 239400 247498 239456
rect 247554 239400 247559 239456
rect 201604 239398 247559 239400
rect 201604 239396 201610 239398
rect 247493 239395 247559 239398
rect 249149 239458 249215 239461
rect 263726 239458 263732 239460
rect 249149 239456 263732 239458
rect 249149 239400 249154 239456
rect 249210 239400 263732 239456
rect 249149 239398 263732 239400
rect 249149 239395 249215 239398
rect 263726 239396 263732 239398
rect 263796 239396 263802 239460
rect 74809 238914 74875 238917
rect 64830 238912 74875 238914
rect 64830 238856 74814 238912
rect 74870 238856 74875 238912
rect 64830 238854 74875 238856
rect 61878 238716 61884 238780
rect 61948 238778 61954 238780
rect 64830 238778 64890 238854
rect 74809 238851 74875 238854
rect 61948 238718 64890 238778
rect 79317 238778 79383 238781
rect 85573 238778 85639 238781
rect 79317 238776 85639 238778
rect 79317 238720 79322 238776
rect 79378 238720 85578 238776
rect 85634 238720 85639 238776
rect 79317 238718 85639 238720
rect 61948 238716 61954 238718
rect 79317 238715 79383 238718
rect 85573 238715 85639 238718
rect 65977 238642 66043 238645
rect 76557 238642 76623 238645
rect 65977 238640 76623 238642
rect 65977 238584 65982 238640
rect 66038 238584 76562 238640
rect 76618 238584 76623 238640
rect 65977 238582 76623 238584
rect 65977 238579 66043 238582
rect 76557 238579 76623 238582
rect 91001 238642 91067 238645
rect 91134 238642 91140 238644
rect 91001 238640 91140 238642
rect 91001 238584 91006 238640
rect 91062 238584 91140 238640
rect 91001 238582 91140 238584
rect 91001 238579 91067 238582
rect 91134 238580 91140 238582
rect 91204 238580 91210 238644
rect 144637 238642 144703 238645
rect 191189 238642 191255 238645
rect 144637 238640 191255 238642
rect 144637 238584 144642 238640
rect 144698 238584 191194 238640
rect 191250 238584 191255 238640
rect 144637 238582 191255 238584
rect 144637 238579 144703 238582
rect 191189 238579 191255 238582
rect 193806 238580 193812 238644
rect 193876 238642 193882 238644
rect 230473 238642 230539 238645
rect 193876 238640 230539 238642
rect 193876 238584 230478 238640
rect 230534 238584 230539 238640
rect 193876 238582 230539 238584
rect 193876 238580 193882 238582
rect 230473 238579 230539 238582
rect 251817 238642 251883 238645
rect 276013 238642 276079 238645
rect 251817 238640 276079 238642
rect 251817 238584 251822 238640
rect 251878 238584 276018 238640
rect 276074 238584 276079 238640
rect 251817 238582 276079 238584
rect 251817 238579 251883 238582
rect 276013 238579 276079 238582
rect 91093 238506 91159 238509
rect 96654 238506 96660 238508
rect 91093 238504 96660 238506
rect 91093 238448 91098 238504
rect 91154 238448 96660 238504
rect 91093 238446 96660 238448
rect 91093 238443 91159 238446
rect 96654 238444 96660 238446
rect 96724 238444 96730 238508
rect 76005 238370 76071 238373
rect 110597 238370 110663 238373
rect 76005 238368 110663 238370
rect 76005 238312 76010 238368
rect 76066 238312 110602 238368
rect 110658 238312 110663 238368
rect 76005 238310 110663 238312
rect 76005 238307 76071 238310
rect 110597 238307 110663 238310
rect 108297 238098 108363 238101
rect 144637 238098 144703 238101
rect 108297 238096 144703 238098
rect 108297 238040 108302 238096
rect 108358 238040 144642 238096
rect 144698 238040 144703 238096
rect 108297 238038 144703 238040
rect 108297 238035 108363 238038
rect 144637 238035 144703 238038
rect 189809 238098 189875 238101
rect 196065 238098 196131 238101
rect 189809 238096 196131 238098
rect 189809 238040 189814 238096
rect 189870 238040 196070 238096
rect 196126 238040 196131 238096
rect 189809 238038 196131 238040
rect 189809 238035 189875 238038
rect 196065 238035 196131 238038
rect 247769 238098 247835 238101
rect 257521 238098 257587 238101
rect 247769 238096 257587 238098
rect 247769 238040 247774 238096
rect 247830 238040 257526 238096
rect 257582 238040 257587 238096
rect 247769 238038 257587 238040
rect 247769 238035 247835 238038
rect 257521 238035 257587 238038
rect 124213 237962 124279 237965
rect 189993 237962 190059 237965
rect 124213 237960 190059 237962
rect 124213 237904 124218 237960
rect 124274 237904 189998 237960
rect 190054 237904 190059 237960
rect 124213 237902 190059 237904
rect 124213 237899 124279 237902
rect 189993 237899 190059 237902
rect 192017 237962 192083 237965
rect 211654 237962 211660 237964
rect 192017 237960 211660 237962
rect 192017 237904 192022 237960
rect 192078 237904 211660 237960
rect 192017 237902 211660 237904
rect 192017 237899 192083 237902
rect 211654 237900 211660 237902
rect 211724 237962 211730 237964
rect 253933 237962 253999 237965
rect 211724 237960 253999 237962
rect 211724 237904 253938 237960
rect 253994 237904 253999 237960
rect 211724 237902 253999 237904
rect 211724 237900 211730 237902
rect 253933 237899 253999 237902
rect 91093 237418 91159 237421
rect 91502 237418 91508 237420
rect 91093 237416 91508 237418
rect 91093 237360 91098 237416
rect 91154 237360 91508 237416
rect 91093 237358 91508 237360
rect 91093 237355 91159 237358
rect 91502 237356 91508 237358
rect 91572 237356 91578 237420
rect 93894 237356 93900 237420
rect 93964 237418 93970 237420
rect 100753 237418 100819 237421
rect 93964 237416 100819 237418
rect 93964 237360 100758 237416
rect 100814 237360 100819 237416
rect 93964 237358 100819 237360
rect 93964 237356 93970 237358
rect 100753 237355 100819 237358
rect 257337 237418 257403 237421
rect 258441 237418 258507 237421
rect 257337 237416 258507 237418
rect 257337 237360 257342 237416
rect 257398 237360 258446 237416
rect 258502 237360 258507 237416
rect 257337 237358 258507 237360
rect 257337 237355 257403 237358
rect 258441 237355 258507 237358
rect 80605 237282 80671 237285
rect 113909 237282 113975 237285
rect 80605 237280 113975 237282
rect 80605 237224 80610 237280
rect 80666 237224 113914 237280
rect 113970 237224 113975 237280
rect 80605 237222 113975 237224
rect 80605 237219 80671 237222
rect 113909 237219 113975 237222
rect 246389 236874 246455 236877
rect 252829 236874 252895 236877
rect 246389 236872 252895 236874
rect 246389 236816 246394 236872
rect 246450 236816 252834 236872
rect 252890 236816 252895 236872
rect 246389 236814 252895 236816
rect 246389 236811 246455 236814
rect 252829 236811 252895 236814
rect 73470 236676 73476 236740
rect 73540 236738 73546 236740
rect 79409 236738 79475 236741
rect 73540 236736 79475 236738
rect 73540 236680 79414 236736
rect 79470 236680 79475 236736
rect 73540 236678 79475 236680
rect 73540 236676 73546 236678
rect 79409 236675 79475 236678
rect 92289 236738 92355 236741
rect 95182 236738 95188 236740
rect 92289 236736 95188 236738
rect 92289 236680 92294 236736
rect 92350 236680 95188 236736
rect 92289 236678 95188 236680
rect 92289 236675 92355 236678
rect 95182 236676 95188 236678
rect 95252 236676 95258 236740
rect 178861 236738 178927 236741
rect 178861 236736 238770 236738
rect 178861 236680 178866 236736
rect 178922 236680 238770 236736
rect 178861 236678 238770 236680
rect 178861 236675 178927 236678
rect 67909 236602 67975 236605
rect 90357 236602 90423 236605
rect 67909 236600 90423 236602
rect 67909 236544 67914 236600
rect 67970 236544 90362 236600
rect 90418 236544 90423 236600
rect 67909 236542 90423 236544
rect 67909 236539 67975 236542
rect 90357 236539 90423 236542
rect 92381 236602 92447 236605
rect 94262 236602 94268 236604
rect 92381 236600 94268 236602
rect 92381 236544 92386 236600
rect 92442 236544 94268 236600
rect 92381 236542 94268 236544
rect 92381 236539 92447 236542
rect 94262 236540 94268 236542
rect 94332 236540 94338 236604
rect 133137 236602 133203 236605
rect 210417 236602 210483 236605
rect 133137 236600 210483 236602
rect 133137 236544 133142 236600
rect 133198 236544 210422 236600
rect 210478 236544 210483 236600
rect 133137 236542 210483 236544
rect 238710 236602 238770 236678
rect 249885 236602 249951 236605
rect 262438 236602 262444 236604
rect 238710 236600 262444 236602
rect 238710 236544 249890 236600
rect 249946 236544 262444 236600
rect 238710 236542 262444 236544
rect 133137 236539 133203 236542
rect 210417 236539 210483 236542
rect 249885 236539 249951 236542
rect 262438 236540 262444 236542
rect 262508 236540 262514 236604
rect 77937 236058 78003 236061
rect 80605 236058 80671 236061
rect 77937 236056 80671 236058
rect 77937 236000 77942 236056
rect 77998 236000 80610 236056
rect 80666 236000 80671 236056
rect 77937 235998 80671 236000
rect 77937 235995 78003 235998
rect 80605 235995 80671 235998
rect 108389 236058 108455 236061
rect 109033 236058 109099 236061
rect 108389 236056 109099 236058
rect 108389 236000 108394 236056
rect 108450 236000 109038 236056
rect 109094 236000 109099 236056
rect 108389 235998 109099 236000
rect 108389 235995 108455 235998
rect 109033 235995 109099 235998
rect 257286 235996 257292 236060
rect 257356 236058 257362 236060
rect 258257 236058 258323 236061
rect 582649 236058 582715 236061
rect 257356 236056 582715 236058
rect 257356 236000 258262 236056
rect 258318 236000 582654 236056
rect 582710 236000 582715 236056
rect 257356 235998 582715 236000
rect 257356 235996 257362 235998
rect 258257 235995 258323 235998
rect 582649 235995 582715 235998
rect 74809 235922 74875 235925
rect 122189 235922 122255 235925
rect 74809 235920 122255 235922
rect 74809 235864 74814 235920
rect 74870 235864 122194 235920
rect 122250 235864 122255 235920
rect 74809 235862 122255 235864
rect 74809 235859 74875 235862
rect 122189 235859 122255 235862
rect 186221 235922 186287 235925
rect 260925 235922 260991 235925
rect 186221 235920 260991 235922
rect 186221 235864 186226 235920
rect 186282 235864 260930 235920
rect 260986 235864 260991 235920
rect 186221 235862 260991 235864
rect 186221 235859 186287 235862
rect 260925 235859 260991 235862
rect 253933 235786 253999 235789
rect 255405 235786 255471 235789
rect 280153 235786 280219 235789
rect 253933 235784 280219 235786
rect 253933 235728 253938 235784
rect 253994 235728 255410 235784
rect 255466 235728 280158 235784
rect 280214 235728 280219 235784
rect 253933 235726 280219 235728
rect 253933 235723 253999 235726
rect 255405 235723 255471 235726
rect 280153 235723 280219 235726
rect 83273 235378 83339 235381
rect 115197 235378 115263 235381
rect 117957 235378 118023 235381
rect 83273 235376 118023 235378
rect 83273 235320 83278 235376
rect 83334 235320 115202 235376
rect 115258 235320 117962 235376
rect 118018 235320 118023 235376
rect 83273 235318 118023 235320
rect 83273 235315 83339 235318
rect 115197 235315 115263 235318
rect 117957 235315 118023 235318
rect 110413 235242 110479 235245
rect 184381 235242 184447 235245
rect 110413 235240 184447 235242
rect 110413 235184 110418 235240
rect 110474 235184 184386 235240
rect 184442 235184 184447 235240
rect 110413 235182 184447 235184
rect 110413 235179 110479 235182
rect 184381 235179 184447 235182
rect 67449 234562 67515 234565
rect 116761 234562 116827 234565
rect 67449 234560 116827 234562
rect 67449 234504 67454 234560
rect 67510 234504 116766 234560
rect 116822 234504 116827 234560
rect 67449 234502 116827 234504
rect 67449 234499 67515 234502
rect 116761 234499 116827 234502
rect 175181 234562 175247 234565
rect 258390 234562 258396 234564
rect 175181 234560 258396 234562
rect 175181 234504 175186 234560
rect 175242 234504 258396 234560
rect 175181 234502 258396 234504
rect 175181 234499 175247 234502
rect 258390 234500 258396 234502
rect 258460 234500 258466 234564
rect 197353 234426 197419 234429
rect 190410 234424 197419 234426
rect 190410 234368 197358 234424
rect 197414 234368 197419 234424
rect 190410 234366 197419 234368
rect 174721 234154 174787 234157
rect 175181 234154 175247 234157
rect 174721 234152 175247 234154
rect 174721 234096 174726 234152
rect 174782 234096 175186 234152
rect 175242 234096 175247 234152
rect 174721 234094 175247 234096
rect 174721 234091 174787 234094
rect 175181 234091 175247 234094
rect 180885 234154 180951 234157
rect 182081 234154 182147 234157
rect 190410 234154 190470 234366
rect 197353 234363 197419 234366
rect 180885 234152 190470 234154
rect 180885 234096 180890 234152
rect 180946 234096 182086 234152
rect 182142 234096 190470 234152
rect 180885 234094 190470 234096
rect 180885 234091 180951 234094
rect 182081 234091 182147 234094
rect 31753 233882 31819 233885
rect 137829 233882 137895 233885
rect 31753 233880 137895 233882
rect 31753 233824 31758 233880
rect 31814 233824 137834 233880
rect 137890 233824 137895 233880
rect 31753 233822 137895 233824
rect 31753 233819 31819 233822
rect 137829 233819 137895 233822
rect 77569 233202 77635 233205
rect 104157 233202 104223 233205
rect 108389 233202 108455 233205
rect 77569 233200 108455 233202
rect 77569 233144 77574 233200
rect 77630 233144 104162 233200
rect 104218 233144 108394 233200
rect 108450 233144 108455 233200
rect 77569 233142 108455 233144
rect 77569 233139 77635 233142
rect 104157 233139 104223 233142
rect 108389 233139 108455 233142
rect 155309 233202 155375 233205
rect 160686 233202 160692 233204
rect 155309 233200 160692 233202
rect 155309 233144 155314 233200
rect 155370 233144 160692 233200
rect 155309 233142 160692 233144
rect 155309 233139 155375 233142
rect 160686 233140 160692 233142
rect 160756 233140 160762 233204
rect 171869 233202 171935 233205
rect 256877 233202 256943 233205
rect 171869 233200 256943 233202
rect 171869 233144 171874 233200
rect 171930 233144 256882 233200
rect 256938 233144 256943 233200
rect 171869 233142 256943 233144
rect 171869 233139 171935 233142
rect 256877 233139 256943 233142
rect 173341 233066 173407 233069
rect 253933 233066 253999 233069
rect 173341 233064 253999 233066
rect 173341 233008 173346 233064
rect 173402 233008 253938 233064
rect 253994 233008 253999 233064
rect 173341 233006 253999 233008
rect 173341 233003 173407 233006
rect 253933 233003 253999 233006
rect 110505 232658 110571 232661
rect 116025 232658 116091 232661
rect 110505 232656 116091 232658
rect 110505 232600 110510 232656
rect 110566 232600 116030 232656
rect 116086 232600 116091 232656
rect 110505 232598 116091 232600
rect 110505 232595 110571 232598
rect 116025 232595 116091 232598
rect 111057 232522 111123 232525
rect 207013 232522 207079 232525
rect 111057 232520 207079 232522
rect 111057 232464 111062 232520
rect 111118 232464 207018 232520
rect 207074 232464 207079 232520
rect 111057 232462 207079 232464
rect 111057 232459 111123 232462
rect 207013 232459 207079 232462
rect 236637 232522 236703 232525
rect 252093 232522 252159 232525
rect 236637 232520 252159 232522
rect 236637 232464 236642 232520
rect 236698 232464 252098 232520
rect 252154 232464 252159 232520
rect 236637 232462 252159 232464
rect 236637 232459 236703 232462
rect 252093 232459 252159 232462
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 180241 231298 180307 231301
rect 266486 231298 266492 231300
rect 180241 231296 266492 231298
rect 180241 231240 180246 231296
rect 180302 231240 266492 231296
rect 180241 231238 266492 231240
rect 180241 231235 180307 231238
rect 266486 231236 266492 231238
rect 266556 231236 266562 231300
rect 115381 231162 115447 231165
rect 217317 231162 217383 231165
rect 115381 231160 217383 231162
rect 115381 231104 115386 231160
rect 115442 231104 217322 231160
rect 217378 231104 217383 231160
rect 115381 231102 217383 231104
rect 115381 231099 115447 231102
rect 217317 231099 217383 231102
rect 58985 230482 59051 230485
rect 166257 230482 166323 230485
rect 166809 230482 166875 230485
rect 58985 230480 161490 230482
rect 58985 230424 58990 230480
rect 59046 230424 161490 230480
rect 58985 230422 161490 230424
rect 58985 230419 59051 230422
rect 161430 230346 161490 230422
rect 166257 230480 171150 230482
rect 166257 230424 166262 230480
rect 166318 230424 166814 230480
rect 166870 230424 171150 230480
rect 166257 230422 171150 230424
rect 166257 230419 166323 230422
rect 166809 230419 166875 230422
rect 168465 230346 168531 230349
rect 169661 230346 169727 230349
rect 161430 230344 169727 230346
rect 161430 230288 168470 230344
rect 168526 230288 169666 230344
rect 169722 230288 169727 230344
rect 161430 230286 169727 230288
rect 171090 230346 171150 230422
rect 269062 230346 269068 230348
rect 171090 230286 269068 230346
rect 168465 230283 168531 230286
rect 169661 230283 169727 230286
rect 269062 230284 269068 230286
rect 269132 230284 269138 230348
rect 207013 229122 207079 229125
rect 210509 229122 210575 229125
rect 207013 229120 210575 229122
rect 207013 229064 207018 229120
rect 207074 229064 210514 229120
rect 210570 229064 210575 229120
rect 207013 229062 210575 229064
rect 207013 229059 207079 229062
rect 210509 229059 210575 229062
rect 177389 228986 177455 228989
rect 254669 228986 254735 228989
rect 177389 228984 254735 228986
rect 177389 228928 177394 228984
rect 177450 228928 254674 228984
rect 254730 228928 254735 228984
rect 177389 228926 254735 228928
rect 177389 228923 177455 228926
rect 254669 228923 254735 228926
rect 192334 228788 192340 228852
rect 192404 228850 192410 228852
rect 231853 228850 231919 228853
rect 192404 228848 231919 228850
rect 192404 228792 231858 228848
rect 231914 228792 231919 228848
rect 192404 228790 231919 228792
rect 192404 228788 192410 228790
rect 231853 228787 231919 228790
rect 61694 228244 61700 228308
rect 61764 228306 61770 228308
rect 119337 228306 119403 228309
rect 61764 228304 119403 228306
rect 61764 228248 119342 228304
rect 119398 228248 119403 228304
rect 61764 228246 119403 228248
rect 61764 228244 61770 228246
rect 119337 228243 119403 228246
rect -960 227884 480 228124
rect 85481 227762 85547 227765
rect 88742 227762 88748 227764
rect 85481 227760 88748 227762
rect 85481 227704 85486 227760
rect 85542 227704 88748 227760
rect 85481 227702 88748 227704
rect 85481 227699 85547 227702
rect 88742 227700 88748 227702
rect 88812 227700 88818 227764
rect 94078 227700 94084 227764
rect 94148 227762 94154 227764
rect 101254 227762 101260 227764
rect 94148 227702 101260 227762
rect 94148 227700 94154 227702
rect 101254 227700 101260 227702
rect 101324 227700 101330 227764
rect 177389 227762 177455 227765
rect 177941 227762 178007 227765
rect 177389 227760 178007 227762
rect 177389 227704 177394 227760
rect 177450 227704 177946 227760
rect 178002 227704 178007 227760
rect 177389 227702 178007 227704
rect 177389 227699 177455 227702
rect 177941 227699 178007 227702
rect 231853 227762 231919 227765
rect 233141 227762 233207 227765
rect 231853 227760 233207 227762
rect 231853 227704 231858 227760
rect 231914 227704 233146 227760
rect 233202 227704 233207 227760
rect 231853 227702 233207 227704
rect 231853 227699 231919 227702
rect 233141 227699 233207 227702
rect 71446 227564 71452 227628
rect 71516 227626 71522 227628
rect 73245 227626 73311 227629
rect 138657 227626 138723 227629
rect 71516 227624 138723 227626
rect 71516 227568 73250 227624
rect 73306 227568 138662 227624
rect 138718 227568 138723 227624
rect 71516 227566 138723 227568
rect 71516 227564 71522 227566
rect 73245 227563 73311 227566
rect 138657 227563 138723 227566
rect 210417 227626 210483 227629
rect 267958 227626 267964 227628
rect 210417 227624 267964 227626
rect 210417 227568 210422 227624
rect 210478 227568 267964 227624
rect 210417 227566 267964 227568
rect 210417 227563 210483 227566
rect 267958 227564 267964 227566
rect 268028 227564 268034 227628
rect 155401 226946 155467 226949
rect 204897 226946 204963 226949
rect 271873 226946 271939 226949
rect 155401 226944 271939 226946
rect 155401 226888 155406 226944
rect 155462 226888 204902 226944
rect 204958 226888 271878 226944
rect 271934 226888 271939 226944
rect 155401 226886 271939 226888
rect 155401 226883 155467 226886
rect 204897 226883 204963 226886
rect 271873 226883 271939 226886
rect 210417 226402 210483 226405
rect 211061 226402 211127 226405
rect 210417 226400 211127 226402
rect 210417 226344 210422 226400
rect 210478 226344 211066 226400
rect 211122 226344 211127 226400
rect 210417 226342 211127 226344
rect 210417 226339 210483 226342
rect 211061 226339 211127 226342
rect 195973 225586 196039 225589
rect 255313 225586 255379 225589
rect 195973 225584 255379 225586
rect 195973 225528 195978 225584
rect 196034 225528 255318 225584
rect 255374 225528 255379 225584
rect 195973 225526 255379 225528
rect 195973 225523 196039 225526
rect 255313 225523 255379 225526
rect 169661 224906 169727 224909
rect 288525 224906 288591 224909
rect 169661 224904 288591 224906
rect 169661 224848 169666 224904
rect 169722 224848 288530 224904
rect 288586 224848 288591 224904
rect 169661 224846 288591 224848
rect 169661 224843 169727 224846
rect 288525 224843 288591 224846
rect 180333 224226 180399 224229
rect 241421 224226 241487 224229
rect 263869 224226 263935 224229
rect 180333 224224 263935 224226
rect 180333 224168 180338 224224
rect 180394 224168 241426 224224
rect 241482 224168 263874 224224
rect 263930 224168 263935 224224
rect 180333 224166 263935 224168
rect 180333 224163 180399 224166
rect 241421 224163 241487 224166
rect 263869 224163 263935 224166
rect 104249 223546 104315 223549
rect 270718 223546 270724 223548
rect 104249 223544 270724 223546
rect 104249 223488 104254 223544
rect 104310 223488 270724 223544
rect 104249 223486 270724 223488
rect 104249 223483 104315 223486
rect 270718 223484 270724 223486
rect 270788 223484 270794 223548
rect 186957 222186 187023 222189
rect 258257 222186 258323 222189
rect 186957 222184 258323 222186
rect 186957 222128 186962 222184
rect 187018 222128 258262 222184
rect 258318 222128 258323 222184
rect 186957 222126 258323 222128
rect 186957 222123 187023 222126
rect 258257 222123 258323 222126
rect 98126 220900 98132 220964
rect 98196 220962 98202 220964
rect 252553 220962 252619 220965
rect 98196 220960 252619 220962
rect 98196 220904 252558 220960
rect 252614 220904 252619 220960
rect 98196 220902 252619 220904
rect 98196 220900 98202 220902
rect 252553 220899 252619 220902
rect 164141 220826 164207 220829
rect 236637 220826 236703 220829
rect 164141 220824 236703 220826
rect 164141 220768 164146 220824
rect 164202 220768 236642 220824
rect 236698 220768 236703 220824
rect 164141 220766 236703 220768
rect 164141 220763 164207 220766
rect 236637 220763 236703 220766
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 82813 217970 82879 217973
rect 186957 217970 187023 217973
rect 82813 217968 187023 217970
rect 82813 217912 82818 217968
rect 82874 217912 186962 217968
rect 187018 217912 187023 217968
rect 82813 217910 187023 217912
rect 82813 217907 82879 217910
rect 186957 217907 187023 217910
rect 217317 217970 217383 217973
rect 244917 217970 244983 217973
rect 217317 217968 244983 217970
rect 217317 217912 217322 217968
rect 217378 217912 244922 217968
rect 244978 217912 244983 217968
rect 217317 217910 244983 217912
rect 217317 217907 217383 217910
rect 244917 217907 244983 217910
rect 186313 216746 186379 216749
rect 186957 216746 187023 216749
rect 186313 216744 187023 216746
rect 186313 216688 186318 216744
rect 186374 216688 186962 216744
rect 187018 216688 187023 216744
rect 186313 216686 187023 216688
rect 186313 216683 186379 216686
rect 186957 216683 187023 216686
rect 213177 216746 213243 216749
rect 215334 216746 215340 216748
rect 213177 216744 215340 216746
rect 213177 216688 213182 216744
rect 213238 216688 215340 216744
rect 213177 216686 215340 216688
rect 213177 216683 213243 216686
rect 215334 216684 215340 216686
rect 215404 216684 215410 216748
rect 2773 215930 2839 215933
rect 188470 215930 188476 215932
rect 2773 215928 188476 215930
rect 2773 215872 2778 215928
rect 2834 215872 188476 215928
rect 2773 215870 188476 215872
rect 2773 215867 2839 215870
rect 188470 215868 188476 215870
rect 188540 215868 188546 215932
rect 196617 215930 196683 215933
rect 205582 215930 205588 215932
rect 196617 215928 205588 215930
rect 196617 215872 196622 215928
rect 196678 215872 205588 215928
rect 196617 215870 205588 215872
rect 196617 215867 196683 215870
rect 205582 215868 205588 215870
rect 205652 215868 205658 215932
rect -960 214978 480 215068
rect 3969 214978 4035 214981
rect -960 214976 4035 214978
rect -960 214920 3974 214976
rect 4030 214920 4035 214976
rect -960 214918 4035 214920
rect -960 214828 480 214918
rect 3969 214915 4035 214918
rect 97942 214508 97948 214572
rect 98012 214570 98018 214572
rect 98821 214570 98887 214573
rect 266721 214570 266787 214573
rect 98012 214568 266787 214570
rect 98012 214512 98826 214568
rect 98882 214512 266726 214568
rect 266782 214512 266787 214568
rect 98012 214510 266787 214512
rect 98012 214508 98018 214510
rect 98821 214507 98887 214510
rect 266721 214507 266787 214510
rect 92974 213148 92980 213212
rect 93044 213210 93050 213212
rect 93526 213210 93532 213212
rect 93044 213150 93532 213210
rect 93044 213148 93050 213150
rect 93526 213148 93532 213150
rect 93596 213210 93602 213212
rect 273437 213210 273503 213213
rect 93596 213208 273503 213210
rect 93596 213152 273442 213208
rect 273498 213152 273503 213208
rect 93596 213150 273503 213152
rect 93596 213148 93602 213150
rect 273437 213147 273503 213150
rect 235993 210354 236059 210357
rect 267774 210354 267780 210356
rect 235993 210352 267780 210354
rect 235993 210296 235998 210352
rect 236054 210296 267780 210352
rect 235993 210294 267780 210296
rect 235993 210291 236059 210294
rect 267774 210292 267780 210294
rect 267844 210292 267850 210356
rect 153837 208314 153903 208317
rect 219566 208314 219572 208316
rect 153837 208312 219572 208314
rect 153837 208256 153842 208312
rect 153898 208256 219572 208312
rect 153837 208254 219572 208256
rect 153837 208251 153903 208254
rect 219566 208252 219572 208254
rect 219636 208314 219642 208316
rect 220077 208314 220143 208317
rect 219636 208312 220143 208314
rect 219636 208256 220082 208312
rect 220138 208256 220143 208312
rect 219636 208254 220143 208256
rect 219636 208252 219642 208254
rect 220077 208251 220143 208254
rect 117313 206274 117379 206277
rect 185577 206274 185643 206277
rect 117313 206272 185643 206274
rect 117313 206216 117318 206272
rect 117374 206216 185582 206272
rect 185638 206216 185643 206272
rect 117313 206214 185643 206216
rect 117313 206211 117379 206214
rect 185577 206211 185643 206214
rect 260925 205730 260991 205733
rect 262070 205730 262076 205732
rect 260925 205728 262076 205730
rect 260925 205672 260930 205728
rect 260986 205672 262076 205728
rect 260925 205670 262076 205672
rect 260925 205667 260991 205670
rect 262070 205668 262076 205670
rect 262140 205668 262146 205732
rect 580349 205730 580415 205733
rect 583520 205730 584960 205820
rect 580349 205728 584960 205730
rect 580349 205672 580354 205728
rect 580410 205672 584960 205728
rect 580349 205670 584960 205672
rect 580349 205667 580415 205670
rect 166206 205532 166212 205596
rect 166276 205594 166282 205596
rect 302233 205594 302299 205597
rect 166276 205592 302299 205594
rect 166276 205536 302238 205592
rect 302294 205536 302299 205592
rect 583520 205580 584960 205670
rect 166276 205534 302299 205536
rect 166276 205532 166282 205534
rect 302233 205531 302299 205534
rect 97758 204308 97764 204372
rect 97828 204370 97834 204372
rect 104985 204370 105051 204373
rect 258165 204370 258231 204373
rect 258717 204370 258783 204373
rect 97828 204368 258783 204370
rect 97828 204312 104990 204368
rect 105046 204312 258170 204368
rect 258226 204312 258722 204368
rect 258778 204312 258783 204368
rect 97828 204310 258783 204312
rect 97828 204308 97834 204310
rect 104985 204307 105051 204310
rect 258165 204307 258231 204310
rect 258717 204307 258783 204310
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 214649 200698 214715 200701
rect 242934 200698 242940 200700
rect 214649 200696 242940 200698
rect 214649 200640 214654 200696
rect 214710 200640 242940 200696
rect 214649 200638 242940 200640
rect 214649 200635 214715 200638
rect 242934 200636 242940 200638
rect 243004 200636 243010 200700
rect 66110 199276 66116 199340
rect 66180 199338 66186 199340
rect 180241 199338 180307 199341
rect 66180 199336 180307 199338
rect 66180 199280 180246 199336
rect 180302 199280 180307 199336
rect 66180 199278 180307 199280
rect 66180 199276 66186 199278
rect 180241 199275 180307 199278
rect 188838 199276 188844 199340
rect 188908 199338 188914 199340
rect 246389 199338 246455 199341
rect 188908 199336 246455 199338
rect 188908 199280 246394 199336
rect 246450 199280 246455 199336
rect 188908 199278 246455 199280
rect 188908 199276 188914 199278
rect 246389 199275 246455 199278
rect 197353 193898 197419 193901
rect 262254 193898 262260 193900
rect 197353 193896 262260 193898
rect 197353 193840 197358 193896
rect 197414 193840 262260 193896
rect 197353 193838 262260 193840
rect 197353 193835 197419 193838
rect 262254 193836 262260 193838
rect 262324 193836 262330 193900
rect 104014 192476 104020 192540
rect 104084 192538 104090 192540
rect 123569 192538 123635 192541
rect 104084 192536 123635 192538
rect 104084 192480 123574 192536
rect 123630 192480 123635 192536
rect 104084 192478 123635 192480
rect 104084 192476 104090 192478
rect 123569 192475 123635 192478
rect 211797 192538 211863 192541
rect 263542 192538 263548 192540
rect 211797 192536 263548 192538
rect 211797 192480 211802 192536
rect 211858 192480 263548 192536
rect 211797 192478 263548 192480
rect 211797 192475 211863 192478
rect 263542 192476 263548 192478
rect 263612 192476 263618 192540
rect 579981 192538 580047 192541
rect 583520 192538 584960 192628
rect 579981 192536 584960 192538
rect 579981 192480 579986 192536
rect 580042 192480 584960 192536
rect 579981 192478 584960 192480
rect 579981 192475 580047 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 42793 188322 42859 188325
rect 168414 188322 168420 188324
rect 42793 188320 168420 188322
rect 42793 188264 42798 188320
rect 42854 188264 168420 188320
rect 42793 188262 168420 188264
rect 42793 188259 42859 188262
rect 168414 188260 168420 188262
rect 168484 188260 168490 188324
rect 86534 185540 86540 185604
rect 86604 185602 86610 185604
rect 120073 185602 120139 185605
rect 86604 185600 120139 185602
rect 86604 185544 120078 185600
rect 120134 185544 120139 185600
rect 86604 185542 120139 185544
rect 86604 185540 86610 185542
rect 120073 185539 120139 185542
rect 153837 185602 153903 185605
rect 188286 185602 188292 185604
rect 153837 185600 188292 185602
rect 153837 185544 153842 185600
rect 153898 185544 188292 185600
rect 153837 185542 188292 185544
rect 153837 185539 153903 185542
rect 188286 185540 188292 185542
rect 188356 185540 188362 185604
rect 188286 181324 188292 181388
rect 188356 181386 188362 181388
rect 277894 181386 277900 181388
rect 188356 181326 277900 181386
rect 188356 181324 188362 181326
rect 277894 181324 277900 181326
rect 277964 181324 277970 181388
rect 192477 180026 192543 180029
rect 200614 180026 200620 180028
rect 192477 180024 200620 180026
rect 192477 179968 192482 180024
rect 192538 179968 200620 180024
rect 192477 179966 200620 179968
rect 192477 179963 192543 179966
rect 200614 179964 200620 179966
rect 200684 179964 200690 180028
rect 63217 179482 63283 179485
rect 188286 179482 188292 179484
rect 63217 179480 188292 179482
rect 63217 179424 63222 179480
rect 63278 179424 188292 179480
rect 63217 179422 188292 179424
rect 63217 179419 63283 179422
rect 188286 179420 188292 179422
rect 188356 179420 188362 179484
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 93669 176764 93735 176765
rect 93669 176760 93716 176764
rect 93780 176762 93786 176764
rect 93669 176704 93674 176760
rect 93669 176700 93716 176704
rect 93780 176702 93826 176762
rect 93780 176700 93786 176702
rect 93669 176699 93735 176700
rect -960 175796 480 176036
rect 86309 175810 86375 175813
rect 86718 175810 86724 175812
rect 86309 175808 86724 175810
rect 86309 175752 86314 175808
rect 86370 175752 86724 175808
rect 86309 175750 86724 175752
rect 86309 175747 86375 175750
rect 86718 175748 86724 175750
rect 86788 175748 86794 175812
rect 86309 175402 86375 175405
rect 210417 175402 210483 175405
rect 86309 175400 210483 175402
rect 86309 175344 86314 175400
rect 86370 175344 210422 175400
rect 210478 175344 210483 175400
rect 86309 175342 210483 175344
rect 86309 175339 86375 175342
rect 210417 175339 210483 175342
rect 193857 174586 193923 174589
rect 255313 174586 255379 174589
rect 193857 174584 255379 174586
rect 193857 174528 193862 174584
rect 193918 174528 255318 174584
rect 255374 174528 255379 174584
rect 193857 174526 255379 174528
rect 193857 174523 193923 174526
rect 255313 174523 255379 174526
rect 86217 172546 86283 172549
rect 217317 172546 217383 172549
rect 86217 172544 217383 172546
rect 86217 172488 86222 172544
rect 86278 172488 217322 172544
rect 217378 172488 217383 172544
rect 86217 172486 217383 172488
rect 86217 172483 86283 172486
rect 217317 172483 217383 172486
rect 209129 171730 209195 171733
rect 226425 171730 226491 171733
rect 209129 171728 226491 171730
rect 209129 171672 209134 171728
rect 209190 171672 226430 171728
rect 226486 171672 226491 171728
rect 209129 171670 226491 171672
rect 209129 171667 209195 171670
rect 226425 171667 226491 171670
rect 142981 169826 143047 169829
rect 235993 169826 236059 169829
rect 142981 169824 236059 169826
rect 142981 169768 142986 169824
rect 143042 169768 235998 169824
rect 236054 169768 236059 169824
rect 142981 169766 236059 169768
rect 142981 169763 143047 169766
rect 235993 169763 236059 169766
rect 196801 169010 196867 169013
rect 216673 169010 216739 169013
rect 196801 169008 216739 169010
rect 196801 168952 196806 169008
rect 196862 168952 216678 169008
rect 216734 168952 216739 169008
rect 196801 168950 216739 168952
rect 196801 168947 196867 168950
rect 216673 168947 216739 168950
rect 89713 167106 89779 167109
rect 219433 167106 219499 167109
rect 220169 167106 220235 167109
rect 89713 167104 220235 167106
rect 89713 167048 89718 167104
rect 89774 167048 219438 167104
rect 219494 167048 220174 167104
rect 220230 167048 220235 167104
rect 89713 167046 220235 167048
rect 89713 167043 89779 167046
rect 219433 167043 219499 167046
rect 220169 167043 220235 167046
rect 200113 166970 200179 166973
rect 200665 166970 200731 166973
rect 266302 166970 266308 166972
rect 200113 166968 266308 166970
rect 200113 166912 200118 166968
rect 200174 166912 200670 166968
rect 200726 166912 266308 166968
rect 200113 166910 266308 166912
rect 200113 166907 200179 166910
rect 200665 166907 200731 166910
rect 266302 166908 266308 166910
rect 266372 166908 266378 166972
rect 582833 165882 582899 165885
rect 583520 165882 584960 165972
rect 582833 165880 584960 165882
rect 582833 165824 582838 165880
rect 582894 165824 584960 165880
rect 582833 165822 584960 165824
rect 582833 165819 582899 165822
rect 76649 165746 76715 165749
rect 192477 165746 192543 165749
rect 76649 165744 192543 165746
rect 76649 165688 76654 165744
rect 76710 165688 192482 165744
rect 192538 165688 192543 165744
rect 583520 165732 584960 165822
rect 76649 165686 192543 165688
rect 76649 165683 76715 165686
rect 192477 165683 192543 165686
rect 153929 164386 153995 164389
rect 237373 164386 237439 164389
rect 153929 164384 237439 164386
rect 153929 164328 153934 164384
rect 153990 164328 237378 164384
rect 237434 164328 237439 164384
rect 153929 164326 237439 164328
rect 153929 164323 153995 164326
rect 237373 164323 237439 164326
rect 75177 163434 75243 163437
rect 95182 163434 95188 163436
rect 75177 163432 95188 163434
rect 75177 163376 75182 163432
rect 75238 163376 95188 163432
rect 75177 163374 95188 163376
rect 75177 163371 75243 163374
rect 95182 163372 95188 163374
rect 95252 163372 95258 163436
rect -960 162890 480 162980
rect 2865 162890 2931 162893
rect -960 162888 2931 162890
rect -960 162832 2870 162888
rect 2926 162832 2931 162888
rect -960 162830 2931 162832
rect -960 162740 480 162830
rect 2865 162827 2931 162830
rect 105537 162890 105603 162893
rect 229093 162890 229159 162893
rect 105537 162888 229159 162890
rect 105537 162832 105542 162888
rect 105598 162832 229098 162888
rect 229154 162832 229159 162888
rect 105537 162830 229159 162832
rect 105537 162827 105603 162830
rect 229093 162827 229159 162830
rect 208393 162754 208459 162757
rect 270493 162754 270559 162757
rect 208393 162752 270559 162754
rect 208393 162696 208398 162752
rect 208454 162696 270498 162752
rect 270554 162696 270559 162752
rect 208393 162694 270559 162696
rect 208393 162691 208459 162694
rect 270493 162691 270559 162694
rect 181989 162210 182055 162213
rect 190453 162210 190519 162213
rect 181989 162208 190519 162210
rect 181989 162152 181994 162208
rect 182050 162152 190458 162208
rect 190514 162152 190519 162208
rect 181989 162150 190519 162152
rect 181989 162147 182055 162150
rect 190453 162147 190519 162150
rect 74717 162074 74783 162077
rect 166809 162074 166875 162077
rect 185761 162074 185827 162077
rect 74717 162072 185827 162074
rect 74717 162016 74722 162072
rect 74778 162016 166814 162072
rect 166870 162016 185766 162072
rect 185822 162016 185827 162072
rect 74717 162014 185827 162016
rect 74717 162011 74783 162014
rect 166809 162011 166875 162014
rect 185761 162011 185827 162014
rect 193121 162074 193187 162077
rect 230473 162074 230539 162077
rect 193121 162072 230539 162074
rect 193121 162016 193126 162072
rect 193182 162016 230478 162072
rect 230534 162016 230539 162072
rect 193121 162014 230539 162016
rect 193121 162011 193187 162014
rect 230473 162011 230539 162014
rect 63309 160714 63375 160717
rect 157333 160714 157399 160717
rect 63309 160712 157399 160714
rect 63309 160656 63314 160712
rect 63370 160656 157338 160712
rect 157394 160656 157399 160712
rect 63309 160654 157399 160656
rect 63309 160651 63375 160654
rect 157333 160651 157399 160654
rect 157333 160306 157399 160309
rect 158069 160306 158135 160309
rect 157333 160304 158135 160306
rect 157333 160248 157338 160304
rect 157394 160248 158074 160304
rect 158130 160248 158135 160304
rect 157333 160246 158135 160248
rect 157333 160243 157399 160246
rect 158069 160243 158135 160246
rect 140129 160170 140195 160173
rect 249885 160170 249951 160173
rect 140129 160168 249951 160170
rect 140129 160112 140134 160168
rect 140190 160112 249890 160168
rect 249946 160112 249951 160168
rect 140129 160110 249951 160112
rect 140129 160107 140195 160110
rect 249885 160107 249951 160110
rect 61745 159354 61811 159357
rect 191833 159354 191899 159357
rect 192569 159354 192635 159357
rect 61745 159352 192635 159354
rect 61745 159296 61750 159352
rect 61806 159296 191838 159352
rect 191894 159296 192574 159352
rect 192630 159296 192635 159352
rect 61745 159294 192635 159296
rect 61745 159291 61811 159294
rect 191833 159291 191899 159294
rect 192569 159291 192635 159294
rect 61745 158810 61811 158813
rect 61929 158810 61995 158813
rect 61745 158808 61995 158810
rect 61745 158752 61750 158808
rect 61806 158752 61934 158808
rect 61990 158752 61995 158808
rect 61745 158750 61995 158752
rect 61745 158747 61811 158750
rect 61929 158747 61995 158750
rect 211889 158810 211955 158813
rect 212441 158810 212507 158813
rect 230473 158810 230539 158813
rect 211889 158808 230539 158810
rect 211889 158752 211894 158808
rect 211950 158752 212446 158808
rect 212502 158752 230478 158808
rect 230534 158752 230539 158808
rect 211889 158750 230539 158752
rect 211889 158747 211955 158750
rect 212441 158747 212507 158750
rect 230473 158747 230539 158750
rect 200205 157994 200271 157997
rect 288433 157994 288499 157997
rect 200205 157992 288499 157994
rect 200205 157936 200210 157992
rect 200266 157936 288438 157992
rect 288494 157936 288499 157992
rect 200205 157934 288499 157936
rect 200205 157931 200271 157934
rect 288433 157931 288499 157934
rect 92749 157450 92815 157453
rect 223573 157450 223639 157453
rect 224769 157450 224835 157453
rect 92749 157448 224835 157450
rect 92749 157392 92754 157448
rect 92810 157392 223578 157448
rect 223634 157392 224774 157448
rect 224830 157392 224835 157448
rect 92749 157390 224835 157392
rect 92749 157387 92815 157390
rect 223573 157387 223639 157390
rect 224769 157387 224835 157390
rect 178861 156226 178927 156229
rect 207657 156226 207723 156229
rect 178861 156224 207723 156226
rect 178861 156168 178866 156224
rect 178922 156168 207662 156224
rect 207718 156168 207723 156224
rect 178861 156166 207723 156168
rect 178861 156163 178927 156166
rect 207657 156163 207723 156166
rect 145649 156090 145715 156093
rect 259545 156090 259611 156093
rect 145649 156088 259611 156090
rect 145649 156032 145654 156088
rect 145710 156032 259550 156088
rect 259606 156032 259611 156088
rect 145649 156030 259611 156032
rect 145649 156027 145715 156030
rect 259545 156027 259611 156030
rect 210417 155954 210483 155957
rect 294045 155954 294111 155957
rect 294689 155954 294755 155957
rect 210417 155952 294755 155954
rect 210417 155896 210422 155952
rect 210478 155896 294050 155952
rect 294106 155896 294694 155952
rect 294750 155896 294755 155952
rect 210417 155894 294755 155896
rect 210417 155891 210483 155894
rect 294045 155891 294111 155894
rect 294689 155891 294755 155894
rect 177389 155410 177455 155413
rect 210509 155410 210575 155413
rect 177389 155408 210575 155410
rect 177389 155352 177394 155408
rect 177450 155352 210514 155408
rect 210570 155352 210575 155408
rect 177389 155350 210575 155352
rect 177389 155347 177455 155350
rect 210509 155347 210575 155350
rect 19333 155274 19399 155277
rect 188337 155274 188403 155277
rect 19333 155272 188403 155274
rect 19333 155216 19338 155272
rect 19394 155216 188342 155272
rect 188398 155216 188403 155272
rect 19333 155214 188403 155216
rect 19333 155211 19399 155214
rect 188337 155211 188403 155214
rect 240225 154458 240291 154461
rect 240777 154458 240843 154461
rect 240225 154456 240843 154458
rect 240225 154400 240230 154456
rect 240286 154400 240782 154456
rect 240838 154400 240843 154456
rect 240225 154398 240843 154400
rect 240225 154395 240291 154398
rect 240777 154395 240843 154398
rect 155401 153778 155467 153781
rect 187693 153778 187759 153781
rect 155401 153776 187759 153778
rect 155401 153720 155406 153776
rect 155462 153720 187698 153776
rect 187754 153720 187759 153776
rect 155401 153718 187759 153720
rect 155401 153715 155467 153718
rect 187693 153715 187759 153718
rect 190310 153716 190316 153780
rect 190380 153778 190386 153780
rect 193857 153778 193923 153781
rect 190380 153776 193923 153778
rect 190380 153720 193862 153776
rect 193918 153720 193923 153776
rect 190380 153718 193923 153720
rect 190380 153716 190386 153718
rect 193857 153715 193923 153718
rect 204989 153778 205055 153781
rect 211153 153778 211219 153781
rect 273529 153778 273595 153781
rect 204989 153776 273595 153778
rect 204989 153720 204994 153776
rect 205050 153720 211158 153776
rect 211214 153720 273534 153776
rect 273590 153720 273595 153776
rect 204989 153718 273595 153720
rect 204989 153715 205055 153718
rect 211153 153715 211219 153718
rect 273529 153715 273595 153718
rect 59077 153234 59143 153237
rect 124949 153234 125015 153237
rect 59077 153232 125015 153234
rect 59077 153176 59082 153232
rect 59138 153176 124954 153232
rect 125010 153176 125015 153232
rect 59077 153174 125015 153176
rect 59077 153171 59143 153174
rect 124949 153171 125015 153174
rect 134701 153234 134767 153237
rect 240225 153234 240291 153237
rect 134701 153232 240291 153234
rect 134701 153176 134706 153232
rect 134762 153176 240230 153232
rect 240286 153176 240291 153232
rect 134701 153174 240291 153176
rect 134701 153171 134767 153174
rect 240225 153171 240291 153174
rect 231945 153098 232011 153101
rect 232497 153098 232563 153101
rect 231945 153096 232563 153098
rect 231945 153040 231950 153096
rect 232006 153040 232502 153096
rect 232558 153040 232563 153096
rect 231945 153038 232563 153040
rect 231945 153035 232011 153038
rect 232497 153035 232563 153038
rect 582649 152690 582715 152693
rect 583520 152690 584960 152780
rect 582649 152688 584960 152690
rect 582649 152632 582654 152688
rect 582710 152632 584960 152688
rect 582649 152630 584960 152632
rect 582649 152627 582715 152630
rect 583520 152540 584960 152630
rect 81433 152418 81499 152421
rect 102133 152418 102199 152421
rect 81433 152416 102199 152418
rect 81433 152360 81438 152416
rect 81494 152360 102138 152416
rect 102194 152360 102199 152416
rect 81433 152358 102199 152360
rect 81433 152355 81499 152358
rect 102133 152355 102199 152358
rect 208485 152418 208551 152421
rect 281717 152418 281783 152421
rect 208485 152416 281783 152418
rect 208485 152360 208490 152416
rect 208546 152360 281722 152416
rect 281778 152360 281783 152416
rect 208485 152358 281783 152360
rect 208485 152355 208551 152358
rect 281717 152355 281783 152358
rect 204345 152010 204411 152013
rect 211797 152010 211863 152013
rect 204345 152008 211863 152010
rect 204345 151952 204350 152008
rect 204406 151952 211802 152008
rect 211858 151952 211863 152008
rect 204345 151950 211863 151952
rect 204345 151947 204411 151950
rect 211797 151947 211863 151950
rect 82813 151874 82879 151877
rect 86309 151874 86375 151877
rect 82813 151872 86375 151874
rect 82813 151816 82818 151872
rect 82874 151816 86314 151872
rect 86370 151816 86375 151872
rect 82813 151814 86375 151816
rect 82813 151811 82879 151814
rect 86309 151811 86375 151814
rect 102869 151874 102935 151877
rect 231945 151874 232011 151877
rect 102869 151872 232011 151874
rect 102869 151816 102874 151872
rect 102930 151816 231950 151872
rect 232006 151816 232011 151872
rect 102869 151814 232011 151816
rect 102869 151811 102935 151814
rect 231945 151811 232011 151814
rect 184473 151058 184539 151061
rect 211889 151058 211955 151061
rect 184473 151056 211955 151058
rect 184473 151000 184478 151056
rect 184534 151000 211894 151056
rect 211950 151000 211955 151056
rect 184473 150998 211955 151000
rect 184473 150995 184539 150998
rect 211889 150995 211955 150998
rect 169293 150650 169359 150653
rect 233233 150650 233299 150653
rect 169293 150648 233299 150650
rect 169293 150592 169298 150648
rect 169354 150592 233238 150648
rect 233294 150592 233299 150648
rect 169293 150590 233299 150592
rect 169293 150587 169359 150590
rect 233233 150587 233299 150590
rect 50889 150514 50955 150517
rect 184289 150514 184355 150517
rect 50889 150512 184355 150514
rect 50889 150456 50894 150512
rect 50950 150456 184294 150512
rect 184350 150456 184355 150512
rect 50889 150454 184355 150456
rect 50889 150451 50955 150454
rect 184289 150451 184355 150454
rect 220169 150514 220235 150517
rect 582925 150514 582991 150517
rect 220169 150512 582991 150514
rect 220169 150456 220174 150512
rect 220230 150456 582930 150512
rect 582986 150456 582991 150512
rect 220169 150454 582991 150456
rect 220169 150451 220235 150454
rect 582925 150451 582991 150454
rect -960 149834 480 149924
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 52269 149698 52335 149701
rect 189073 149698 189139 149701
rect 189625 149698 189691 149701
rect 52269 149696 189691 149698
rect 52269 149640 52274 149696
rect 52330 149640 189078 149696
rect 189134 149640 189630 149696
rect 189686 149640 189691 149696
rect 52269 149638 189691 149640
rect 52269 149635 52335 149638
rect 189073 149635 189139 149638
rect 189625 149635 189691 149638
rect 198825 149698 198891 149701
rect 207749 149698 207815 149701
rect 198825 149696 207815 149698
rect 198825 149640 198830 149696
rect 198886 149640 207754 149696
rect 207810 149640 207815 149696
rect 198825 149638 207815 149640
rect 198825 149635 198891 149638
rect 207749 149635 207815 149638
rect 66662 149092 66668 149156
rect 66732 149154 66738 149156
rect 67541 149154 67607 149157
rect 66732 149152 67607 149154
rect 66732 149096 67546 149152
rect 67602 149096 67607 149152
rect 66732 149094 67607 149096
rect 66732 149092 66738 149094
rect 67541 149091 67607 149094
rect 191741 149154 191807 149157
rect 240317 149154 240383 149157
rect 240777 149154 240843 149157
rect 191741 149152 240843 149154
rect 191741 149096 191746 149152
rect 191802 149096 240322 149152
rect 240378 149096 240782 149152
rect 240838 149096 240843 149152
rect 191741 149094 240843 149096
rect 191741 149091 191807 149094
rect 240317 149091 240383 149094
rect 240777 149091 240843 149094
rect 211061 148474 211127 148477
rect 224902 148474 224908 148476
rect 211061 148472 224908 148474
rect 211061 148416 211066 148472
rect 211122 148416 224908 148472
rect 211061 148414 224908 148416
rect 211061 148411 211127 148414
rect 224902 148412 224908 148414
rect 224972 148412 224978 148476
rect 87597 148338 87663 148341
rect 101581 148338 101647 148341
rect 87597 148336 101647 148338
rect 87597 148280 87602 148336
rect 87658 148280 101586 148336
rect 101642 148280 101647 148336
rect 87597 148278 101647 148280
rect 87597 148275 87663 148278
rect 101581 148275 101647 148278
rect 193806 148276 193812 148340
rect 193876 148338 193882 148340
rect 215293 148338 215359 148341
rect 193876 148336 215359 148338
rect 193876 148280 215298 148336
rect 215354 148280 215359 148336
rect 193876 148278 215359 148280
rect 193876 148276 193882 148278
rect 215293 148275 215359 148278
rect 173249 148066 173315 148069
rect 207013 148066 207079 148069
rect 173249 148064 207079 148066
rect 173249 148008 173254 148064
rect 173310 148008 207018 148064
rect 207074 148008 207079 148064
rect 173249 148006 207079 148008
rect 173249 148003 173315 148006
rect 207013 148003 207079 148006
rect 102777 147930 102843 147933
rect 193029 147930 193095 147933
rect 102777 147928 193095 147930
rect 102777 147872 102782 147928
rect 102838 147872 193034 147928
rect 193090 147872 193095 147928
rect 102777 147870 193095 147872
rect 102777 147867 102843 147870
rect 193029 147867 193095 147870
rect 188981 147794 189047 147797
rect 289813 147794 289879 147797
rect 188981 147792 289879 147794
rect 188981 147736 188986 147792
rect 189042 147736 289818 147792
rect 289874 147736 289879 147792
rect 188981 147734 289879 147736
rect 188981 147731 189047 147734
rect 289813 147731 289879 147734
rect 192937 146978 193003 146981
rect 245101 146978 245167 146981
rect 192937 146976 245167 146978
rect 192937 146920 192942 146976
rect 192998 146920 245106 146976
rect 245162 146920 245167 146976
rect 192937 146918 245167 146920
rect 192937 146915 193003 146918
rect 245101 146915 245167 146918
rect 181529 146570 181595 146573
rect 226609 146570 226675 146573
rect 181529 146568 226675 146570
rect 181529 146512 181534 146568
rect 181590 146512 226614 146568
rect 226670 146512 226675 146568
rect 181529 146510 226675 146512
rect 181529 146507 181595 146510
rect 226609 146507 226675 146510
rect 70393 146434 70459 146437
rect 71630 146434 71636 146436
rect 70393 146432 71636 146434
rect 70393 146376 70398 146432
rect 70454 146376 71636 146432
rect 70393 146374 71636 146376
rect 70393 146371 70459 146374
rect 71630 146372 71636 146374
rect 71700 146434 71706 146436
rect 196525 146434 196591 146437
rect 71700 146432 196591 146434
rect 71700 146376 196530 146432
rect 196586 146376 196591 146432
rect 71700 146374 196591 146376
rect 71700 146372 71706 146374
rect 196525 146371 196591 146374
rect 187693 145890 187759 145893
rect 191649 145890 191715 145893
rect 187693 145888 191715 145890
rect 187693 145832 187698 145888
rect 187754 145832 191654 145888
rect 191710 145832 191715 145888
rect 187693 145830 191715 145832
rect 187693 145827 187759 145830
rect 191649 145827 191715 145830
rect 177481 145754 177547 145757
rect 204897 145754 204963 145757
rect 177481 145752 204963 145754
rect 177481 145696 177486 145752
rect 177542 145696 204902 145752
rect 204958 145696 204963 145752
rect 177481 145694 204963 145696
rect 177481 145691 177547 145694
rect 204897 145691 204963 145694
rect 93945 145618 94011 145621
rect 169109 145618 169175 145621
rect 93945 145616 169175 145618
rect 93945 145560 93950 145616
rect 94006 145560 169114 145616
rect 169170 145560 169175 145616
rect 93945 145558 169175 145560
rect 93945 145555 94011 145558
rect 169109 145555 169175 145558
rect 191649 145618 191715 145621
rect 252185 145618 252251 145621
rect 191649 145616 252251 145618
rect 191649 145560 191654 145616
rect 191710 145560 252190 145616
rect 252246 145560 252251 145616
rect 191649 145558 252251 145560
rect 191649 145555 191715 145558
rect 252185 145555 252251 145558
rect 72877 145076 72943 145077
rect 72877 145074 72924 145076
rect 72832 145072 72924 145074
rect 72832 145016 72882 145072
rect 72832 145014 72924 145016
rect 72877 145012 72924 145014
rect 72988 145012 72994 145076
rect 86309 145074 86375 145077
rect 159541 145074 159607 145077
rect 86309 145072 159607 145074
rect 86309 145016 86314 145072
rect 86370 145016 159546 145072
rect 159602 145016 159607 145072
rect 86309 145014 159607 145016
rect 72877 145011 72943 145012
rect 86309 145011 86375 145014
rect 159541 145011 159607 145014
rect 153929 144938 153995 144941
rect 227989 144938 228055 144941
rect 153929 144936 228055 144938
rect 153929 144880 153934 144936
rect 153990 144880 227994 144936
rect 228050 144880 228055 144936
rect 153929 144878 228055 144880
rect 153929 144875 153995 144878
rect 227989 144875 228055 144878
rect 86861 144802 86927 144805
rect 89846 144802 89852 144804
rect 86861 144800 89852 144802
rect 86861 144744 86866 144800
rect 86922 144744 89852 144800
rect 86861 144742 89852 144744
rect 86861 144739 86927 144742
rect 89846 144740 89852 144742
rect 89916 144740 89922 144804
rect 97533 144802 97599 144805
rect 99966 144802 99972 144804
rect 97533 144800 99972 144802
rect 97533 144744 97538 144800
rect 97594 144744 99972 144800
rect 97533 144742 99972 144744
rect 97533 144739 97599 144742
rect 99966 144740 99972 144742
rect 100036 144740 100042 144804
rect 182173 144802 182239 144805
rect 183461 144802 183527 144805
rect 197905 144804 197971 144805
rect 197854 144802 197860 144804
rect 182173 144800 183527 144802
rect 182173 144744 182178 144800
rect 182234 144744 183466 144800
rect 183522 144744 183527 144800
rect 182173 144742 183527 144744
rect 197814 144742 197860 144802
rect 197924 144800 197971 144804
rect 197966 144744 197971 144800
rect 182173 144739 182239 144742
rect 183461 144739 183527 144742
rect 197854 144740 197860 144742
rect 197924 144740 197971 144744
rect 197905 144739 197971 144740
rect 222837 144802 222903 144805
rect 223614 144802 223620 144804
rect 222837 144800 223620 144802
rect 222837 144744 222842 144800
rect 222898 144744 223620 144800
rect 222837 144742 223620 144744
rect 222837 144739 222903 144742
rect 223614 144740 223620 144742
rect 223684 144740 223690 144804
rect 191097 144258 191163 144261
rect 224493 144258 224559 144261
rect 191097 144256 224559 144258
rect 191097 144200 191102 144256
rect 191158 144200 224498 144256
rect 224554 144200 224559 144256
rect 191097 144198 224559 144200
rect 191097 144195 191163 144198
rect 224493 144195 224559 144198
rect 185761 144122 185827 144125
rect 201309 144122 201375 144125
rect 185761 144120 201375 144122
rect 185761 144064 185766 144120
rect 185822 144064 201314 144120
rect 201370 144064 201375 144120
rect 185761 144062 201375 144064
rect 185761 144059 185827 144062
rect 201309 144059 201375 144062
rect 210509 144122 210575 144125
rect 285949 144122 286015 144125
rect 210509 144120 286015 144122
rect 210509 144064 210514 144120
rect 210570 144064 285954 144120
rect 286010 144064 286015 144120
rect 210509 144062 286015 144064
rect 210509 144059 210575 144062
rect 285949 144059 286015 144062
rect 183461 143714 183527 143717
rect 215845 143714 215911 143717
rect 183461 143712 215911 143714
rect 183461 143656 183466 143712
rect 183522 143656 215850 143712
rect 215906 143656 215911 143712
rect 183461 143654 215911 143656
rect 183461 143651 183527 143654
rect 215845 143651 215911 143654
rect 54937 143578 55003 143581
rect 185577 143578 185643 143581
rect 54937 143576 185643 143578
rect 54937 143520 54942 143576
rect 54998 143520 185582 143576
rect 185638 143520 185643 143576
rect 54937 143518 185643 143520
rect 54937 143515 55003 143518
rect 185577 143515 185643 143518
rect 83457 142626 83523 142629
rect 83457 142624 195990 142626
rect 83457 142568 83462 142624
rect 83518 142568 195990 142624
rect 83457 142566 195990 142568
rect 83457 142563 83523 142566
rect 76005 142490 76071 142493
rect 194593 142490 194659 142493
rect 76005 142488 194659 142490
rect 76005 142432 76010 142488
rect 76066 142432 194598 142488
rect 194654 142432 194659 142488
rect 76005 142430 194659 142432
rect 195930 142490 195990 142566
rect 212349 142490 212415 142493
rect 224350 142490 224356 142492
rect 195930 142488 224356 142490
rect 195930 142432 212354 142488
rect 212410 142432 224356 142488
rect 195930 142430 224356 142432
rect 76005 142427 76071 142430
rect 194593 142427 194659 142430
rect 212349 142427 212415 142430
rect 224350 142428 224356 142430
rect 224420 142428 224426 142492
rect 73797 142354 73863 142357
rect 196566 142354 196572 142356
rect 73797 142352 196572 142354
rect 73797 142296 73802 142352
rect 73858 142296 196572 142352
rect 73797 142294 196572 142296
rect 73797 142291 73863 142294
rect 196566 142292 196572 142294
rect 196636 142354 196642 142356
rect 196709 142354 196775 142357
rect 196636 142352 196775 142354
rect 196636 142296 196714 142352
rect 196770 142296 196775 142352
rect 196636 142294 196775 142296
rect 196636 142292 196642 142294
rect 196709 142291 196775 142294
rect 224217 142354 224283 142357
rect 232497 142354 232563 142357
rect 224217 142352 232563 142354
rect 224217 142296 224222 142352
rect 224278 142296 232502 142352
rect 232558 142296 232563 142352
rect 224217 142294 232563 142296
rect 224217 142291 224283 142294
rect 232497 142291 232563 142294
rect 202873 142218 202939 142221
rect 203190 142218 203196 142220
rect 202873 142216 203196 142218
rect 202873 142160 202878 142216
rect 202934 142160 203196 142216
rect 202873 142158 203196 142160
rect 202873 142155 202939 142158
rect 203190 142156 203196 142158
rect 203260 142218 203266 142220
rect 203885 142218 203951 142221
rect 203260 142216 203951 142218
rect 203260 142160 203890 142216
rect 203946 142160 203951 142216
rect 203260 142158 203951 142160
rect 203260 142156 203266 142158
rect 203885 142155 203951 142158
rect 218237 142218 218303 142221
rect 323577 142218 323643 142221
rect 218237 142216 323643 142218
rect 218237 142160 218242 142216
rect 218298 142160 323582 142216
rect 323638 142160 323643 142216
rect 218237 142158 323643 142160
rect 218237 142155 218303 142158
rect 323577 142155 323643 142158
rect 79961 141538 80027 141541
rect 173249 141538 173315 141541
rect 79961 141536 173315 141538
rect 79961 141480 79966 141536
rect 80022 141480 173254 141536
rect 173310 141480 173315 141536
rect 79961 141478 173315 141480
rect 79961 141475 80027 141478
rect 173249 141475 173315 141478
rect 207657 141538 207723 141541
rect 222837 141538 222903 141541
rect 207657 141536 222903 141538
rect 207657 141480 207662 141536
rect 207718 141480 222842 141536
rect 222898 141480 222903 141536
rect 207657 141478 222903 141480
rect 207657 141475 207723 141478
rect 222837 141475 222903 141478
rect 53557 141402 53623 141405
rect 71405 141402 71471 141405
rect 53557 141400 71471 141402
rect 53557 141344 53562 141400
rect 53618 141344 71410 141400
rect 71466 141344 71471 141400
rect 53557 141342 71471 141344
rect 53557 141339 53623 141342
rect 71405 141339 71471 141342
rect 80605 141402 80671 141405
rect 83406 141402 83412 141404
rect 80605 141400 83412 141402
rect 80605 141344 80610 141400
rect 80666 141344 83412 141400
rect 80605 141342 83412 141344
rect 80605 141339 80671 141342
rect 83406 141340 83412 141342
rect 83476 141402 83482 141404
rect 207841 141402 207907 141405
rect 208117 141402 208183 141405
rect 83476 141400 208183 141402
rect 83476 141344 207846 141400
rect 207902 141344 208122 141400
rect 208178 141344 208183 141400
rect 83476 141342 208183 141344
rect 83476 141340 83482 141342
rect 207841 141339 207907 141342
rect 208117 141339 208183 141342
rect 193070 141068 193076 141132
rect 193140 141130 193146 141132
rect 195237 141130 195303 141133
rect 193140 141128 195303 141130
rect 193140 141072 195242 141128
rect 195298 141072 195303 141128
rect 193140 141070 195303 141072
rect 193140 141068 193146 141070
rect 195237 141067 195303 141070
rect 222193 141130 222259 141133
rect 223205 141130 223271 141133
rect 222193 141128 223271 141130
rect 222193 141072 222198 141128
rect 222254 141072 223210 141128
rect 223266 141072 223271 141128
rect 222193 141070 223271 141072
rect 222193 141067 222259 141070
rect 223205 141067 223271 141070
rect 193213 140858 193279 140861
rect 206553 140858 206619 140861
rect 193213 140856 206619 140858
rect 193213 140800 193218 140856
rect 193274 140800 206558 140856
rect 206614 140800 206619 140856
rect 193213 140798 206619 140800
rect 193213 140795 193279 140798
rect 206553 140795 206619 140798
rect 223389 140858 223455 140861
rect 238017 140858 238083 140861
rect 223389 140856 238083 140858
rect 223389 140800 223394 140856
rect 223450 140800 238022 140856
rect 238078 140800 238083 140856
rect 223389 140798 238083 140800
rect 223389 140795 223455 140798
rect 238017 140795 238083 140798
rect 222837 140722 222903 140725
rect 226374 140722 226380 140724
rect 222837 140720 226380 140722
rect 222837 140664 222842 140720
rect 222898 140664 226380 140720
rect 222837 140662 226380 140664
rect 222837 140659 222903 140662
rect 226374 140660 226380 140662
rect 226444 140660 226450 140724
rect 209037 140586 209103 140589
rect 209814 140586 209820 140588
rect 209037 140584 209820 140586
rect 209037 140528 209042 140584
rect 209098 140528 209820 140584
rect 209037 140526 209820 140528
rect 209037 140523 209103 140526
rect 209814 140524 209820 140526
rect 209884 140524 209890 140588
rect 210141 140586 210207 140589
rect 215385 140586 215451 140589
rect 210141 140584 215451 140586
rect 210141 140528 210146 140584
rect 210202 140528 215390 140584
rect 215446 140528 215451 140584
rect 210141 140526 215451 140528
rect 210141 140523 210207 140526
rect 215385 140523 215451 140526
rect 194961 140450 195027 140453
rect 195094 140450 195100 140452
rect 194961 140448 195100 140450
rect 194961 140392 194966 140448
rect 195022 140392 195100 140448
rect 194961 140390 195100 140392
rect 194961 140387 195027 140390
rect 195094 140388 195100 140390
rect 195164 140388 195170 140452
rect 86861 140178 86927 140181
rect 193397 140178 193463 140181
rect 86861 140176 193463 140178
rect 86861 140120 86866 140176
rect 86922 140120 193402 140176
rect 193458 140120 193463 140176
rect 86861 140118 193463 140120
rect 86861 140115 86927 140118
rect 193397 140115 193463 140118
rect 65926 139980 65932 140044
rect 65996 140042 66002 140044
rect 86309 140042 86375 140045
rect 65996 140040 86375 140042
rect 65996 139984 86314 140040
rect 86370 139984 86375 140040
rect 65996 139982 86375 139984
rect 65996 139980 66002 139982
rect 86309 139979 86375 139982
rect 192845 139906 192911 139909
rect 228357 139906 228423 139909
rect 192845 139904 193660 139906
rect 192845 139848 192850 139904
rect 192906 139848 193660 139904
rect 192845 139846 193660 139848
rect 224940 139904 228423 139906
rect 224940 139848 228362 139904
rect 228418 139848 228423 139904
rect 224940 139846 228423 139848
rect 192845 139843 192911 139846
rect 228357 139843 228423 139846
rect 68686 139572 68692 139636
rect 68756 139634 68762 139636
rect 70485 139634 70551 139637
rect 68756 139632 70551 139634
rect 68756 139576 70490 139632
rect 70546 139576 70551 139632
rect 68756 139574 70551 139576
rect 68756 139572 68762 139574
rect 70485 139571 70551 139574
rect 53465 139498 53531 139501
rect 53741 139498 53807 139501
rect 95969 139498 96035 139501
rect 53465 139496 96035 139498
rect 53465 139440 53470 139496
rect 53526 139440 53746 139496
rect 53802 139440 95974 139496
rect 96030 139440 96035 139496
rect 53465 139438 96035 139440
rect 53465 139435 53531 139438
rect 53741 139435 53807 139438
rect 95969 139435 96035 139438
rect 583017 139362 583083 139365
rect 583520 139362 584960 139452
rect 583017 139360 584960 139362
rect 583017 139304 583022 139360
rect 583078 139304 584960 139360
rect 583017 139302 584960 139304
rect 583017 139299 583083 139302
rect 583520 139212 584960 139302
rect 193070 139028 193076 139092
rect 193140 139090 193146 139092
rect 226701 139090 226767 139093
rect 193140 139030 193660 139090
rect 224940 139088 226767 139090
rect 224940 139032 226706 139088
rect 226762 139032 226767 139088
rect 224940 139030 226767 139032
rect 193140 139028 193146 139030
rect 226701 139027 226767 139030
rect 235993 138954 236059 138957
rect 224910 138952 236059 138954
rect 224910 138896 235998 138952
rect 236054 138896 236059 138952
rect 224910 138894 236059 138896
rect 78029 138682 78095 138685
rect 115289 138682 115355 138685
rect 78029 138680 115355 138682
rect 78029 138624 78034 138680
rect 78090 138624 115294 138680
rect 115350 138624 115355 138680
rect 78029 138622 115355 138624
rect 78029 138619 78095 138622
rect 115289 138619 115355 138622
rect 72918 138348 72924 138412
rect 72988 138410 72994 138412
rect 73153 138410 73219 138413
rect 72988 138408 73219 138410
rect 72988 138352 73158 138408
rect 73214 138352 73219 138408
rect 72988 138350 73219 138352
rect 72988 138348 72994 138350
rect 73153 138347 73219 138350
rect 64505 138274 64571 138277
rect 93761 138274 93827 138277
rect 64505 138272 93827 138274
rect 64505 138216 64510 138272
rect 64566 138216 93766 138272
rect 93822 138216 93827 138272
rect 64505 138214 93827 138216
rect 64505 138211 64571 138214
rect 93761 138211 93827 138214
rect 193029 138274 193095 138277
rect 193029 138272 193660 138274
rect 193029 138216 193034 138272
rect 193090 138216 193660 138272
rect 224910 138244 224970 138894
rect 235993 138891 236059 138894
rect 193029 138214 193660 138216
rect 193029 138211 193095 138214
rect 55029 138138 55095 138141
rect 94681 138138 94747 138141
rect 55029 138136 94747 138138
rect 55029 138080 55034 138136
rect 55090 138080 94686 138136
rect 94742 138080 94747 138136
rect 55029 138078 94747 138080
rect 55029 138075 55095 138078
rect 94681 138075 94747 138078
rect 70209 138002 70275 138005
rect 71814 138002 71820 138004
rect 70209 138000 71820 138002
rect 70209 137944 70214 138000
rect 70270 137944 71820 138000
rect 70209 137942 71820 137944
rect 70209 137939 70275 137942
rect 71814 137940 71820 137942
rect 71884 137940 71890 138004
rect 88517 138002 88583 138005
rect 155953 138002 156019 138005
rect 156413 138002 156479 138005
rect 88517 138000 156479 138002
rect 88517 137944 88522 138000
rect 88578 137944 155958 138000
rect 156014 137944 156418 138000
rect 156474 137944 156479 138000
rect 88517 137942 156479 137944
rect 88517 137939 88583 137942
rect 155953 137939 156019 137942
rect 156413 137939 156479 137942
rect 152641 137866 152707 137869
rect 191097 137866 191163 137869
rect 152641 137864 191163 137866
rect 152641 137808 152646 137864
rect 152702 137808 191102 137864
rect 191158 137808 191163 137864
rect 152641 137806 191163 137808
rect 152641 137803 152707 137806
rect 191097 137803 191163 137806
rect 87045 137596 87111 137597
rect 87045 137592 87092 137596
rect 87156 137594 87162 137596
rect 87045 137536 87050 137592
rect 87045 137532 87092 137536
rect 87156 137534 87202 137594
rect 87156 137532 87162 137534
rect 87045 137531 87111 137532
rect 70158 137396 70164 137460
rect 70228 137458 70234 137460
rect 72325 137458 72391 137461
rect 79317 137458 79383 137461
rect 70228 137456 72391 137458
rect 70228 137400 72330 137456
rect 72386 137400 72391 137456
rect 70228 137398 72391 137400
rect 70228 137396 70234 137398
rect 72325 137395 72391 137398
rect 72558 137456 79383 137458
rect 72558 137400 79322 137456
rect 79378 137400 79383 137456
rect 72558 137398 79383 137400
rect 70158 137260 70164 137324
rect 70228 137322 70234 137324
rect 72558 137322 72618 137398
rect 79317 137395 79383 137398
rect 70228 137262 72618 137322
rect 74257 137322 74323 137325
rect 87689 137322 87755 137325
rect 74257 137320 87755 137322
rect 74257 137264 74262 137320
rect 74318 137264 87694 137320
rect 87750 137264 87755 137320
rect 74257 137262 87755 137264
rect 70228 137260 70234 137262
rect 74257 137259 74323 137262
rect 87689 137259 87755 137262
rect 156413 137322 156479 137325
rect 169201 137322 169267 137325
rect 156413 137320 169267 137322
rect 156413 137264 156418 137320
rect 156474 137264 169206 137320
rect 169262 137264 169267 137320
rect 156413 137262 169267 137264
rect 156413 137259 156479 137262
rect 169201 137259 169267 137262
rect 79041 136914 79107 136917
rect 82077 136914 82143 136917
rect 79041 136912 82143 136914
rect -960 136778 480 136868
rect 79041 136856 79046 136912
rect 79102 136856 82082 136912
rect 82138 136856 82143 136912
rect 79041 136854 82143 136856
rect 79041 136851 79107 136854
rect 82077 136851 82143 136854
rect 2865 136778 2931 136781
rect -960 136776 2931 136778
rect -960 136720 2870 136776
rect 2926 136720 2931 136776
rect -960 136718 2931 136720
rect -960 136628 480 136718
rect 2865 136715 2931 136718
rect 81893 136778 81959 136781
rect 95141 136778 95207 136781
rect 81893 136776 95207 136778
rect 81893 136720 81898 136776
rect 81954 136720 95146 136776
rect 95202 136720 95207 136776
rect 81893 136718 95207 136720
rect 81893 136715 81959 136718
rect 95141 136715 95207 136718
rect 189809 136778 189875 136781
rect 193630 136778 193690 137428
rect 226701 137186 226767 137189
rect 224940 137184 226767 137186
rect 224940 137128 226706 137184
rect 226762 137128 226767 137184
rect 224940 137126 226767 137128
rect 226701 137123 226767 137126
rect 189809 136776 193690 136778
rect 189809 136720 189814 136776
rect 189870 136720 193690 136776
rect 189809 136718 193690 136720
rect 189809 136715 189875 136718
rect 69422 136580 69428 136644
rect 69492 136642 69498 136644
rect 76649 136642 76715 136645
rect 226609 136642 226675 136645
rect 259494 136642 259500 136644
rect 69492 136640 76715 136642
rect 69492 136584 76654 136640
rect 76710 136584 76715 136640
rect 69492 136582 76715 136584
rect 69492 136580 69498 136582
rect 76649 136579 76715 136582
rect 224910 136640 259500 136642
rect 224910 136584 226614 136640
rect 226670 136584 259500 136640
rect 224910 136582 259500 136584
rect 191557 136370 191623 136373
rect 191557 136368 193660 136370
rect 191557 136312 191562 136368
rect 191618 136312 193660 136368
rect 224910 136340 224970 136582
rect 226609 136579 226675 136582
rect 259494 136580 259500 136582
rect 259564 136580 259570 136644
rect 191557 136310 193660 136312
rect 191557 136307 191623 136310
rect 81065 136234 81131 136237
rect 151261 136234 151327 136237
rect 81065 136232 151327 136234
rect 81065 136176 81070 136232
rect 81126 136176 151266 136232
rect 151322 136176 151327 136232
rect 81065 136174 151327 136176
rect 81065 136171 81131 136174
rect 151261 136171 151327 136174
rect 67817 136098 67883 136101
rect 160185 136098 160251 136101
rect 67817 136096 160251 136098
rect 67817 136040 67822 136096
rect 67878 136040 160190 136096
rect 160246 136040 160251 136096
rect 67817 136038 160251 136040
rect 67817 136035 67883 136038
rect 160185 136035 160251 136038
rect 87045 135962 87111 135965
rect 182173 135962 182239 135965
rect 87045 135960 182239 135962
rect 87045 135904 87050 135960
rect 87106 135904 182178 135960
rect 182234 135904 182239 135960
rect 87045 135902 182239 135904
rect 87045 135899 87111 135902
rect 182173 135899 182239 135902
rect 191557 135554 191623 135557
rect 226701 135554 226767 135557
rect 191557 135552 193660 135554
rect 191557 135496 191562 135552
rect 191618 135496 193660 135552
rect 191557 135494 193660 135496
rect 224940 135552 226767 135554
rect 224940 135496 226706 135552
rect 226762 135496 226767 135552
rect 224940 135494 226767 135496
rect 191557 135491 191623 135494
rect 226701 135491 226767 135494
rect 72366 135084 72372 135148
rect 72436 135146 72442 135148
rect 73061 135146 73127 135149
rect 72436 135144 73127 135146
rect 72436 135088 73066 135144
rect 73122 135088 73127 135144
rect 72436 135086 73127 135088
rect 72436 135084 72442 135086
rect 73061 135083 73127 135086
rect 3417 134874 3483 134877
rect 70301 134874 70367 134877
rect 3417 134872 70367 134874
rect 3417 134816 3422 134872
rect 3478 134816 70306 134872
rect 70362 134816 70367 134872
rect 3417 134814 70367 134816
rect 3417 134811 3483 134814
rect 70301 134811 70367 134814
rect 69657 134738 69723 134741
rect 69430 134736 69723 134738
rect 69430 134680 69662 134736
rect 69718 134680 69723 134736
rect 69430 134678 69723 134680
rect 69430 134436 69490 134678
rect 69657 134675 69723 134678
rect 190453 134738 190519 134741
rect 226425 134738 226491 134741
rect 226609 134738 226675 134741
rect 190453 134736 193660 134738
rect 190453 134680 190458 134736
rect 190514 134680 193660 134736
rect 190453 134678 193660 134680
rect 224940 134736 226675 134738
rect 224940 134680 226430 134736
rect 226486 134680 226614 134736
rect 226670 134680 226675 134736
rect 224940 134678 226675 134680
rect 190453 134675 190519 134678
rect 226425 134675 226491 134678
rect 226609 134675 226675 134678
rect 189165 134602 189231 134605
rect 190310 134602 190316 134604
rect 189165 134600 190316 134602
rect 189165 134544 189170 134600
rect 189226 134544 190316 134600
rect 189165 134542 190316 134544
rect 189165 134539 189231 134542
rect 190310 134540 190316 134542
rect 190380 134540 190386 134604
rect 97901 133922 97967 133925
rect 94668 133920 97967 133922
rect 94668 133864 97906 133920
rect 97962 133864 97967 133920
rect 94668 133862 97967 133864
rect 97901 133859 97967 133862
rect 191189 133922 191255 133925
rect 191189 133920 193660 133922
rect 191189 133864 191194 133920
rect 191250 133864 193660 133920
rect 191189 133862 193660 133864
rect 191189 133859 191255 133862
rect 65977 133650 66043 133653
rect 226701 133650 226767 133653
rect 65977 133648 68908 133650
rect 65977 133592 65982 133648
rect 66038 133592 68908 133648
rect 65977 133590 68908 133592
rect 224940 133648 226767 133650
rect 224940 133592 226706 133648
rect 226762 133592 226767 133648
rect 224940 133590 226767 133592
rect 65977 133587 66043 133590
rect 226701 133587 226767 133590
rect 224350 133452 224356 133516
rect 224420 133514 224426 133516
rect 284937 133514 285003 133517
rect 224420 133512 287070 133514
rect 224420 133456 284942 133512
rect 284998 133456 287070 133512
rect 224420 133454 287070 133456
rect 224420 133452 224426 133454
rect 284937 133451 285003 133454
rect 69422 133316 69428 133380
rect 69492 133316 69498 133380
rect 69430 132804 69490 133316
rect 164141 133106 164207 133109
rect 182817 133106 182883 133109
rect 164141 133104 182883 133106
rect 94638 132562 94698 133076
rect 164141 133048 164146 133104
rect 164202 133048 182822 133104
rect 182878 133048 182883 133104
rect 164141 133046 182883 133048
rect 287010 133106 287070 133454
rect 317413 133106 317479 133109
rect 287010 133104 317479 133106
rect 287010 133048 317418 133104
rect 317474 133048 317479 133104
rect 287010 133046 317479 133048
rect 164141 133043 164207 133046
rect 182817 133043 182883 133046
rect 317413 133043 317479 133046
rect 226609 132834 226675 132837
rect 224940 132832 226675 132834
rect 105537 132562 105603 132565
rect 94638 132560 105603 132562
rect 94638 132504 105542 132560
rect 105598 132504 105603 132560
rect 94638 132502 105603 132504
rect 105537 132499 105603 132502
rect 190310 132500 190316 132564
rect 190380 132562 190386 132564
rect 193630 132562 193690 132804
rect 224940 132776 226614 132832
rect 226670 132776 226675 132832
rect 224940 132774 226675 132776
rect 226609 132771 226675 132774
rect 190380 132502 193690 132562
rect 190380 132500 190386 132502
rect 97901 132290 97967 132293
rect 94668 132288 97967 132290
rect 94668 132232 97906 132288
rect 97962 132232 97967 132288
rect 94668 132230 97967 132232
rect 97901 132227 97967 132230
rect 66897 132018 66963 132021
rect 66897 132016 68908 132018
rect 66897 131960 66902 132016
rect 66958 131960 68908 132016
rect 66897 131958 68908 131960
rect 66897 131955 66963 131958
rect 192702 131956 192708 132020
rect 192772 132018 192778 132020
rect 226701 132018 226767 132021
rect 192772 131958 193660 132018
rect 224940 132016 226767 132018
rect 224940 131960 226706 132016
rect 226762 131960 226767 132016
rect 224940 131958 226767 131960
rect 192772 131956 192778 131958
rect 226701 131955 226767 131958
rect 94681 131882 94747 131885
rect 193213 131882 193279 131885
rect 94681 131880 193279 131882
rect 94681 131824 94686 131880
rect 94742 131824 193218 131880
rect 193274 131824 193279 131880
rect 94681 131822 193279 131824
rect 94681 131819 94747 131822
rect 193213 131819 193279 131822
rect 97533 131474 97599 131477
rect 94668 131472 97599 131474
rect 94668 131416 97538 131472
rect 97594 131416 97599 131472
rect 94668 131414 97599 131416
rect 97533 131411 97599 131414
rect 188889 131474 188955 131477
rect 192702 131474 192708 131476
rect 188889 131472 192708 131474
rect 188889 131416 188894 131472
rect 188950 131416 192708 131472
rect 188889 131414 192708 131416
rect 188889 131411 188955 131414
rect 192702 131412 192708 131414
rect 192772 131412 192778 131476
rect 193213 131474 193279 131477
rect 193438 131474 193444 131476
rect 193213 131472 193444 131474
rect 193213 131416 193218 131472
rect 193274 131416 193444 131472
rect 193213 131414 193444 131416
rect 193213 131411 193279 131414
rect 193438 131412 193444 131414
rect 193508 131412 193514 131476
rect 66805 131202 66871 131205
rect 66805 131200 68908 131202
rect 66805 131144 66810 131200
rect 66866 131144 68908 131200
rect 66805 131142 68908 131144
rect 66805 131139 66871 131142
rect 188286 131140 188292 131204
rect 188356 131202 188362 131204
rect 188356 131142 193660 131202
rect 188356 131140 188362 131142
rect 96613 130930 96679 130933
rect 97717 130930 97783 130933
rect 226701 130930 226767 130933
rect 94668 130928 97783 130930
rect 94668 130872 96618 130928
rect 96674 130872 97722 130928
rect 97778 130872 97783 130928
rect 94668 130870 97783 130872
rect 224940 130928 226767 130930
rect 224940 130872 226706 130928
rect 226762 130872 226767 130928
rect 224940 130870 226767 130872
rect 96613 130867 96679 130870
rect 97717 130867 97783 130870
rect 226701 130867 226767 130870
rect 66805 130658 66871 130661
rect 66805 130656 68908 130658
rect 66805 130600 66810 130656
rect 66866 130600 68908 130656
rect 66805 130598 68908 130600
rect 66805 130595 66871 130598
rect 97533 130114 97599 130117
rect 226793 130114 226859 130117
rect 94668 130112 97599 130114
rect 94668 130056 97538 130112
rect 97594 130056 97599 130112
rect 224940 130112 226859 130114
rect 94668 130054 97599 130056
rect 97533 130051 97599 130054
rect 66713 129842 66779 129845
rect 190361 129842 190427 129845
rect 193630 129842 193690 130084
rect 224940 130056 226798 130112
rect 226854 130056 226859 130112
rect 224940 130054 226859 130056
rect 226793 130051 226859 130054
rect 66713 129840 68908 129842
rect 66713 129784 66718 129840
rect 66774 129784 68908 129840
rect 66713 129782 68908 129784
rect 190361 129840 193690 129842
rect 190361 129784 190366 129840
rect 190422 129784 193690 129840
rect 190361 129782 193690 129784
rect 66713 129779 66779 129782
rect 190361 129779 190427 129782
rect 225045 129706 225111 129709
rect 224910 129704 225111 129706
rect 224910 129648 225050 129704
rect 225106 129648 225111 129704
rect 224910 129646 225111 129648
rect 100702 129298 100708 129300
rect 94668 129238 100708 129298
rect 100702 129236 100708 129238
rect 100772 129236 100778 129300
rect 191741 129298 191807 129301
rect 224910 129298 224970 129646
rect 225045 129643 225111 129646
rect 227897 129298 227963 129301
rect 191741 129296 193660 129298
rect 191741 129240 191746 129296
rect 191802 129240 193660 129296
rect 224910 129296 227963 129298
rect 224910 129268 227902 129296
rect 191741 129238 193660 129240
rect 224940 129240 227902 129268
rect 227958 129240 227963 129296
rect 224940 129238 227963 129240
rect 191741 129235 191807 129238
rect 227897 129235 227963 129238
rect 66805 129026 66871 129029
rect 105537 129026 105603 129029
rect 128997 129026 129063 129029
rect 66805 129024 68908 129026
rect 66805 128968 66810 129024
rect 66866 128968 68908 129024
rect 66805 128966 68908 128968
rect 105537 129024 129063 129026
rect 105537 128968 105542 129024
rect 105598 128968 129002 129024
rect 129058 128968 129063 129024
rect 105537 128966 129063 128968
rect 66805 128963 66871 128966
rect 105537 128963 105603 128966
rect 128997 128963 129063 128966
rect 224350 128964 224356 129028
rect 224420 129026 224426 129028
rect 226609 129026 226675 129029
rect 259453 129026 259519 129029
rect 224420 128966 224970 129026
rect 224420 128964 224426 128966
rect 97901 128482 97967 128485
rect 94668 128480 97967 128482
rect 94668 128424 97906 128480
rect 97962 128424 97967 128480
rect 94668 128422 97967 128424
rect 97901 128419 97967 128422
rect 191649 128482 191715 128485
rect 224910 128482 224970 128966
rect 226609 129024 259519 129026
rect 226609 128968 226614 129024
rect 226670 128968 259458 129024
rect 259514 128968 259519 129024
rect 226609 128966 259519 128968
rect 226609 128963 226675 128966
rect 259453 128963 259519 128966
rect 226425 128482 226491 128485
rect 191649 128480 193660 128482
rect 191649 128424 191654 128480
rect 191710 128424 193660 128480
rect 224910 128480 226491 128482
rect 224910 128452 226430 128480
rect 191649 128422 193660 128424
rect 224940 128424 226430 128452
rect 226486 128424 226491 128480
rect 224940 128422 226491 128424
rect 191649 128419 191715 128422
rect 226425 128419 226491 128422
rect 68553 128210 68619 128213
rect 68553 128208 68908 128210
rect 68553 128152 68558 128208
rect 68614 128152 68908 128208
rect 68553 128150 68908 128152
rect 68553 128147 68619 128150
rect 67725 127666 67791 127669
rect 95417 127666 95483 127669
rect 67725 127664 68908 127666
rect 67725 127608 67730 127664
rect 67786 127608 68908 127664
rect 67725 127606 68908 127608
rect 94668 127664 95483 127666
rect 94668 127608 95422 127664
rect 95478 127608 95483 127664
rect 94668 127606 95483 127608
rect 67725 127603 67791 127606
rect 95417 127603 95483 127606
rect 191741 127666 191807 127669
rect 191741 127664 193660 127666
rect 191741 127608 191746 127664
rect 191802 127608 193660 127664
rect 191741 127606 193660 127608
rect 191741 127603 191807 127606
rect 226701 127394 226767 127397
rect 224940 127392 226767 127394
rect 224940 127336 226706 127392
rect 226762 127336 226767 127392
rect 224940 127334 226767 127336
rect 226701 127331 226767 127334
rect 97625 127122 97691 127125
rect 94668 127120 97691 127122
rect 94668 127064 97630 127120
rect 97686 127064 97691 127120
rect 94668 127062 97691 127064
rect 97625 127059 97691 127062
rect 227897 126986 227963 126989
rect 281625 126986 281691 126989
rect 227897 126984 281691 126986
rect 227897 126928 227902 126984
rect 227958 126928 281630 126984
rect 281686 126928 281691 126984
rect 227897 126926 281691 126928
rect 227897 126923 227963 126926
rect 281625 126923 281691 126926
rect 66805 126850 66871 126853
rect 66805 126848 68908 126850
rect 66805 126792 66810 126848
rect 66866 126792 68908 126848
rect 66805 126790 68908 126792
rect 66805 126787 66871 126790
rect 191557 126578 191623 126581
rect 226701 126578 226767 126581
rect 191557 126576 193660 126578
rect 191557 126520 191562 126576
rect 191618 126520 193660 126576
rect 191557 126518 193660 126520
rect 224940 126576 226767 126578
rect 224940 126520 226706 126576
rect 226762 126520 226767 126576
rect 224940 126518 226767 126520
rect 191557 126515 191623 126518
rect 226701 126515 226767 126518
rect 95969 126442 96035 126445
rect 95969 126440 103530 126442
rect 95969 126384 95974 126440
rect 96030 126384 103530 126440
rect 95969 126382 103530 126384
rect 95969 126379 96035 126382
rect 97901 126306 97967 126309
rect 94668 126304 97967 126306
rect 94668 126248 97906 126304
rect 97962 126248 97967 126304
rect 94668 126246 97967 126248
rect 103470 126306 103530 126382
rect 184749 126306 184815 126309
rect 103470 126304 184815 126306
rect 103470 126248 184754 126304
rect 184810 126248 184815 126304
rect 103470 126246 184815 126248
rect 97901 126243 97967 126246
rect 184749 126243 184815 126246
rect 66069 126034 66135 126037
rect 583109 126034 583175 126037
rect 583520 126034 584960 126124
rect 66069 126032 68908 126034
rect 66069 125976 66074 126032
rect 66130 125976 68908 126032
rect 66069 125974 68908 125976
rect 583109 126032 584960 126034
rect 583109 125976 583114 126032
rect 583170 125976 584960 126032
rect 583109 125974 584960 125976
rect 66069 125971 66135 125974
rect 583109 125971 583175 125974
rect 583520 125884 584960 125974
rect 184749 125762 184815 125765
rect 190269 125762 190335 125765
rect 227897 125762 227963 125765
rect 184749 125760 193660 125762
rect 184749 125704 184754 125760
rect 184810 125704 190274 125760
rect 190330 125704 193660 125760
rect 184749 125702 193660 125704
rect 224940 125760 227963 125762
rect 224940 125704 227902 125760
rect 227958 125704 227963 125760
rect 224940 125702 227963 125704
rect 184749 125699 184815 125702
rect 190269 125699 190335 125702
rect 227897 125699 227963 125702
rect 97809 125490 97875 125493
rect 94668 125488 97875 125490
rect 94668 125432 97814 125488
rect 97870 125432 97875 125488
rect 94668 125430 97875 125432
rect 97809 125427 97875 125430
rect 68878 124674 68938 125188
rect 192477 124946 192543 124949
rect 192477 124944 193660 124946
rect 192477 124888 192482 124944
rect 192538 124888 193660 124944
rect 192477 124886 193660 124888
rect 192477 124883 192543 124886
rect 100753 124810 100819 124813
rect 102225 124810 102291 124813
rect 169293 124810 169359 124813
rect 100753 124808 169359 124810
rect 100753 124752 100758 124808
rect 100814 124752 102230 124808
rect 102286 124752 169298 124808
rect 169354 124752 169359 124808
rect 100753 124750 169359 124752
rect 100753 124747 100819 124750
rect 102225 124747 102291 124750
rect 169293 124747 169359 124750
rect 97901 124674 97967 124677
rect 226609 124674 226675 124677
rect 64830 124614 68938 124674
rect 94668 124672 97967 124674
rect 94668 124616 97906 124672
rect 97962 124616 97967 124672
rect 94668 124614 97967 124616
rect 224940 124672 226675 124674
rect 224940 124616 226614 124672
rect 226670 124616 226675 124672
rect 224940 124614 226675 124616
rect 63217 124402 63283 124405
rect 64830 124402 64890 124614
rect 97901 124611 97967 124614
rect 226609 124611 226675 124614
rect 63217 124400 64890 124402
rect 63217 124344 63222 124400
rect 63278 124344 64890 124400
rect 63217 124342 64890 124344
rect 66805 124402 66871 124405
rect 66805 124400 68908 124402
rect 66805 124344 66810 124400
rect 66866 124344 68908 124400
rect 66805 124342 68908 124344
rect 63217 124339 63283 124342
rect 66805 124339 66871 124342
rect 97901 124130 97967 124133
rect 94668 124128 97967 124130
rect 94668 124072 97906 124128
rect 97962 124072 97967 124128
rect 94668 124070 97967 124072
rect 97901 124067 97967 124070
rect 124949 124130 125015 124133
rect 124949 124128 180810 124130
rect 124949 124072 124954 124128
rect 125010 124072 180810 124128
rect 124949 124070 180810 124072
rect 124949 124067 125015 124070
rect 66989 123858 67055 123861
rect 180750 123858 180810 124070
rect 192334 123858 192340 123860
rect 66989 123856 68908 123858
rect -960 123572 480 123812
rect 66989 123800 66994 123856
rect 67050 123800 68908 123856
rect 66989 123798 68908 123800
rect 180750 123798 192340 123858
rect 66989 123795 67055 123798
rect 192334 123796 192340 123798
rect 192404 123858 192410 123860
rect 192937 123858 193003 123861
rect 227621 123858 227687 123861
rect 192404 123856 193660 123858
rect 192404 123800 192942 123856
rect 192998 123800 193660 123856
rect 192404 123798 193660 123800
rect 224940 123856 227687 123858
rect 224940 123800 227626 123856
rect 227682 123800 227687 123856
rect 224940 123798 227687 123800
rect 192404 123796 192410 123798
rect 192937 123795 193003 123798
rect 227621 123795 227687 123798
rect 97165 123314 97231 123317
rect 94668 123312 97231 123314
rect 94668 123256 97170 123312
rect 97226 123256 97231 123312
rect 94668 123254 97231 123256
rect 97165 123251 97231 123254
rect 66897 123042 66963 123045
rect 191741 123042 191807 123045
rect 226701 123042 226767 123045
rect 66897 123040 68908 123042
rect 66897 122984 66902 123040
rect 66958 122984 68908 123040
rect 66897 122982 68908 122984
rect 191741 123040 193660 123042
rect 191741 122984 191746 123040
rect 191802 122984 193660 123040
rect 191741 122982 193660 122984
rect 224940 123040 226767 123042
rect 224940 122984 226706 123040
rect 226762 122984 226767 123040
rect 224940 122982 226767 122984
rect 66897 122979 66963 122982
rect 191741 122979 191807 122982
rect 226701 122979 226767 122982
rect 97349 122498 97415 122501
rect 94668 122496 97415 122498
rect 94668 122440 97354 122496
rect 97410 122440 97415 122496
rect 94668 122438 97415 122440
rect 97349 122435 97415 122438
rect 66345 122226 66411 122229
rect 191741 122226 191807 122229
rect 226517 122226 226583 122229
rect 66345 122224 68908 122226
rect 66345 122168 66350 122224
rect 66406 122168 68908 122224
rect 66345 122166 68908 122168
rect 191741 122224 193660 122226
rect 191741 122168 191746 122224
rect 191802 122168 193660 122224
rect 191741 122166 193660 122168
rect 224940 122224 226583 122226
rect 224940 122168 226522 122224
rect 226578 122168 226583 122224
rect 224940 122166 226583 122168
rect 66345 122163 66411 122166
rect 191741 122163 191807 122166
rect 226517 122163 226583 122166
rect 97901 121682 97967 121685
rect 94668 121680 97967 121682
rect 94668 121624 97906 121680
rect 97962 121624 97967 121680
rect 94668 121622 97967 121624
rect 97901 121619 97967 121622
rect 66805 121410 66871 121413
rect 191189 121410 191255 121413
rect 66805 121408 68908 121410
rect 66805 121352 66810 121408
rect 66866 121352 68908 121408
rect 66805 121350 68908 121352
rect 191189 121408 193660 121410
rect 191189 121352 191194 121408
rect 191250 121352 193660 121408
rect 191189 121350 193660 121352
rect 66805 121347 66871 121350
rect 191189 121347 191255 121350
rect 224902 121348 224908 121412
rect 224972 121348 224978 121412
rect 224910 121108 224970 121348
rect 97073 120866 97139 120869
rect 94668 120864 97139 120866
rect 94668 120808 97078 120864
rect 97134 120808 97139 120864
rect 94668 120806 97139 120808
rect 97073 120803 97139 120806
rect 66897 120594 66963 120597
rect 66897 120592 68908 120594
rect 66897 120536 66902 120592
rect 66958 120536 68908 120592
rect 66897 120534 68908 120536
rect 66897 120531 66963 120534
rect 95325 120322 95391 120325
rect 96061 120322 96127 120325
rect 94668 120320 96127 120322
rect 94668 120264 95330 120320
rect 95386 120264 96066 120320
rect 96122 120264 96127 120320
rect 94668 120262 96127 120264
rect 95325 120259 95391 120262
rect 96061 120259 96127 120262
rect 191005 120322 191071 120325
rect 226701 120322 226767 120325
rect 191005 120320 193660 120322
rect 191005 120264 191010 120320
rect 191066 120264 193660 120320
rect 191005 120262 193660 120264
rect 224940 120320 226767 120322
rect 224940 120264 226706 120320
rect 226762 120264 226767 120320
rect 224940 120262 226767 120264
rect 191005 120259 191071 120262
rect 226701 120259 226767 120262
rect 66805 120050 66871 120053
rect 66805 120048 68908 120050
rect 66805 119992 66810 120048
rect 66866 119992 68908 120048
rect 66805 119990 68908 119992
rect 66805 119987 66871 119990
rect 97901 119506 97967 119509
rect 94668 119504 97967 119506
rect 94668 119448 97906 119504
rect 97962 119448 97967 119504
rect 94668 119446 97967 119448
rect 97901 119443 97967 119446
rect 191741 119506 191807 119509
rect 226374 119506 226380 119508
rect 191741 119504 193660 119506
rect 191741 119448 191746 119504
rect 191802 119448 193660 119504
rect 191741 119446 193660 119448
rect 224940 119446 226380 119506
rect 191741 119443 191807 119446
rect 226374 119444 226380 119446
rect 226444 119444 226450 119508
rect 106774 119308 106780 119372
rect 106844 119370 106850 119372
rect 127617 119370 127683 119373
rect 106844 119368 127683 119370
rect 106844 119312 127622 119368
rect 127678 119312 127683 119368
rect 106844 119310 127683 119312
rect 106844 119308 106850 119310
rect 127617 119307 127683 119310
rect 66897 119234 66963 119237
rect 66897 119232 68908 119234
rect 66897 119176 66902 119232
rect 66958 119176 68908 119232
rect 66897 119174 68908 119176
rect 66897 119171 66963 119174
rect 97901 118690 97967 118693
rect 94668 118688 97967 118690
rect 94668 118632 97906 118688
rect 97962 118632 97967 118688
rect 94668 118630 97967 118632
rect 97901 118627 97967 118630
rect 191741 118690 191807 118693
rect 191741 118688 193660 118690
rect 191741 118632 191746 118688
rect 191802 118632 193660 118688
rect 191741 118630 193660 118632
rect 191741 118627 191807 118630
rect 67817 118418 67883 118421
rect 226517 118418 226583 118421
rect 67817 118416 68908 118418
rect 67817 118360 67822 118416
rect 67878 118360 68908 118416
rect 67817 118358 68908 118360
rect 224940 118416 226583 118418
rect 224940 118360 226522 118416
rect 226578 118360 226583 118416
rect 224940 118358 226583 118360
rect 67817 118355 67883 118358
rect 226517 118355 226583 118358
rect 127617 118010 127683 118013
rect 144177 118010 144243 118013
rect 127617 118008 144243 118010
rect 127617 117952 127622 118008
rect 127678 117952 144182 118008
rect 144238 117952 144243 118008
rect 127617 117950 144243 117952
rect 127617 117947 127683 117950
rect 144177 117947 144243 117950
rect 102777 117874 102843 117877
rect 94668 117872 102843 117874
rect 94668 117816 102782 117872
rect 102838 117816 102843 117872
rect 94668 117814 102843 117816
rect 102777 117811 102843 117814
rect 66621 117602 66687 117605
rect 191097 117602 191163 117605
rect 226609 117602 226675 117605
rect 66621 117600 68908 117602
rect 66621 117544 66626 117600
rect 66682 117544 68908 117600
rect 66621 117542 68908 117544
rect 191097 117600 193660 117602
rect 191097 117544 191102 117600
rect 191158 117544 193660 117600
rect 191097 117542 193660 117544
rect 224940 117600 226675 117602
rect 224940 117544 226614 117600
rect 226670 117544 226675 117600
rect 224940 117542 226675 117544
rect 66621 117539 66687 117542
rect 191097 117539 191163 117542
rect 226609 117539 226675 117542
rect 65926 116996 65932 117060
rect 65996 117058 66002 117060
rect 97901 117058 97967 117061
rect 65996 116998 68908 117058
rect 94668 117056 97967 117058
rect 94668 117000 97906 117056
rect 97962 117000 97967 117056
rect 94668 116998 97967 117000
rect 65996 116996 66002 116998
rect 97901 116995 97967 116998
rect 191557 116786 191623 116789
rect 227621 116786 227687 116789
rect 191557 116784 193660 116786
rect 191557 116728 191562 116784
rect 191618 116728 193660 116784
rect 191557 116726 193660 116728
rect 224940 116784 227687 116786
rect 224940 116728 227626 116784
rect 227682 116728 227687 116784
rect 224940 116726 227687 116728
rect 191557 116723 191623 116726
rect 227621 116723 227687 116726
rect 97349 116514 97415 116517
rect 94668 116512 97415 116514
rect 94668 116456 97354 116512
rect 97410 116456 97415 116512
rect 94668 116454 97415 116456
rect 97349 116451 97415 116454
rect 171961 116514 172027 116517
rect 189809 116514 189875 116517
rect 171961 116512 189875 116514
rect 171961 116456 171966 116512
rect 172022 116456 189814 116512
rect 189870 116456 189875 116512
rect 171961 116454 189875 116456
rect 171961 116451 172027 116454
rect 189809 116451 189875 116454
rect 66621 116242 66687 116245
rect 66621 116240 68908 116242
rect 66621 116184 66626 116240
rect 66682 116184 68908 116240
rect 66621 116182 68908 116184
rect 66621 116179 66687 116182
rect 189717 115970 189783 115973
rect 226701 115970 226767 115973
rect 189717 115968 193660 115970
rect 189717 115912 189722 115968
rect 189778 115912 193660 115968
rect 189717 115910 193660 115912
rect 224940 115968 226767 115970
rect 224940 115912 226706 115968
rect 226762 115912 226767 115968
rect 224940 115910 226767 115912
rect 189717 115907 189783 115910
rect 226701 115907 226767 115910
rect 97901 115698 97967 115701
rect 94668 115696 97967 115698
rect 94668 115640 97906 115696
rect 97962 115640 97967 115696
rect 94668 115638 97967 115640
rect 97901 115635 97967 115638
rect 66805 115426 66871 115429
rect 66805 115424 68908 115426
rect 66805 115368 66810 115424
rect 66866 115368 68908 115424
rect 66805 115366 68908 115368
rect 66805 115363 66871 115366
rect 191741 115154 191807 115157
rect 191741 115152 193660 115154
rect 191741 115096 191746 115152
rect 191802 115096 193660 115152
rect 191741 115094 193660 115096
rect 191741 115091 191807 115094
rect 97809 114882 97875 114885
rect 225137 114882 225203 114885
rect 226149 114882 226215 114885
rect 94668 114880 97875 114882
rect 94668 114824 97814 114880
rect 97870 114824 97875 114880
rect 94668 114822 97875 114824
rect 224940 114880 226215 114882
rect 224940 114824 225142 114880
rect 225198 114824 226154 114880
rect 226210 114824 226215 114880
rect 224940 114822 226215 114824
rect 97809 114819 97875 114822
rect 225137 114819 225203 114822
rect 226149 114819 226215 114822
rect 66897 114610 66963 114613
rect 66897 114608 68908 114610
rect 66897 114552 66902 114608
rect 66958 114552 68908 114608
rect 66897 114550 68908 114552
rect 66897 114547 66963 114550
rect 97257 114066 97323 114069
rect 94668 114064 97323 114066
rect 94668 114008 97262 114064
rect 97318 114008 97323 114064
rect 94668 114006 97323 114008
rect 97257 114003 97323 114006
rect 191833 114066 191899 114069
rect 226425 114066 226491 114069
rect 191833 114064 193660 114066
rect 191833 114008 191838 114064
rect 191894 114008 193660 114064
rect 191833 114006 193660 114008
rect 224940 114064 226491 114066
rect 224940 114008 226430 114064
rect 226486 114008 226491 114064
rect 224940 114006 226491 114008
rect 191833 114003 191899 114006
rect 226425 114003 226491 114006
rect 66805 113794 66871 113797
rect 225045 113794 225111 113797
rect 66805 113792 68908 113794
rect 66805 113736 66810 113792
rect 66866 113736 68908 113792
rect 66805 113734 68908 113736
rect 224910 113792 225111 113794
rect 224910 113736 225050 113792
rect 225106 113736 225111 113792
rect 224910 113734 225111 113736
rect 66805 113731 66871 113734
rect 97533 113522 97599 113525
rect 94668 113520 97599 113522
rect 94668 113464 97538 113520
rect 97594 113464 97599 113520
rect 94668 113462 97599 113464
rect 97533 113459 97599 113462
rect 66897 113250 66963 113253
rect 191741 113250 191807 113253
rect 66897 113248 68908 113250
rect 66897 113192 66902 113248
rect 66958 113192 68908 113248
rect 66897 113190 68908 113192
rect 191741 113248 193660 113250
rect 191741 113192 191746 113248
rect 191802 113192 193660 113248
rect 224910 113220 224970 113734
rect 225045 113731 225111 113734
rect 191741 113190 193660 113192
rect 66897 113187 66963 113190
rect 191741 113187 191807 113190
rect 582925 112842 582991 112845
rect 583520 112842 584960 112932
rect 582925 112840 584960 112842
rect 582925 112784 582930 112840
rect 582986 112784 584960 112840
rect 582925 112782 584960 112784
rect 582925 112779 582991 112782
rect 97901 112706 97967 112709
rect 94668 112704 97967 112706
rect 94668 112648 97906 112704
rect 97962 112648 97967 112704
rect 583520 112692 584960 112782
rect 94668 112646 97967 112648
rect 97901 112643 97967 112646
rect 66805 112434 66871 112437
rect 191741 112434 191807 112437
rect 66805 112432 68908 112434
rect 66805 112376 66810 112432
rect 66866 112376 68908 112432
rect 66805 112374 68908 112376
rect 191741 112432 193660 112434
rect 191741 112376 191746 112432
rect 191802 112376 193660 112432
rect 191741 112374 193660 112376
rect 66805 112371 66871 112374
rect 191741 112371 191807 112374
rect 226333 112162 226399 112165
rect 224940 112160 226399 112162
rect 224940 112104 226338 112160
rect 226394 112104 226399 112160
rect 224940 112102 226399 112104
rect 226333 112099 226399 112102
rect 96705 111890 96771 111893
rect 94668 111888 96771 111890
rect 94668 111832 96710 111888
rect 96766 111832 96771 111888
rect 94668 111830 96771 111832
rect 96705 111827 96771 111830
rect 97349 111890 97415 111893
rect 104985 111890 105051 111893
rect 97349 111888 105051 111890
rect 97349 111832 97354 111888
rect 97410 111832 104990 111888
rect 105046 111832 105051 111888
rect 97349 111830 105051 111832
rect 97349 111827 97415 111830
rect 104985 111827 105051 111830
rect 66805 111618 66871 111621
rect 66805 111616 68908 111618
rect 66805 111560 66810 111616
rect 66866 111560 68908 111616
rect 66805 111558 68908 111560
rect 66805 111555 66871 111558
rect 226701 111346 226767 111349
rect 224940 111344 226767 111346
rect 96797 111074 96863 111077
rect 94668 111072 96863 111074
rect 94668 111016 96802 111072
rect 96858 111016 96863 111072
rect 94668 111014 96863 111016
rect 96797 111011 96863 111014
rect 66897 110802 66963 110805
rect 189073 110802 189139 110805
rect 193630 110802 193690 111316
rect 224940 111288 226706 111344
rect 226762 111288 226767 111344
rect 224940 111286 226767 111288
rect 226701 111283 226767 111286
rect 66897 110800 68908 110802
rect -960 110666 480 110756
rect 66897 110744 66902 110800
rect 66958 110744 68908 110800
rect 66897 110742 68908 110744
rect 189073 110800 193690 110802
rect 189073 110744 189078 110800
rect 189134 110744 193690 110800
rect 189073 110742 193690 110744
rect 66897 110739 66963 110742
rect 189073 110739 189139 110742
rect 2865 110666 2931 110669
rect -960 110664 2931 110666
rect -960 110608 2870 110664
rect 2926 110608 2931 110664
rect -960 110606 2931 110608
rect -960 110516 480 110606
rect 2865 110603 2931 110606
rect 191741 110530 191807 110533
rect 226333 110530 226399 110533
rect 191741 110528 193660 110530
rect 191741 110472 191746 110528
rect 191802 110472 193660 110528
rect 191741 110470 193660 110472
rect 224940 110528 226399 110530
rect 224940 110472 226338 110528
rect 226394 110472 226399 110528
rect 224940 110470 226399 110472
rect 191741 110467 191807 110470
rect 226333 110467 226399 110470
rect 66897 110258 66963 110261
rect 97809 110258 97875 110261
rect 66897 110256 68908 110258
rect 66897 110200 66902 110256
rect 66958 110200 68908 110256
rect 66897 110198 68908 110200
rect 94668 110256 97875 110258
rect 94668 110200 97814 110256
rect 97870 110200 97875 110256
rect 94668 110198 97875 110200
rect 66897 110195 66963 110198
rect 97809 110195 97875 110198
rect 97901 109714 97967 109717
rect 94668 109712 97967 109714
rect 94668 109656 97906 109712
rect 97962 109656 97967 109712
rect 94668 109654 97967 109656
rect 97901 109651 97967 109654
rect 190637 109714 190703 109717
rect 190637 109712 193660 109714
rect 190637 109656 190642 109712
rect 190698 109656 193660 109712
rect 190637 109654 193660 109656
rect 190637 109651 190703 109654
rect 66478 109380 66484 109444
rect 66548 109442 66554 109444
rect 66548 109382 68908 109442
rect 66548 109380 66554 109382
rect 94078 109108 94084 109172
rect 94148 109108 94154 109172
rect 224910 109170 224970 109684
rect 225045 109170 225111 109173
rect 224910 109168 225111 109170
rect 224910 109112 225050 109168
rect 225106 109112 225111 109168
rect 224910 109110 225111 109112
rect 94086 108868 94146 109108
rect 225045 109107 225111 109110
rect 191741 108898 191807 108901
rect 191741 108896 193660 108898
rect 191741 108840 191746 108896
rect 191802 108840 193660 108896
rect 191741 108838 193660 108840
rect 191741 108835 191807 108838
rect 66069 108626 66135 108629
rect 226517 108626 226583 108629
rect 66069 108624 68908 108626
rect 66069 108568 66074 108624
rect 66130 108568 68908 108624
rect 66069 108566 68908 108568
rect 224940 108624 226583 108626
rect 224940 108568 226522 108624
rect 226578 108568 226583 108624
rect 224940 108566 226583 108568
rect 66069 108563 66135 108566
rect 226517 108563 226583 108566
rect 227662 108354 227668 108356
rect 224910 108294 227668 108354
rect 97901 108082 97967 108085
rect 94668 108080 97967 108082
rect 94668 108024 97906 108080
rect 97962 108024 97967 108080
rect 94668 108022 97967 108024
rect 97901 108019 97967 108022
rect 66805 107810 66871 107813
rect 188429 107810 188495 107813
rect 188838 107810 188844 107812
rect 66805 107808 68908 107810
rect 66805 107752 66810 107808
rect 66866 107752 68908 107808
rect 66805 107750 68908 107752
rect 188429 107808 188844 107810
rect 188429 107752 188434 107808
rect 188490 107752 188844 107808
rect 188429 107750 188844 107752
rect 66805 107747 66871 107750
rect 188429 107747 188495 107750
rect 188838 107748 188844 107750
rect 188908 107810 188914 107812
rect 188908 107750 193660 107810
rect 224910 107780 224970 108294
rect 227662 108292 227668 108294
rect 227732 108354 227738 108356
rect 270534 108354 270540 108356
rect 227732 108294 270540 108354
rect 227732 108292 227738 108294
rect 270534 108292 270540 108294
rect 270604 108292 270610 108356
rect 188908 107748 188914 107750
rect 97901 107266 97967 107269
rect 94668 107264 97967 107266
rect 94668 107208 97906 107264
rect 97962 107208 97967 107264
rect 94668 107206 97967 107208
rect 97901 107203 97967 107206
rect 66662 106932 66668 106996
rect 66732 106994 66738 106996
rect 66805 106994 66871 106997
rect 190821 106994 190887 106997
rect 226701 106994 226767 106997
rect 66732 106992 68908 106994
rect 66732 106936 66810 106992
rect 66866 106936 68908 106992
rect 66732 106934 68908 106936
rect 190821 106992 193660 106994
rect 190821 106936 190826 106992
rect 190882 106936 193660 106992
rect 190821 106934 193660 106936
rect 224940 106992 226767 106994
rect 224940 106936 226706 106992
rect 226762 106936 226767 106992
rect 224940 106934 226767 106936
rect 66732 106932 66738 106934
rect 66805 106931 66871 106934
rect 190821 106931 190887 106934
rect 226701 106931 226767 106934
rect 97901 106722 97967 106725
rect 94668 106720 97967 106722
rect 94668 106664 97906 106720
rect 97962 106664 97967 106720
rect 94668 106662 97967 106664
rect 97901 106659 97967 106662
rect 66621 106450 66687 106453
rect 66621 106448 68908 106450
rect 66621 106392 66626 106448
rect 66682 106392 68908 106448
rect 66621 106390 68908 106392
rect 66621 106387 66687 106390
rect 94262 106116 94268 106180
rect 94332 106116 94338 106180
rect 191189 106178 191255 106181
rect 191189 106176 193660 106178
rect 191189 106120 191194 106176
rect 191250 106120 193660 106176
rect 191189 106118 193660 106120
rect 94270 105876 94330 106116
rect 191189 106115 191255 106118
rect 226333 105906 226399 105909
rect 224940 105904 226399 105906
rect 224940 105848 226338 105904
rect 226394 105848 226399 105904
rect 224940 105846 226399 105848
rect 226333 105843 226399 105846
rect 66621 105634 66687 105637
rect 66621 105632 68908 105634
rect 66621 105576 66626 105632
rect 66682 105576 68908 105632
rect 66621 105574 68908 105576
rect 66621 105571 66687 105574
rect 98494 105090 98500 105092
rect 94668 105030 98500 105090
rect 98494 105028 98500 105030
rect 98564 105028 98570 105092
rect 191741 105090 191807 105093
rect 226701 105090 226767 105093
rect 191741 105088 193660 105090
rect 191741 105032 191746 105088
rect 191802 105032 193660 105088
rect 191741 105030 193660 105032
rect 224940 105088 226767 105090
rect 224940 105032 226706 105088
rect 226762 105032 226767 105088
rect 224940 105030 226767 105032
rect 191741 105027 191807 105030
rect 226701 105027 226767 105030
rect 66805 104818 66871 104821
rect 66805 104816 68908 104818
rect 66805 104760 66810 104816
rect 66866 104760 68908 104816
rect 66805 104758 68908 104760
rect 66805 104755 66871 104758
rect 97901 104274 97967 104277
rect 94668 104272 97967 104274
rect 94668 104216 97906 104272
rect 97962 104216 97967 104272
rect 94668 104214 97967 104216
rect 97901 104211 97967 104214
rect 193213 104274 193279 104277
rect 226701 104274 226767 104277
rect 193213 104272 193660 104274
rect 193213 104216 193218 104272
rect 193274 104216 193660 104272
rect 193213 104214 193660 104216
rect 224940 104272 226767 104274
rect 224940 104216 226706 104272
rect 226762 104216 226767 104272
rect 224940 104214 226767 104216
rect 193213 104211 193279 104214
rect 226701 104211 226767 104214
rect 67265 104002 67331 104005
rect 67265 104000 68908 104002
rect 67265 103944 67270 104000
rect 67326 103944 68908 104000
rect 67265 103942 68908 103944
rect 67265 103939 67331 103942
rect 98637 103594 98703 103597
rect 104014 103594 104020 103596
rect 98637 103592 104020 103594
rect 98637 103536 98642 103592
rect 98698 103536 104020 103592
rect 98637 103534 104020 103536
rect 98637 103531 98703 103534
rect 104014 103532 104020 103534
rect 104084 103532 104090 103596
rect 97901 103458 97967 103461
rect 94668 103456 97967 103458
rect 94668 103400 97906 103456
rect 97962 103400 97967 103456
rect 94668 103398 97967 103400
rect 97901 103395 97967 103398
rect 191005 103458 191071 103461
rect 226701 103458 226767 103461
rect 191005 103456 193660 103458
rect 191005 103400 191010 103456
rect 191066 103400 193660 103456
rect 191005 103398 193660 103400
rect 224940 103456 226767 103458
rect 224940 103400 226706 103456
rect 226762 103400 226767 103456
rect 224940 103398 226767 103400
rect 191005 103395 191071 103398
rect 226701 103395 226767 103398
rect 65885 103186 65951 103189
rect 65885 103184 68908 103186
rect 65885 103128 65890 103184
rect 65946 103128 68908 103184
rect 65885 103126 68908 103128
rect 65885 103123 65951 103126
rect 97901 102914 97967 102917
rect 94668 102912 97967 102914
rect 94668 102856 97906 102912
rect 97962 102856 97967 102912
rect 94668 102854 97967 102856
rect 97901 102851 97967 102854
rect 66437 102642 66503 102645
rect 193121 102642 193187 102645
rect 66437 102640 68908 102642
rect 66437 102584 66442 102640
rect 66498 102584 68908 102640
rect 66437 102582 68908 102584
rect 193121 102640 193844 102642
rect 193121 102584 193126 102640
rect 193182 102612 193844 102640
rect 193182 102584 193874 102612
rect 193121 102582 193874 102584
rect 66437 102579 66503 102582
rect 193121 102579 193187 102582
rect 100017 102234 100083 102237
rect 171869 102234 171935 102237
rect 172421 102234 172487 102237
rect 193814 102236 193874 102582
rect 226701 102370 226767 102373
rect 224940 102368 226767 102370
rect 224940 102312 226706 102368
rect 226762 102312 226767 102368
rect 224940 102310 226767 102312
rect 226701 102307 226767 102310
rect 100017 102232 172487 102234
rect 100017 102176 100022 102232
rect 100078 102176 171874 102232
rect 171930 102176 172426 102232
rect 172482 102176 172487 102232
rect 100017 102174 172487 102176
rect 100017 102171 100083 102174
rect 171869 102171 171935 102174
rect 172421 102171 172487 102174
rect 193806 102172 193812 102236
rect 193876 102172 193882 102236
rect 97901 102098 97967 102101
rect 94668 102096 97967 102098
rect 94668 102040 97906 102096
rect 97962 102040 97967 102096
rect 94668 102038 97967 102040
rect 97901 102035 97967 102038
rect 66713 101826 66779 101829
rect 66713 101824 68908 101826
rect 66713 101768 66718 101824
rect 66774 101768 68908 101824
rect 66713 101766 68908 101768
rect 66713 101763 66779 101766
rect 191741 101554 191807 101557
rect 226333 101554 226399 101557
rect 191741 101552 193660 101554
rect 191741 101496 191746 101552
rect 191802 101496 193660 101552
rect 191741 101494 193660 101496
rect 224940 101552 226399 101554
rect 224940 101496 226338 101552
rect 226394 101496 226399 101552
rect 224940 101494 226399 101496
rect 191741 101491 191807 101494
rect 226333 101491 226399 101494
rect 97901 101282 97967 101285
rect 94668 101280 97967 101282
rect 94668 101224 97906 101280
rect 97962 101224 97967 101280
rect 94668 101222 97967 101224
rect 97901 101219 97967 101222
rect 66805 101010 66871 101013
rect 66805 101008 68908 101010
rect 66805 100952 66810 101008
rect 66866 100952 68908 101008
rect 66805 100950 68908 100952
rect 66805 100947 66871 100950
rect 191649 100738 191715 100741
rect 227897 100738 227963 100741
rect 191649 100736 193660 100738
rect 191649 100680 191654 100736
rect 191710 100680 193660 100736
rect 191649 100678 193660 100680
rect 224940 100736 227963 100738
rect 224940 100680 227902 100736
rect 227958 100680 227963 100736
rect 224940 100678 227963 100680
rect 191649 100675 191715 100678
rect 227897 100675 227963 100678
rect 97533 100466 97599 100469
rect 94668 100464 97599 100466
rect 94668 100408 97538 100464
rect 97594 100408 97599 100464
rect 94668 100406 97599 100408
rect 97533 100403 97599 100406
rect 67449 100194 67515 100197
rect 67449 100192 68908 100194
rect 67449 100136 67454 100192
rect 67510 100136 68908 100192
rect 67449 100134 68908 100136
rect 67449 100131 67515 100134
rect 66805 99650 66871 99653
rect 97901 99650 97967 99653
rect 66805 99648 68908 99650
rect 66805 99592 66810 99648
rect 66866 99592 68908 99648
rect 66805 99590 68908 99592
rect 94668 99648 97967 99650
rect 94668 99592 97906 99648
rect 97962 99592 97967 99648
rect 94668 99590 97967 99592
rect 66805 99587 66871 99590
rect 97901 99587 97967 99590
rect 189809 99650 189875 99653
rect 193630 99650 193690 99892
rect 189809 99648 193690 99650
rect 189809 99592 189814 99648
rect 189870 99592 193690 99648
rect 189809 99590 193690 99592
rect 189809 99587 189875 99590
rect 190177 99514 190243 99517
rect 191649 99514 191715 99517
rect 224358 99516 224418 99620
rect 190177 99512 191715 99514
rect 190177 99456 190182 99512
rect 190238 99456 191654 99512
rect 191710 99456 191715 99512
rect 190177 99454 191715 99456
rect 190177 99451 190243 99454
rect 191649 99451 191715 99454
rect 224350 99452 224356 99516
rect 224420 99514 224426 99516
rect 226333 99514 226399 99517
rect 224420 99512 226399 99514
rect 224420 99456 226338 99512
rect 226394 99456 226399 99512
rect 224420 99454 226399 99456
rect 224420 99452 224426 99454
rect 226333 99451 226399 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 98913 99106 98979 99109
rect 94668 99104 98979 99106
rect 94668 99048 98918 99104
rect 98974 99048 98979 99104
rect 94668 99046 98979 99048
rect 98913 99043 98979 99046
rect 66805 98834 66871 98837
rect 226701 98834 226767 98837
rect 66805 98832 68908 98834
rect 66805 98776 66810 98832
rect 66866 98776 68908 98832
rect 224940 98832 226767 98834
rect 66805 98774 68908 98776
rect 66805 98771 66871 98774
rect 94773 98562 94839 98565
rect 193630 98562 193690 98804
rect 224940 98776 226706 98832
rect 226762 98776 226767 98832
rect 224940 98774 226767 98776
rect 226701 98771 226767 98774
rect 94773 98560 193690 98562
rect 94773 98504 94778 98560
rect 94834 98504 193690 98560
rect 94773 98502 193690 98504
rect 94773 98499 94839 98502
rect 97901 98290 97967 98293
rect 94668 98288 97967 98290
rect 94668 98232 97906 98288
rect 97962 98232 97967 98288
rect 94668 98230 97967 98232
rect 97901 98227 97967 98230
rect 67357 98018 67423 98021
rect 191741 98018 191807 98021
rect 226609 98018 226675 98021
rect 67357 98016 68908 98018
rect 67357 97960 67362 98016
rect 67418 97960 68908 98016
rect 67357 97958 68908 97960
rect 191741 98016 193660 98018
rect 191741 97960 191746 98016
rect 191802 97960 193660 98016
rect 191741 97958 193660 97960
rect 224940 98016 226675 98018
rect 224940 97960 226614 98016
rect 226670 97960 226675 98016
rect 224940 97958 226675 97960
rect 67357 97955 67423 97958
rect 191741 97955 191807 97958
rect 226609 97955 226675 97958
rect -960 97610 480 97700
rect 3049 97610 3115 97613
rect -960 97608 3115 97610
rect -960 97552 3054 97608
rect 3110 97552 3115 97608
rect -960 97550 3115 97552
rect -960 97460 480 97550
rect 3049 97547 3115 97550
rect 67357 97202 67423 97205
rect 67541 97202 67607 97205
rect 67357 97200 68908 97202
rect 67357 97144 67362 97200
rect 67418 97144 67546 97200
rect 67602 97144 68908 97200
rect 67357 97142 68908 97144
rect 67357 97139 67423 97142
rect 67541 97139 67607 97142
rect 94638 96930 94698 97444
rect 191649 97202 191715 97205
rect 226374 97202 226380 97204
rect 191649 97200 193660 97202
rect 191649 97144 191654 97200
rect 191710 97144 193660 97200
rect 191649 97142 193660 97144
rect 224940 97142 226380 97202
rect 191649 97139 191715 97142
rect 226374 97140 226380 97142
rect 226444 97202 226450 97204
rect 226977 97202 227043 97205
rect 226444 97200 227043 97202
rect 226444 97144 226982 97200
rect 227038 97144 227043 97200
rect 226444 97142 227043 97144
rect 226444 97140 226450 97142
rect 226977 97139 227043 97142
rect 189942 96930 189948 96932
rect 94638 96870 189948 96930
rect 189942 96868 189948 96870
rect 190012 96868 190018 96932
rect 96705 96658 96771 96661
rect 94668 96656 96771 96658
rect 94668 96600 96710 96656
rect 96766 96600 96771 96656
rect 94668 96598 96771 96600
rect 96705 96595 96771 96598
rect 66110 96324 66116 96388
rect 66180 96386 66186 96388
rect 66180 96326 68908 96386
rect 66180 96324 66186 96326
rect 97206 96114 97212 96116
rect 94668 96054 97212 96114
rect 97206 96052 97212 96054
rect 97276 96052 97282 96116
rect 67541 95842 67607 95845
rect 67541 95840 68908 95842
rect 67541 95784 67546 95840
rect 67602 95784 68908 95840
rect 67541 95782 68908 95784
rect 67541 95779 67607 95782
rect 94814 95780 94820 95844
rect 94884 95842 94890 95844
rect 126973 95842 127039 95845
rect 94884 95840 127039 95842
rect 94884 95784 126978 95840
rect 127034 95784 127039 95840
rect 94884 95782 127039 95784
rect 94884 95780 94890 95782
rect 126973 95779 127039 95782
rect 172421 95842 172487 95845
rect 191649 95842 191715 95845
rect 193630 95842 193690 96356
rect 226701 96114 226767 96117
rect 224940 96112 226767 96114
rect 224940 96056 226706 96112
rect 226762 96056 226767 96112
rect 224940 96054 226767 96056
rect 226701 96051 226767 96054
rect 172421 95840 193690 95842
rect 172421 95784 172426 95840
rect 172482 95784 191654 95840
rect 191710 95784 193690 95840
rect 172421 95782 193690 95784
rect 264237 95842 264303 95845
rect 273294 95842 273300 95844
rect 264237 95840 273300 95842
rect 264237 95784 264242 95840
rect 264298 95784 273300 95840
rect 264237 95782 273300 95784
rect 172421 95779 172487 95782
rect 191649 95779 191715 95782
rect 264237 95779 264303 95782
rect 273294 95780 273300 95782
rect 273364 95780 273370 95844
rect 97901 95298 97967 95301
rect 94668 95296 97967 95298
rect 94668 95240 97906 95296
rect 97962 95240 97967 95296
rect 94668 95238 97967 95240
rect 97901 95235 97967 95238
rect 173801 95298 173867 95301
rect 227989 95298 228055 95301
rect 173801 95296 193660 95298
rect 173801 95240 173806 95296
rect 173862 95240 193660 95296
rect 173801 95238 193660 95240
rect 224940 95296 228055 95298
rect 224940 95240 227994 95296
rect 228050 95240 228055 95296
rect 224940 95238 228055 95240
rect 173801 95235 173867 95238
rect 227989 95235 228055 95238
rect 226425 95162 226491 95165
rect 227069 95162 227135 95165
rect 224910 95160 227135 95162
rect 224910 95104 226430 95160
rect 226486 95104 227074 95160
rect 227130 95104 227135 95160
rect 224910 95102 227135 95104
rect 66805 95026 66871 95029
rect 66805 95024 68908 95026
rect 66805 94968 66810 95024
rect 66866 94968 68908 95024
rect 66805 94966 68908 94968
rect 66805 94963 66871 94966
rect 97533 94482 97599 94485
rect 94668 94480 97599 94482
rect 94668 94424 97538 94480
rect 97594 94424 97599 94480
rect 94668 94422 97599 94424
rect 97533 94419 97599 94422
rect 164141 94482 164207 94485
rect 191741 94482 191807 94485
rect 164141 94480 193660 94482
rect 164141 94424 164146 94480
rect 164202 94424 191746 94480
rect 191802 94424 193660 94480
rect 224910 94452 224970 95102
rect 226425 95099 226491 95102
rect 227069 95099 227135 95102
rect 225137 94754 225203 94757
rect 258073 94754 258139 94757
rect 225137 94752 258139 94754
rect 225137 94696 225142 94752
rect 225198 94696 258078 94752
rect 258134 94696 258139 94752
rect 225137 94694 258139 94696
rect 225137 94691 225203 94694
rect 258073 94691 258139 94694
rect 164141 94422 193660 94424
rect 164141 94419 164207 94422
rect 191741 94419 191807 94422
rect 69430 94076 69490 94180
rect 69422 94012 69428 94076
rect 69492 94012 69498 94076
rect 97901 93666 97967 93669
rect 94668 93664 97967 93666
rect 94668 93608 97906 93664
rect 97962 93608 97967 93664
rect 94668 93606 97967 93608
rect 97901 93603 97967 93606
rect 191097 93666 191163 93669
rect 227161 93666 227227 93669
rect 191097 93664 193660 93666
rect 191097 93608 191102 93664
rect 191158 93608 193660 93664
rect 191097 93606 193660 93608
rect 224940 93664 227227 93666
rect 224940 93608 227166 93664
rect 227222 93608 227227 93664
rect 224940 93606 227227 93608
rect 191097 93603 191163 93606
rect 227161 93603 227227 93606
rect 67173 93394 67239 93397
rect 199193 93394 199259 93397
rect 200614 93394 200620 93396
rect 67173 93392 68908 93394
rect 67173 93336 67178 93392
rect 67234 93364 68908 93392
rect 199193 93392 200620 93394
rect 67234 93336 68938 93364
rect 67173 93334 68938 93336
rect 67173 93331 67239 93334
rect 68878 92850 68938 93334
rect 199193 93336 199198 93392
rect 199254 93336 200620 93392
rect 199193 93334 200620 93336
rect 199193 93331 199259 93334
rect 200614 93332 200620 93334
rect 200684 93332 200690 93396
rect 208945 93394 209011 93397
rect 209814 93394 209820 93396
rect 208945 93392 209820 93394
rect 208945 93336 208950 93392
rect 209006 93336 209820 93392
rect 208945 93334 209820 93336
rect 208945 93331 209011 93334
rect 209814 93332 209820 93334
rect 209884 93332 209890 93396
rect 102317 93258 102383 93261
rect 162761 93258 162827 93261
rect 189073 93258 189139 93261
rect 102317 93256 189139 93258
rect 102317 93200 102322 93256
rect 102378 93200 162766 93256
rect 162822 93200 189078 93256
rect 189134 93200 189139 93256
rect 102317 93198 189139 93200
rect 102317 93195 102383 93198
rect 162761 93195 162827 93198
rect 189073 93195 189139 93198
rect 101673 93122 101739 93125
rect 187693 93122 187759 93125
rect 101673 93120 187759 93122
rect 101673 93064 101678 93120
rect 101734 93064 187698 93120
rect 187754 93064 187759 93120
rect 101673 93062 187759 93064
rect 101673 93059 101739 93062
rect 187693 93059 187759 93062
rect 188797 93122 188863 93125
rect 213269 93122 213335 93125
rect 188797 93120 213335 93122
rect 188797 93064 188802 93120
rect 188858 93064 213274 93120
rect 213330 93064 213335 93120
rect 188797 93062 213335 93064
rect 188797 93059 188863 93062
rect 213269 93059 213335 93062
rect 97349 92850 97415 92853
rect 68510 92790 68938 92850
rect 94668 92848 97415 92850
rect 94668 92792 97354 92848
rect 97410 92792 97415 92848
rect 94668 92790 97415 92792
rect 68510 92717 68570 92790
rect 97349 92787 97415 92790
rect 68510 92712 68619 92717
rect 68510 92656 68558 92712
rect 68614 92656 68619 92712
rect 68510 92654 68619 92656
rect 68553 92651 68619 92654
rect 68686 92652 68692 92716
rect 68756 92714 68762 92716
rect 71175 92714 71241 92717
rect 68756 92712 71241 92714
rect 68756 92656 71180 92712
rect 71236 92656 71241 92712
rect 68756 92654 71241 92656
rect 68756 92652 68762 92654
rect 71175 92651 71241 92654
rect 72366 92652 72372 92716
rect 72436 92714 72442 92716
rect 72831 92714 72897 92717
rect 72436 92712 72897 92714
rect 72436 92656 72836 92712
rect 72892 92656 72897 92712
rect 72436 92654 72897 92656
rect 72436 92652 72442 92654
rect 72831 92651 72897 92654
rect 68870 92516 68876 92580
rect 68940 92578 68946 92580
rect 69013 92578 69079 92581
rect 69703 92578 69769 92581
rect 68940 92576 69769 92578
rect 68940 92520 69018 92576
rect 69074 92520 69708 92576
rect 69764 92520 69769 92576
rect 68940 92518 69769 92520
rect 68940 92516 68946 92518
rect 69013 92515 69079 92518
rect 69703 92515 69769 92518
rect 189073 92578 189139 92581
rect 190269 92578 190335 92581
rect 191097 92578 191163 92581
rect 189073 92576 191163 92578
rect 189073 92520 189078 92576
rect 189134 92520 190274 92576
rect 190330 92520 191102 92576
rect 191158 92520 191163 92576
rect 189073 92518 191163 92520
rect 189073 92515 189139 92518
rect 190269 92515 190335 92518
rect 191097 92515 191163 92518
rect 192334 92516 192340 92580
rect 192404 92578 192410 92580
rect 193121 92578 193187 92581
rect 192404 92576 193187 92578
rect 192404 92520 193126 92576
rect 193182 92520 193187 92576
rect 192404 92518 193187 92520
rect 192404 92516 192410 92518
rect 193121 92515 193187 92518
rect 71446 92380 71452 92444
rect 71516 92442 71522 92444
rect 73337 92442 73403 92445
rect 71516 92440 73403 92442
rect 71516 92384 73342 92440
rect 73398 92384 73403 92440
rect 71516 92382 73403 92384
rect 71516 92380 71522 92382
rect 73337 92379 73403 92382
rect 91001 92442 91067 92445
rect 91686 92442 91692 92444
rect 91001 92440 91692 92442
rect 91001 92384 91006 92440
rect 91062 92384 91692 92440
rect 91001 92382 91692 92384
rect 91001 92379 91067 92382
rect 91686 92380 91692 92382
rect 91756 92380 91762 92444
rect 91829 92442 91895 92445
rect 92974 92442 92980 92444
rect 91829 92440 92980 92442
rect 91829 92384 91834 92440
rect 91890 92384 92980 92440
rect 91829 92382 92980 92384
rect 91829 92379 91895 92382
rect 92974 92380 92980 92382
rect 93044 92380 93050 92444
rect 175181 92442 175247 92445
rect 196525 92442 196591 92445
rect 175181 92440 196591 92442
rect 175181 92384 175186 92440
rect 175242 92384 196530 92440
rect 196586 92384 196591 92440
rect 175181 92382 196591 92384
rect 175181 92379 175247 92382
rect 196525 92379 196591 92382
rect 197997 92442 198063 92445
rect 201534 92442 201540 92444
rect 197997 92440 201540 92442
rect 197997 92384 198002 92440
rect 198058 92384 201540 92440
rect 197997 92382 201540 92384
rect 197997 92379 198063 92382
rect 201534 92380 201540 92382
rect 201604 92380 201610 92444
rect 206093 92442 206159 92445
rect 211654 92442 211660 92444
rect 206093 92440 211660 92442
rect 206093 92384 206098 92440
rect 206154 92384 211660 92440
rect 206093 92382 211660 92384
rect 206093 92379 206159 92382
rect 211654 92380 211660 92382
rect 211724 92380 211730 92444
rect 61878 92244 61884 92308
rect 61948 92306 61954 92308
rect 61948 92246 64890 92306
rect 61948 92244 61954 92246
rect 64830 92170 64890 92246
rect 72918 92244 72924 92308
rect 72988 92306 72994 92308
rect 73705 92306 73771 92309
rect 92749 92306 92815 92309
rect 113173 92306 113239 92309
rect 72988 92304 84210 92306
rect 72988 92248 73710 92304
rect 73766 92248 84210 92304
rect 72988 92246 84210 92248
rect 72988 92244 72994 92246
rect 73705 92243 73771 92246
rect 74809 92170 74875 92173
rect 64830 92168 74875 92170
rect 64830 92112 74814 92168
rect 74870 92112 74875 92168
rect 64830 92110 74875 92112
rect 84150 92170 84210 92246
rect 92749 92304 113239 92306
rect 92749 92248 92754 92304
rect 92810 92248 113178 92304
rect 113234 92248 113239 92304
rect 92749 92246 113239 92248
rect 92749 92243 92815 92246
rect 113173 92243 113239 92246
rect 185669 92306 185735 92309
rect 224350 92306 224356 92308
rect 185669 92304 224356 92306
rect 185669 92248 185674 92304
rect 185730 92248 224356 92304
rect 185669 92246 224356 92248
rect 185669 92243 185735 92246
rect 224350 92244 224356 92246
rect 224420 92244 224426 92308
rect 158621 92170 158687 92173
rect 84150 92168 158687 92170
rect 84150 92112 158626 92168
rect 158682 92112 158687 92168
rect 84150 92110 158687 92112
rect 74809 92107 74875 92110
rect 158621 92107 158687 92110
rect 184841 92170 184907 92173
rect 200757 92170 200823 92173
rect 184841 92168 200823 92170
rect 184841 92112 184846 92168
rect 184902 92112 200762 92168
rect 200818 92112 200823 92168
rect 184841 92110 200823 92112
rect 184841 92107 184907 92110
rect 200757 92107 200823 92110
rect 205541 92170 205607 92173
rect 251766 92170 251772 92172
rect 205541 92168 251772 92170
rect 205541 92112 205546 92168
rect 205602 92112 251772 92168
rect 205541 92110 251772 92112
rect 205541 92107 205607 92110
rect 251766 92108 251772 92110
rect 251836 92108 251842 92172
rect 92381 92034 92447 92037
rect 94814 92034 94820 92036
rect 92381 92032 94820 92034
rect 92381 91976 92386 92032
rect 92442 91976 94820 92032
rect 92381 91974 94820 91976
rect 92381 91971 92447 91974
rect 94814 91972 94820 91974
rect 94884 91972 94890 92036
rect 251766 91700 251772 91764
rect 251836 91762 251842 91764
rect 334617 91762 334683 91765
rect 251836 91760 334683 91762
rect 251836 91704 334622 91760
rect 334678 91704 334683 91760
rect 251836 91702 334683 91704
rect 251836 91700 251842 91702
rect 334617 91699 334683 91702
rect 82629 91218 82695 91221
rect 83457 91218 83523 91221
rect 82629 91216 83523 91218
rect 82629 91160 82634 91216
rect 82690 91160 83462 91216
rect 83518 91160 83523 91216
rect 82629 91158 83523 91160
rect 82629 91155 82695 91158
rect 83457 91155 83523 91158
rect 200205 91082 200271 91085
rect 200941 91082 201007 91085
rect 219157 91084 219223 91085
rect 219157 91082 219204 91084
rect 74490 91080 201007 91082
rect 74490 91024 200210 91080
rect 200266 91024 200946 91080
rect 201002 91024 201007 91080
rect 74490 91022 201007 91024
rect 219076 91080 219204 91082
rect 219268 91082 219274 91084
rect 220077 91082 220143 91085
rect 219268 91080 220143 91082
rect 219076 91024 219162 91080
rect 219268 91024 220082 91080
rect 220138 91024 220143 91080
rect 219076 91022 219204 91024
rect 56409 90946 56475 90949
rect 74349 90946 74415 90949
rect 74490 90946 74550 91022
rect 200205 91019 200271 91022
rect 200941 91019 201007 91022
rect 219157 91020 219204 91022
rect 219268 91022 220143 91024
rect 219268 91020 219274 91022
rect 219157 91019 219223 91020
rect 220077 91019 220143 91022
rect 224309 91082 224375 91085
rect 258165 91082 258231 91085
rect 224309 91080 258231 91082
rect 224309 91024 224314 91080
rect 224370 91024 258170 91080
rect 258226 91024 258231 91080
rect 224309 91022 258231 91024
rect 224309 91019 224375 91022
rect 258165 91019 258231 91022
rect 56409 90944 74550 90946
rect 56409 90888 56414 90944
rect 56470 90888 74354 90944
rect 74410 90888 74550 90944
rect 56409 90886 74550 90888
rect 56409 90883 56475 90886
rect 74349 90883 74415 90886
rect 108389 90538 108455 90541
rect 203701 90538 203767 90541
rect 108389 90536 203767 90538
rect 108389 90480 108394 90536
rect 108450 90480 203706 90536
rect 203762 90480 203767 90536
rect 108389 90478 203767 90480
rect 108389 90475 108455 90478
rect 203701 90475 203767 90478
rect 107009 90402 107075 90405
rect 204437 90402 204503 90405
rect 107009 90400 204503 90402
rect 107009 90344 107014 90400
rect 107070 90344 204442 90400
rect 204498 90344 204503 90400
rect 107009 90342 204503 90344
rect 107009 90339 107075 90342
rect 204437 90339 204503 90342
rect 219433 90402 219499 90405
rect 239397 90402 239463 90405
rect 219433 90400 239463 90402
rect 219433 90344 219438 90400
rect 219494 90344 239402 90400
rect 239458 90344 239463 90400
rect 219433 90342 239463 90344
rect 219433 90339 219499 90342
rect 239397 90339 239463 90342
rect 205633 90268 205699 90269
rect 205582 90266 205588 90268
rect 205506 90206 205588 90266
rect 205652 90266 205699 90268
rect 206829 90266 206895 90269
rect 215293 90268 215359 90269
rect 215293 90266 215340 90268
rect 205652 90264 206895 90266
rect 205694 90208 206834 90264
rect 206890 90208 206895 90264
rect 205582 90204 205588 90206
rect 205652 90206 206895 90208
rect 215212 90264 215340 90266
rect 215404 90266 215410 90268
rect 216397 90266 216463 90269
rect 215404 90264 216463 90266
rect 215212 90208 215298 90264
rect 215404 90208 216402 90264
rect 216458 90208 216463 90264
rect 215212 90206 215340 90208
rect 205652 90204 205699 90206
rect 205633 90203 205699 90204
rect 206829 90203 206895 90206
rect 215293 90204 215340 90206
rect 215404 90206 216463 90208
rect 215404 90204 215410 90206
rect 215293 90203 215359 90204
rect 216397 90203 216463 90206
rect 94773 89858 94839 89861
rect 95182 89858 95188 89860
rect 94773 89856 95188 89858
rect 94773 89800 94778 89856
rect 94834 89800 95188 89856
rect 94773 89798 95188 89800
rect 94773 89795 94839 89798
rect 95182 89796 95188 89798
rect 95252 89796 95258 89860
rect 82997 89722 83063 89725
rect 186313 89722 186379 89725
rect 210325 89722 210391 89725
rect 82997 89720 210391 89722
rect 82997 89664 83002 89720
rect 83058 89664 186318 89720
rect 186374 89664 210330 89720
rect 210386 89664 210391 89720
rect 82997 89662 210391 89664
rect 82997 89659 83063 89662
rect 186313 89659 186379 89662
rect 210325 89659 210391 89662
rect 211613 89722 211679 89725
rect 260925 89722 260991 89725
rect 211613 89720 260991 89722
rect 211613 89664 211618 89720
rect 211674 89664 260930 89720
rect 260986 89664 260991 89720
rect 211613 89662 260991 89664
rect 211613 89659 211679 89662
rect 260925 89659 260991 89662
rect 70158 89524 70164 89588
rect 70228 89586 70234 89588
rect 84653 89586 84719 89589
rect 84837 89586 84903 89589
rect 70228 89584 84903 89586
rect 70228 89528 84658 89584
rect 84714 89528 84842 89584
rect 84898 89528 84903 89584
rect 70228 89526 84903 89528
rect 70228 89524 70234 89526
rect 84653 89523 84719 89526
rect 84837 89523 84903 89526
rect 87229 89586 87295 89589
rect 122925 89586 122991 89589
rect 215201 89586 215267 89589
rect 87229 89584 215267 89586
rect 87229 89528 87234 89584
rect 87290 89528 122930 89584
rect 122986 89528 215206 89584
rect 215262 89528 215267 89584
rect 87229 89526 215267 89528
rect 87229 89523 87295 89526
rect 122925 89523 122991 89526
rect 215201 89523 215267 89526
rect 219801 89586 219867 89589
rect 254577 89586 254643 89589
rect 219801 89584 254643 89586
rect 219801 89528 219806 89584
rect 219862 89528 254582 89584
rect 254638 89528 254643 89584
rect 219801 89526 254643 89528
rect 219801 89523 219867 89526
rect 254577 89523 254643 89526
rect 81525 89450 81591 89453
rect 95233 89450 95299 89453
rect 81525 89448 95299 89450
rect 81525 89392 81530 89448
rect 81586 89392 95238 89448
rect 95294 89392 95299 89448
rect 81525 89390 95299 89392
rect 81525 89387 81591 89390
rect 95233 89387 95299 89390
rect 189717 89450 189783 89453
rect 225045 89450 225111 89453
rect 189717 89448 225111 89450
rect 189717 89392 189722 89448
rect 189778 89392 225050 89448
rect 225106 89392 225111 89448
rect 189717 89390 225111 89392
rect 189717 89387 189783 89390
rect 225045 89387 225111 89390
rect 50981 88226 51047 88229
rect 71773 88226 71839 88229
rect 72601 88226 72667 88229
rect 50981 88224 72667 88226
rect 50981 88168 50986 88224
rect 51042 88168 71778 88224
rect 71834 88168 72606 88224
rect 72662 88168 72667 88224
rect 50981 88166 72667 88168
rect 50981 88163 51047 88166
rect 71773 88163 71839 88166
rect 72601 88163 72667 88166
rect 82077 88226 82143 88229
rect 115197 88226 115263 88229
rect 209221 88226 209287 88229
rect 82077 88224 209287 88226
rect 82077 88168 82082 88224
rect 82138 88168 115202 88224
rect 115258 88168 209226 88224
rect 209282 88168 209287 88224
rect 82077 88166 209287 88168
rect 82077 88163 82143 88166
rect 115197 88163 115263 88166
rect 209221 88163 209287 88166
rect 78029 88090 78095 88093
rect 107009 88090 107075 88093
rect 78029 88088 107075 88090
rect 78029 88032 78034 88088
rect 78090 88032 107014 88088
rect 107070 88032 107075 88088
rect 78029 88030 107075 88032
rect 78029 88027 78095 88030
rect 107009 88027 107075 88030
rect 203701 88090 203767 88093
rect 284385 88090 284451 88093
rect 203701 88088 287070 88090
rect 203701 88032 203706 88088
rect 203762 88032 284390 88088
rect 284446 88032 287070 88088
rect 203701 88030 287070 88032
rect 203701 88027 203767 88030
rect 284385 88027 284451 88030
rect 84101 87954 84167 87957
rect 98821 87954 98887 87957
rect 84101 87952 98887 87954
rect 84101 87896 84106 87952
rect 84162 87896 98826 87952
rect 98882 87896 98887 87952
rect 84101 87894 98887 87896
rect 84101 87891 84167 87894
rect 98821 87891 98887 87894
rect 187693 87954 187759 87957
rect 227662 87954 227668 87956
rect 187693 87952 227668 87954
rect 187693 87896 187698 87952
rect 187754 87896 227668 87952
rect 187693 87894 227668 87896
rect 187693 87891 187759 87894
rect 227662 87892 227668 87894
rect 227732 87892 227738 87956
rect 287010 87546 287070 88030
rect 582833 87546 582899 87549
rect 287010 87544 582899 87546
rect 287010 87488 582838 87544
rect 582894 87488 582899 87544
rect 287010 87486 582899 87488
rect 582833 87483 582899 87486
rect 72601 86866 72667 86869
rect 197077 86866 197143 86869
rect 72601 86864 197143 86866
rect 72601 86808 72606 86864
rect 72662 86808 197082 86864
rect 197138 86808 197143 86864
rect 72601 86806 197143 86808
rect 72601 86803 72667 86806
rect 197077 86803 197143 86806
rect 68553 86730 68619 86733
rect 102317 86730 102383 86733
rect 68553 86728 102383 86730
rect 68553 86672 68558 86728
rect 68614 86672 102322 86728
rect 102378 86672 102383 86728
rect 68553 86670 102383 86672
rect 68553 86667 68619 86670
rect 102317 86667 102383 86670
rect 189942 86668 189948 86732
rect 190012 86730 190018 86732
rect 226374 86730 226380 86732
rect 190012 86670 226380 86730
rect 190012 86668 190018 86670
rect 226374 86668 226380 86670
rect 226444 86668 226450 86732
rect 76373 86594 76439 86597
rect 95969 86594 96035 86597
rect 76373 86592 96035 86594
rect 76373 86536 76378 86592
rect 76434 86536 95974 86592
rect 96030 86536 96035 86592
rect 76373 86534 96035 86536
rect 76373 86531 76439 86534
rect 95969 86531 96035 86534
rect 192702 86124 192708 86188
rect 192772 86186 192778 86188
rect 273253 86186 273319 86189
rect 192772 86184 273319 86186
rect 192772 86128 273258 86184
rect 273314 86128 273319 86184
rect 192772 86126 273319 86128
rect 192772 86124 192778 86126
rect 273253 86123 273319 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 64689 85506 64755 85509
rect 193806 85506 193812 85508
rect 64689 85504 193812 85506
rect 64689 85448 64694 85504
rect 64750 85448 193812 85504
rect 64689 85446 193812 85448
rect 64689 85443 64755 85446
rect 193806 85444 193812 85446
rect 193876 85506 193882 85508
rect 194542 85506 194548 85508
rect 193876 85446 194548 85506
rect 193876 85444 193882 85446
rect 194542 85444 194548 85446
rect 194612 85444 194618 85508
rect 91277 85370 91343 85373
rect 219157 85370 219223 85373
rect 91277 85368 219223 85370
rect 91277 85312 91282 85368
rect 91338 85312 219162 85368
rect 219218 85312 219223 85368
rect 91277 85310 219223 85312
rect 91277 85307 91343 85310
rect 219157 85307 219223 85310
rect 66478 85172 66484 85236
rect 66548 85234 66554 85236
rect 101397 85234 101463 85237
rect 66548 85232 101463 85234
rect 66548 85176 101402 85232
rect 101458 85176 101463 85232
rect 66548 85174 101463 85176
rect 66548 85172 66554 85174
rect 101397 85171 101463 85174
rect -960 84690 480 84780
rect 194542 84764 194548 84828
rect 194612 84826 194618 84828
rect 310513 84826 310579 84829
rect 194612 84824 310579 84826
rect 194612 84768 310518 84824
rect 310574 84768 310579 84824
rect 194612 84766 310579 84768
rect 194612 84764 194618 84766
rect 310513 84763 310579 84766
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 98913 84146 98979 84149
rect 226701 84146 226767 84149
rect 98913 84144 226767 84146
rect 98913 84088 98918 84144
rect 98974 84088 226706 84144
rect 226762 84088 226767 84144
rect 98913 84086 226767 84088
rect 98913 84083 98979 84086
rect 226701 84083 226767 84086
rect 69606 83948 69612 84012
rect 69676 84010 69682 84012
rect 120717 84010 120783 84013
rect 69676 84008 120783 84010
rect 69676 83952 120722 84008
rect 120778 83952 120783 84008
rect 69676 83950 120783 83952
rect 69676 83948 69682 83950
rect 120717 83947 120783 83950
rect 90357 83466 90423 83469
rect 96613 83466 96679 83469
rect 90357 83464 96679 83466
rect 90357 83408 90362 83464
rect 90418 83408 96618 83464
rect 96674 83408 96679 83464
rect 90357 83406 96679 83408
rect 90357 83403 90423 83406
rect 96613 83403 96679 83406
rect 89897 82786 89963 82789
rect 220077 82786 220143 82789
rect 89897 82784 220143 82786
rect 89897 82728 89902 82784
rect 89958 82728 220082 82784
rect 220138 82728 220143 82784
rect 89897 82726 220143 82728
rect 89897 82723 89963 82726
rect 220077 82723 220143 82726
rect 69013 82106 69079 82109
rect 181437 82106 181503 82109
rect 69013 82104 181503 82106
rect 69013 82048 69018 82104
rect 69074 82048 181442 82104
rect 181498 82048 181503 82104
rect 69013 82046 181503 82048
rect 69013 82043 69079 82046
rect 181437 82043 181503 82046
rect 195094 82044 195100 82108
rect 195164 82106 195170 82108
rect 291837 82106 291903 82109
rect 195164 82104 291903 82106
rect 195164 82048 291842 82104
rect 291898 82048 291903 82104
rect 195164 82046 291903 82048
rect 195164 82044 195170 82046
rect 291837 82043 291903 82046
rect 178033 81426 178099 81429
rect 179321 81426 179387 81429
rect 209865 81426 209931 81429
rect 211061 81426 211127 81429
rect 178033 81424 211127 81426
rect 178033 81368 178038 81424
rect 178094 81368 179326 81424
rect 179382 81368 209870 81424
rect 209926 81368 211066 81424
rect 211122 81368 211127 81424
rect 178033 81366 211127 81368
rect 178033 81363 178099 81366
rect 179321 81363 179387 81366
rect 209865 81363 209931 81366
rect 211061 81363 211127 81366
rect 56593 80746 56659 80749
rect 180057 80746 180123 80749
rect 56593 80744 180123 80746
rect 56593 80688 56598 80744
rect 56654 80688 180062 80744
rect 180118 80688 180123 80744
rect 56593 80686 180123 80688
rect 56593 80683 56659 80686
rect 180057 80683 180123 80686
rect 211061 80746 211127 80749
rect 582925 80746 582991 80749
rect 211061 80744 582991 80746
rect 211061 80688 211066 80744
rect 211122 80688 582930 80744
rect 582986 80688 582991 80744
rect 211061 80686 582991 80688
rect 211061 80683 211127 80686
rect 582925 80683 582991 80686
rect 79317 79386 79383 79389
rect 126329 79386 126395 79389
rect 79317 79384 126395 79386
rect 79317 79328 79322 79384
rect 79378 79328 126334 79384
rect 126390 79328 126395 79384
rect 79317 79326 126395 79328
rect 79317 79323 79383 79326
rect 126329 79323 126395 79326
rect 196566 79324 196572 79388
rect 196636 79386 196642 79388
rect 262213 79386 262279 79389
rect 196636 79384 262279 79386
rect 196636 79328 262218 79384
rect 262274 79328 262279 79384
rect 196636 79326 262279 79328
rect 196636 79324 196642 79326
rect 262213 79323 262279 79326
rect 66161 78570 66227 78573
rect 188429 78570 188495 78573
rect 66161 78568 188495 78570
rect 66161 78512 66166 78568
rect 66222 78512 188434 78568
rect 188490 78512 188495 78568
rect 66161 78510 188495 78512
rect 66161 78507 66227 78510
rect 188429 78507 188495 78510
rect 202873 77890 202939 77893
rect 203517 77890 203583 77893
rect 231853 77890 231919 77893
rect 232589 77890 232655 77893
rect 202873 77888 232655 77890
rect 202873 77832 202878 77888
rect 202934 77832 203522 77888
rect 203578 77832 231858 77888
rect 231914 77832 232594 77888
rect 232650 77832 232655 77888
rect 202873 77830 232655 77832
rect 202873 77827 202939 77830
rect 203517 77827 203583 77830
rect 231853 77827 231919 77830
rect 232589 77827 232655 77830
rect 95141 77210 95207 77213
rect 203517 77210 203583 77213
rect 95141 77208 203583 77210
rect 95141 77152 95146 77208
rect 95202 77152 203522 77208
rect 203578 77152 203583 77208
rect 95141 77150 203583 77152
rect 95141 77147 95207 77150
rect 203517 77147 203583 77150
rect 97206 75788 97212 75852
rect 97276 75850 97282 75852
rect 227989 75850 228055 75853
rect 97276 75848 228055 75850
rect 97276 75792 227994 75848
rect 228050 75792 228055 75848
rect 97276 75790 228055 75792
rect 97276 75788 97282 75790
rect 227989 75787 228055 75790
rect 70393 73810 70459 73813
rect 173157 73810 173223 73813
rect 70393 73808 173223 73810
rect 70393 73752 70398 73808
rect 70454 73752 173162 73808
rect 173218 73752 173223 73808
rect 70393 73750 173223 73752
rect 70393 73747 70459 73750
rect 173157 73747 173223 73750
rect 193213 73810 193279 73813
rect 269113 73810 269179 73813
rect 193213 73808 269179 73810
rect 193213 73752 193218 73808
rect 193274 73752 269118 73808
rect 269174 73752 269179 73808
rect 193213 73750 269179 73752
rect 193213 73747 193279 73750
rect 269113 73747 269179 73750
rect 188337 73130 188403 73133
rect 231117 73130 231183 73133
rect 188337 73128 231183 73130
rect 188337 73072 188342 73128
rect 188398 73072 231122 73128
rect 231178 73072 231183 73128
rect 188337 73070 231183 73072
rect 188337 73067 188403 73070
rect 231117 73067 231183 73070
rect 583017 72994 583083 72997
rect 583520 72994 584960 73084
rect 583017 72992 584960 72994
rect 583017 72936 583022 72992
rect 583078 72936 584960 72992
rect 583017 72934 584960 72936
rect 583017 72931 583083 72934
rect 583520 72844 584960 72934
rect 74533 72450 74599 72453
rect 168230 72450 168236 72452
rect 74533 72448 168236 72450
rect 74533 72392 74538 72448
rect 74594 72392 168236 72448
rect 74533 72390 168236 72392
rect 74533 72387 74599 72390
rect 168230 72388 168236 72390
rect 168300 72388 168306 72452
rect 106273 71770 106339 71773
rect 212533 71770 212599 71773
rect 106273 71768 212599 71770
rect -960 71634 480 71724
rect 106273 71712 106278 71768
rect 106334 71712 212538 71768
rect 212594 71712 212599 71768
rect 106273 71710 212599 71712
rect 106273 71707 106339 71710
rect 212533 71707 212599 71710
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 92473 71090 92539 71093
rect 163589 71090 163655 71093
rect 92473 71088 163655 71090
rect 92473 71032 92478 71088
rect 92534 71032 163594 71088
rect 163650 71032 163655 71088
rect 92473 71030 163655 71032
rect 92473 71027 92539 71030
rect 163589 71027 163655 71030
rect 212533 70410 212599 70413
rect 213177 70410 213243 70413
rect 212533 70408 213243 70410
rect 212533 70352 212538 70408
rect 212594 70352 213182 70408
rect 213238 70352 213243 70408
rect 212533 70350 213243 70352
rect 212533 70347 212599 70350
rect 213177 70347 213243 70350
rect 59261 70274 59327 70277
rect 186957 70274 187023 70277
rect 59261 70272 187023 70274
rect 59261 70216 59266 70272
rect 59322 70216 186962 70272
rect 187018 70216 187023 70272
rect 59261 70214 187023 70216
rect 59261 70211 59327 70214
rect 186957 70211 187023 70214
rect 93853 68234 93919 68237
rect 127617 68234 127683 68237
rect 93853 68232 127683 68234
rect 93853 68176 93858 68232
rect 93914 68176 127622 68232
rect 127678 68176 127683 68232
rect 93853 68174 127683 68176
rect 93853 68171 93919 68174
rect 127617 68171 127683 68174
rect 94497 67554 94563 67557
rect 222285 67554 222351 67557
rect 94497 67552 222351 67554
rect 94497 67496 94502 67552
rect 94558 67496 222290 67552
rect 222346 67496 222351 67552
rect 94497 67494 222351 67496
rect 94497 67491 94563 67494
rect 222285 67491 222351 67494
rect 582741 59666 582807 59669
rect 583520 59666 584960 59756
rect 582741 59664 584960 59666
rect 582741 59608 582746 59664
rect 582802 59608 584960 59664
rect 582741 59606 584960 59608
rect 582741 59603 582807 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 66253 55858 66319 55861
rect 105486 55858 105492 55860
rect 66253 55856 105492 55858
rect 66253 55800 66258 55856
rect 66314 55800 105492 55856
rect 66253 55798 105492 55800
rect 66253 55795 66319 55798
rect 105486 55796 105492 55798
rect 105556 55796 105562 55860
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 53833 44842 53899 44845
rect 141366 44842 141372 44844
rect 53833 44840 141372 44842
rect 53833 44784 53838 44840
rect 53894 44784 141372 44840
rect 53833 44782 141372 44784
rect 53833 44779 53899 44782
rect 141366 44780 141372 44782
rect 141436 44780 141442 44844
rect 46933 43482 46999 43485
rect 144126 43482 144132 43484
rect 46933 43480 144132 43482
rect 46933 43424 46938 43480
rect 46994 43424 144132 43480
rect 46933 43422 144132 43424
rect 46933 43419 46999 43422
rect 144126 43420 144132 43422
rect 144196 43420 144202 43484
rect 203190 40564 203196 40628
rect 203260 40626 203266 40628
rect 306373 40626 306439 40629
rect 203260 40624 306439 40626
rect 203260 40568 306378 40624
rect 306434 40568 306439 40624
rect 203260 40566 306439 40568
rect 203260 40564 203266 40566
rect 306373 40563 306439 40566
rect 582925 33146 582991 33149
rect 583520 33146 584960 33236
rect 582925 33144 584960 33146
rect 582925 33088 582930 33144
rect 582986 33088 584960 33144
rect 582925 33086 584960 33088
rect 582925 33083 582991 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 35893 30970 35959 30973
rect 166206 30970 166212 30972
rect 35893 30968 166212 30970
rect 35893 30912 35898 30968
rect 35954 30912 166212 30968
rect 35893 30910 166212 30912
rect 35893 30907 35959 30910
rect 166206 30908 166212 30910
rect 166276 30908 166282 30972
rect 55213 28250 55279 28253
rect 106774 28250 106780 28252
rect 55213 28248 106780 28250
rect 55213 28192 55218 28248
rect 55274 28192 106780 28248
rect 55213 28190 106780 28192
rect 55213 28187 55279 28190
rect 106774 28188 106780 28190
rect 106844 28188 106850 28252
rect 85665 26890 85731 26893
rect 175774 26890 175780 26892
rect 85665 26888 175780 26890
rect 85665 26832 85670 26888
rect 85726 26832 175780 26888
rect 85665 26830 175780 26832
rect 85665 26827 85731 26830
rect 175774 26828 175780 26830
rect 175844 26828 175850 26892
rect 582649 19818 582715 19821
rect 583520 19818 584960 19908
rect 582649 19816 584960 19818
rect 582649 19760 582654 19816
rect 582710 19760 584960 19816
rect 582649 19758 584960 19760
rect 582649 19755 582715 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 98177 15874 98243 15877
rect 124806 15874 124812 15876
rect 98177 15872 124812 15874
rect 98177 15816 98182 15872
rect 98238 15816 124812 15872
rect 98177 15814 124812 15816
rect 98177 15811 98243 15814
rect 124806 15812 124812 15814
rect 124876 15812 124882 15876
rect 582833 6626 582899 6629
rect 583520 6626 584960 6716
rect 582833 6624 584960 6626
rect -960 6490 480 6580
rect 582833 6568 582838 6624
rect 582894 6568 584960 6624
rect 582833 6566 584960 6568
rect 582833 6563 582899 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 26509 6218 26575 6221
rect 186814 6218 186820 6220
rect 26509 6216 186820 6218
rect 26509 6160 26514 6216
rect 26570 6160 186820 6216
rect 26509 6158 186820 6160
rect 26509 6155 26575 6158
rect 186814 6156 186820 6158
rect 186884 6156 186890 6220
rect 224861 4858 224927 4861
rect 254669 4858 254735 4861
rect 224861 4856 254735 4858
rect 224861 4800 224866 4856
rect 224922 4800 254674 4856
rect 254730 4800 254735 4856
rect 224861 4798 254735 4800
rect 224861 4795 224927 4798
rect 254669 4795 254735 4798
rect 226977 3362 227043 3365
rect 265341 3362 265407 3365
rect 226977 3360 265407 3362
rect 226977 3304 226982 3360
rect 227038 3304 265346 3360
rect 265402 3304 265407 3360
rect 226977 3302 265407 3304
rect 226977 3299 227043 3302
rect 265341 3299 265407 3302
rect 291837 3362 291903 3365
rect 301957 3362 302023 3365
rect 291837 3360 302023 3362
rect 291837 3304 291842 3360
rect 291898 3304 301962 3360
rect 302018 3304 302023 3360
rect 291837 3302 302023 3304
rect 291837 3299 291903 3302
rect 301957 3299 302023 3302
<< via3 >>
rect 72924 699816 72988 699820
rect 72924 699760 72974 699816
rect 72974 699760 72988 699816
rect 72924 699756 72988 699760
rect 162716 619652 162780 619716
rect 180012 609996 180076 610060
rect 184060 608772 184124 608836
rect 192340 607276 192404 607340
rect 258396 603060 258460 603124
rect 244596 601836 244660 601900
rect 259500 601700 259564 601764
rect 154436 600884 154500 600948
rect 219940 600748 220004 600812
rect 232452 600612 232516 600676
rect 193444 600476 193508 600540
rect 263548 600476 263612 600540
rect 215340 600400 215404 600404
rect 215340 600344 215354 600400
rect 215354 600344 215404 600400
rect 215340 600340 215404 600344
rect 218652 600340 218716 600404
rect 230980 600340 231044 600404
rect 276244 600340 276308 600404
rect 212396 599448 212460 599452
rect 212396 599392 212446 599448
rect 212446 599392 212460 599448
rect 212396 599388 212460 599392
rect 226380 599448 226444 599452
rect 226380 599392 226394 599448
rect 226394 599392 226444 599448
rect 226380 599388 226444 599392
rect 238524 599388 238588 599452
rect 204852 599116 204916 599180
rect 222700 599116 222764 599180
rect 229692 599116 229756 599180
rect 237420 599116 237484 599180
rect 241652 599116 241716 599180
rect 262260 599116 262324 599180
rect 194548 599040 194612 599044
rect 194548 598984 194598 599040
rect 194598 598984 194612 599040
rect 194548 598980 194612 598984
rect 197124 599040 197188 599044
rect 197124 598984 197174 599040
rect 197174 598984 197188 599040
rect 197124 598980 197188 598984
rect 201540 599040 201604 599044
rect 201540 598984 201590 599040
rect 201590 598984 201604 599040
rect 201540 598980 201604 598984
rect 203012 599040 203076 599044
rect 203012 598984 203062 599040
rect 203062 598984 203076 599040
rect 203012 598980 203076 598984
rect 207060 599040 207124 599044
rect 207060 598984 207110 599040
rect 207110 598984 207124 599040
rect 207060 598980 207124 598984
rect 210740 599040 210804 599044
rect 210740 598984 210790 599040
rect 210790 598984 210804 599040
rect 210740 598980 210804 598984
rect 219572 598980 219636 599044
rect 220860 599040 220924 599044
rect 220860 598984 220910 599040
rect 220910 598984 220924 599040
rect 220860 598980 220924 598984
rect 223804 599040 223868 599044
rect 223804 598984 223854 599040
rect 223854 598984 223868 599040
rect 223804 598980 223868 598984
rect 223988 598980 224052 599044
rect 228220 598980 228284 599044
rect 230612 599040 230676 599044
rect 230612 598984 230662 599040
rect 230662 598984 230676 599040
rect 230612 598980 230676 598984
rect 233188 599040 233252 599044
rect 233188 598984 233238 599040
rect 233238 598984 233252 599040
rect 233188 598980 233252 598984
rect 234660 599040 234724 599044
rect 234660 598984 234710 599040
rect 234710 598984 234724 599040
rect 234660 598980 234724 598984
rect 236500 598980 236564 599044
rect 240732 599040 240796 599044
rect 240732 598984 240746 599040
rect 240746 598984 240796 599040
rect 240732 598980 240796 598984
rect 242940 598980 243004 599044
rect 247724 599040 247788 599044
rect 247724 598984 247774 599040
rect 247774 598984 247788 599040
rect 247724 598980 247788 598984
rect 249932 598980 249996 599044
rect 252508 598980 252572 599044
rect 193260 598436 193324 598500
rect 192340 598164 192404 598228
rect 193444 596804 193508 596868
rect 188292 596320 188356 596324
rect 188292 596264 188306 596320
rect 188306 596264 188356 596320
rect 188292 596260 188356 596264
rect 270540 596260 270604 596324
rect 193260 595444 193324 595508
rect 258396 594764 258460 594828
rect 269068 592588 269132 592652
rect 267780 590684 267844 590748
rect 193812 590140 193876 590204
rect 281580 589868 281644 589932
rect 159772 587964 159836 588028
rect 265756 587148 265820 587212
rect 266308 586468 266372 586532
rect 75684 580892 75748 580956
rect 70900 580816 70964 580820
rect 70900 580760 70950 580816
rect 70950 580760 70964 580816
rect 70900 580756 70964 580760
rect 79916 580816 79980 580820
rect 79916 580760 79966 580816
rect 79966 580760 79980 580816
rect 79916 580756 79980 580760
rect 84700 580816 84764 580820
rect 84700 580760 84714 580816
rect 84714 580760 84764 580816
rect 84700 580756 84764 580760
rect 89300 580816 89364 580820
rect 89300 580760 89314 580816
rect 89314 580760 89364 580816
rect 89300 580756 89364 580760
rect 66668 578580 66732 578644
rect 156644 578852 156708 578916
rect 178540 572732 178604 572796
rect 255268 570556 255332 570620
rect 172100 568652 172164 568716
rect 166764 565796 166828 565860
rect 260972 563348 261036 563412
rect 263732 563076 263796 563140
rect 67772 561988 67836 562052
rect 170812 560356 170876 560420
rect 186820 558180 186884 558244
rect 148180 554780 148244 554844
rect 96660 553420 96724 553484
rect 158484 552196 158548 552260
rect 104940 551924 105004 551988
rect 253980 551720 254044 551784
rect 69428 551108 69492 551172
rect 96660 551244 96724 551308
rect 69428 549476 69492 549540
rect 101260 549340 101324 549404
rect 96844 547028 96908 547092
rect 67956 543356 68020 543420
rect 188476 542404 188540 542468
rect 72924 539548 72988 539612
rect 161244 539548 161308 539612
rect 69612 539064 69676 539068
rect 69612 539008 69662 539064
rect 69662 539008 69676 539064
rect 69612 539004 69676 539008
rect 255268 539276 255332 539340
rect 251220 539004 251284 539068
rect 253980 537372 254044 537436
rect 69612 536208 69676 536212
rect 69612 536152 69662 536208
rect 69662 536152 69676 536208
rect 69612 536148 69676 536152
rect 88196 535468 88260 535532
rect 196020 535468 196084 535532
rect 238524 531932 238588 531996
rect 218652 530708 218716 530772
rect 230612 530708 230676 530772
rect 69796 530572 69860 530636
rect 82860 530572 82924 530636
rect 111748 530572 111812 530636
rect 96660 529212 96724 529276
rect 248460 528532 248524 528596
rect 66116 526356 66180 526420
rect 219940 526356 220004 526420
rect 159956 523636 160020 523700
rect 249748 523636 249812 523700
rect 219572 522412 219636 522476
rect 229692 522276 229756 522340
rect 67956 521596 68020 521660
rect 68876 521596 68940 521660
rect 77156 520916 77220 520980
rect 96844 519420 96908 519484
rect 232452 518876 232516 518940
rect 69612 516700 69676 516764
rect 184060 515340 184124 515404
rect 244412 515340 244476 515404
rect 72740 512620 72804 512684
rect 166212 512620 166276 512684
rect 211660 511396 211724 511460
rect 230980 511396 231044 511460
rect 245700 511396 245764 511460
rect 210740 511260 210804 511324
rect 226380 509764 226444 509828
rect 253060 509764 253124 509828
rect 222700 505684 222764 505748
rect 150940 502964 151004 503028
rect 75684 500108 75748 500172
rect 188476 498748 188540 498812
rect 204852 498748 204916 498812
rect 161060 497388 161124 497452
rect 244596 496572 244660 496636
rect 223804 489908 223868 489972
rect 251220 489092 251284 489156
rect 168972 486508 169036 486572
rect 197124 486372 197188 486436
rect 254532 486372 254596 486436
rect 252508 484392 252572 484396
rect 252508 484336 252558 484392
rect 252558 484336 252572 484392
rect 252508 484332 252572 484336
rect 252692 483788 252756 483852
rect 237420 483652 237484 483716
rect 89300 482836 89364 482900
rect 220860 482156 220924 482220
rect 249932 481748 249996 481812
rect 285628 481612 285692 481676
rect 240732 481536 240796 481540
rect 240732 481480 240782 481536
rect 240782 481480 240796 481536
rect 240732 481476 240796 481480
rect 262444 478076 262508 478140
rect 178724 476716 178788 476780
rect 249380 476172 249444 476236
rect 187556 475356 187620 475420
rect 186820 474132 186884 474196
rect 181484 471820 181548 471884
rect 173572 471276 173636 471340
rect 173756 469236 173820 469300
rect 180012 469236 180076 469300
rect 162532 468420 162596 468484
rect 68876 467936 68940 467940
rect 68876 467880 68926 467936
rect 68926 467880 68940 467936
rect 68876 467876 68940 467880
rect 190316 467060 190380 467124
rect 203012 467060 203076 467124
rect 66116 466516 66180 466580
rect 255268 466516 255332 466580
rect 170996 465836 171060 465900
rect 201540 465836 201604 465900
rect 236500 465836 236564 465900
rect 67772 465700 67836 465764
rect 91324 465700 91388 465764
rect 223988 465700 224052 465764
rect 215340 464476 215404 464540
rect 176516 464340 176580 464404
rect 223804 464340 223868 464404
rect 104204 462844 104268 462908
rect 177620 462844 177684 462908
rect 207060 462844 207124 462908
rect 188844 459036 188908 459100
rect 233188 459036 233252 459100
rect 234660 458900 234724 458964
rect 184796 458764 184860 458828
rect 114324 457404 114388 457468
rect 180564 456316 180628 456380
rect 228220 456180 228284 456244
rect 247724 456044 247788 456108
rect 250300 455364 250364 455428
rect 112300 454684 112364 454748
rect 284340 454004 284404 454068
rect 173572 453868 173636 453932
rect 173572 453732 173636 453796
rect 273300 452432 273364 452436
rect 273300 452376 273314 452432
rect 273314 452376 273364 452432
rect 273300 452372 273364 452376
rect 247172 450604 247236 450668
rect 193076 450332 193140 450396
rect 177804 449380 177868 449444
rect 245700 449984 245764 449988
rect 245700 449928 245750 449984
rect 245750 449928 245764 449984
rect 245700 449924 245764 449928
rect 247724 449652 247788 449716
rect 253980 448760 254044 448764
rect 253980 448704 253994 448760
rect 253994 448704 254044 448760
rect 253980 448700 254044 448704
rect 70900 448624 70964 448628
rect 70900 448568 70914 448624
rect 70914 448568 70964 448624
rect 70900 448564 70964 448568
rect 254532 448564 254596 448628
rect 191788 448428 191852 448492
rect 69612 447748 69676 447812
rect 253060 446796 253124 446860
rect 193076 446524 193140 446588
rect 176516 444212 176580 444276
rect 176332 443532 176396 443596
rect 277348 441628 277412 441692
rect 252876 440948 252940 441012
rect 163452 438092 163516 438156
rect 255268 437548 255332 437612
rect 73476 436460 73540 436524
rect 79180 436324 79244 436388
rect 75132 436188 75196 436252
rect 81020 436188 81084 436252
rect 71084 436052 71148 436116
rect 94452 436052 94516 436116
rect 106044 436052 106108 436116
rect 102732 434556 102796 434620
rect 69244 434344 69308 434348
rect 69244 434288 69294 434344
rect 69294 434288 69308 434344
rect 69244 434284 69308 434288
rect 95188 434284 95252 434348
rect 100156 434344 100220 434348
rect 100156 434288 100206 434344
rect 100206 434288 100220 434344
rect 100156 434284 100220 434288
rect 92796 434208 92860 434212
rect 92796 434152 92810 434208
rect 92810 434152 92860 434208
rect 92796 434148 92860 434152
rect 80652 434012 80716 434076
rect 67956 433876 68020 433940
rect 78444 433740 78508 433804
rect 86724 433740 86788 433804
rect 98500 433740 98564 433804
rect 74764 433664 74828 433668
rect 74764 433608 74814 433664
rect 74814 433608 74828 433664
rect 74764 433604 74828 433608
rect 75868 433604 75932 433668
rect 78260 433604 78324 433668
rect 81940 433664 82004 433668
rect 81940 433608 81954 433664
rect 81954 433608 82004 433664
rect 81940 433604 82004 433608
rect 82492 433604 82556 433668
rect 83044 433604 83108 433668
rect 84516 433664 84580 433668
rect 84516 433608 84566 433664
rect 84566 433608 84580 433664
rect 84516 433604 84580 433608
rect 85804 433604 85868 433668
rect 87092 433604 87156 433668
rect 89668 433604 89732 433668
rect 90220 433604 90284 433668
rect 91508 433664 91572 433668
rect 91508 433608 91558 433664
rect 91558 433608 91572 433664
rect 91508 433604 91572 433608
rect 92980 433664 93044 433668
rect 92980 433608 93030 433664
rect 93030 433608 93044 433664
rect 92980 433604 93044 433608
rect 97948 433604 98012 433668
rect 99972 433604 100036 433668
rect 100708 433664 100772 433668
rect 100708 433608 100722 433664
rect 100722 433608 100772 433664
rect 100708 433604 100772 433608
rect 106412 433604 106476 433668
rect 109540 433664 109604 433668
rect 109540 433608 109554 433664
rect 109554 433608 109604 433664
rect 109540 433604 109604 433608
rect 111012 433604 111076 433668
rect 148180 433196 148244 433260
rect 69428 433060 69492 433124
rect 253060 430884 253124 430948
rect 253980 430884 254044 430948
rect 148180 429252 148244 429316
rect 113220 428164 113284 428228
rect 114508 427076 114572 427140
rect 170812 427076 170876 427140
rect 172100 423676 172164 423740
rect 66116 423268 66180 423332
rect 67956 422180 68020 422244
rect 155724 419596 155788 419660
rect 172284 419596 172348 419660
rect 287100 418236 287164 418300
rect 188292 417420 188356 417484
rect 280292 416740 280356 416804
rect 254532 415108 254596 415172
rect 150940 413884 151004 413948
rect 181484 406268 181548 406332
rect 191972 406268 192036 406332
rect 66668 402596 66732 402660
rect 112116 402596 112180 402660
rect 254716 402596 254780 402660
rect 162716 401644 162780 401708
rect 162716 401508 162780 401572
rect 113036 400148 113100 400212
rect 184796 397972 184860 398036
rect 66300 397292 66364 397356
rect 114324 396340 114388 396404
rect 252876 396748 252940 396812
rect 276428 395252 276492 395316
rect 112852 393892 112916 393956
rect 180748 393348 180812 393412
rect 180748 393136 180812 393140
rect 180748 393080 180762 393136
rect 180762 393080 180812 393136
rect 180748 393076 180812 393080
rect 254716 391988 254780 392052
rect 111932 391580 111996 391644
rect 113036 391580 113100 391644
rect 72740 390900 72804 390964
rect 84516 390900 84580 390964
rect 100156 390900 100220 390964
rect 104204 390960 104268 390964
rect 104204 390904 104254 390960
rect 104254 390904 104268 390960
rect 104204 390900 104268 390904
rect 104940 390900 105004 390964
rect 114508 391444 114572 391508
rect 111932 390960 111996 390964
rect 111932 390904 111982 390960
rect 111982 390904 111996 390960
rect 111932 390900 111996 390904
rect 79916 390764 79980 390828
rect 82860 390764 82924 390828
rect 191972 390688 192036 390692
rect 191972 390632 192022 390688
rect 192022 390632 192036 390688
rect 191972 390628 192036 390632
rect 84700 390492 84764 390556
rect 112852 390492 112916 390556
rect 77156 390416 77220 390420
rect 77156 390360 77206 390416
rect 77206 390360 77220 390416
rect 77156 390356 77220 390360
rect 91324 390356 91388 390420
rect 96660 390356 96724 390420
rect 190316 389812 190380 389876
rect 88196 389268 88260 389332
rect 249748 389268 249812 389332
rect 251036 389268 251100 389332
rect 244228 388996 244292 389060
rect 248644 389056 248708 389060
rect 248644 389000 248658 389056
rect 248658 389000 248708 389056
rect 248644 388996 248708 389000
rect 249380 388996 249444 389060
rect 72740 388860 72804 388924
rect 169708 388724 169772 388788
rect 101260 388588 101324 388652
rect 78260 388452 78324 388516
rect 80652 388452 80716 388516
rect 82492 388452 82556 388516
rect 247172 388512 247236 388516
rect 247172 388456 247222 388512
rect 247222 388456 247236 388512
rect 247172 388452 247236 388456
rect 83964 388316 84028 388380
rect 96660 387772 96724 387836
rect 75132 387636 75196 387700
rect 89668 387228 89732 387292
rect 247724 386956 247788 387020
rect 169708 386276 169772 386340
rect 170812 386276 170876 386340
rect 100708 385732 100772 385796
rect 74764 385052 74828 385116
rect 180748 383828 180812 383892
rect 180932 383556 180996 383620
rect 102732 382876 102796 382940
rect 242940 382876 243004 382940
rect 265940 382332 266004 382396
rect 258396 381652 258460 381716
rect 265756 381516 265820 381580
rect 276428 379340 276492 379404
rect 254532 378660 254596 378724
rect 287100 377980 287164 378044
rect 258396 377300 258460 377364
rect 267964 376620 268028 376684
rect 270540 375940 270604 376004
rect 188844 375396 188908 375460
rect 180748 374096 180812 374100
rect 180748 374040 180762 374096
rect 180762 374040 180812 374096
rect 180748 374036 180812 374040
rect 180748 373764 180812 373828
rect 241652 373356 241716 373420
rect 260972 373220 261036 373284
rect 187556 372676 187620 372740
rect 161060 371860 161124 371924
rect 262260 371860 262324 371924
rect 111012 370636 111076 370700
rect 92796 370500 92860 370564
rect 248460 370500 248524 370564
rect 280292 369744 280356 369748
rect 280292 369688 280306 369744
rect 280306 369688 280356 369744
rect 280292 369684 280356 369688
rect 70900 369004 70964 369068
rect 248644 369004 248708 369068
rect 180748 364440 180812 364444
rect 180748 364384 180762 364440
rect 180762 364384 180812 364440
rect 180748 364380 180812 364384
rect 180748 364108 180812 364172
rect 263732 362204 263796 362268
rect 266860 361660 266924 361724
rect 273484 360844 273548 360908
rect 271092 360164 271156 360228
rect 252508 360028 252572 360092
rect 273300 359348 273364 359412
rect 68876 357308 68940 357372
rect 269068 356628 269132 356692
rect 180748 354920 180812 354924
rect 180748 354864 180762 354920
rect 180762 354864 180812 354920
rect 180748 354860 180812 354864
rect 180748 354588 180812 354652
rect 259500 352548 259564 352612
rect 266308 351052 266372 351116
rect 159772 349828 159836 349892
rect 262260 349828 262324 349892
rect 124812 349692 124876 349756
rect 277532 349692 277596 349756
rect 262444 348468 262508 348532
rect 166764 346428 166828 346492
rect 253060 346292 253124 346356
rect 244228 344252 244292 344316
rect 177620 340912 177684 340916
rect 177620 340856 177634 340912
rect 177634 340856 177684 340912
rect 177620 340852 177684 340856
rect 177620 340172 177684 340236
rect 245700 339764 245764 339828
rect 81940 339492 82004 339556
rect 263548 338676 263612 338740
rect 158484 337996 158548 338060
rect 177988 337920 178052 337924
rect 177988 337864 178038 337920
rect 178038 337864 178052 337920
rect 177988 337860 178052 337864
rect 178724 337180 178788 337244
rect 144132 336772 144196 336836
rect 172284 334732 172348 334796
rect 178540 334656 178604 334660
rect 178540 334600 178590 334656
rect 178590 334600 178604 334656
rect 178540 334596 178604 334600
rect 263548 334596 263612 334660
rect 168972 333296 169036 333300
rect 168972 333240 169022 333296
rect 169022 333240 169036 333296
rect 168972 333236 169036 333240
rect 258396 333236 258460 333300
rect 173756 331876 173820 331940
rect 259684 331740 259748 331804
rect 266308 330380 266372 330444
rect 270540 329156 270604 329220
rect 255268 329020 255332 329084
rect 170996 327796 171060 327860
rect 173572 327660 173636 327724
rect 276244 327660 276308 327724
rect 259500 327116 259564 327180
rect 280292 325756 280356 325820
rect 274588 324940 274652 325004
rect 184796 323580 184860 323644
rect 162532 321540 162596 321604
rect 166396 321540 166460 321604
rect 104940 320588 105004 320652
rect 106044 320588 106108 320652
rect 267780 320104 267844 320108
rect 267780 320048 267830 320104
rect 267830 320048 267844 320104
rect 267780 320044 267844 320048
rect 78444 319364 78508 319428
rect 267780 319364 267844 319428
rect 86724 318004 86788 318068
rect 160692 317596 160756 317660
rect 161244 317596 161308 317660
rect 90220 316644 90284 316708
rect 109540 315284 109604 315348
rect 196020 314876 196084 314940
rect 187556 314060 187620 314124
rect 78260 313924 78324 313988
rect 85804 313924 85868 313988
rect 94452 313924 94516 313988
rect 104940 313924 105004 313988
rect 98500 312428 98564 312492
rect 87460 311204 87524 311268
rect 256740 311204 256804 311268
rect 87092 311068 87156 311132
rect 106412 311068 106476 311132
rect 148180 310388 148244 310452
rect 173020 309300 173084 309364
rect 194548 309028 194612 309092
rect 97948 308484 98012 308548
rect 281580 308348 281644 308412
rect 71084 307668 71148 307732
rect 86540 307668 86604 307732
rect 269620 307668 269684 307732
rect 109540 306988 109604 307052
rect 260972 306988 261036 307052
rect 185348 306716 185412 306780
rect 86172 306580 86236 306644
rect 156644 306308 156708 306372
rect 273300 305764 273364 305828
rect 245700 305628 245764 305692
rect 262444 305628 262508 305692
rect 95188 304268 95252 304332
rect 75868 304132 75932 304196
rect 92980 304132 93044 304196
rect 113220 304132 113284 304196
rect 180564 304132 180628 304196
rect 277164 304132 277228 304196
rect 188476 303724 188540 303788
rect 263732 303724 263796 303788
rect 66116 303588 66180 303652
rect 83044 303588 83108 303652
rect 186820 303588 186884 303652
rect 184060 302500 184124 302564
rect 179276 302288 179340 302292
rect 179276 302232 179326 302288
rect 179326 302232 179340 302288
rect 179276 302228 179340 302232
rect 166212 301744 166276 301748
rect 166212 301688 166262 301744
rect 166262 301688 166276 301744
rect 166212 301684 166276 301688
rect 159772 301548 159836 301612
rect 269620 301412 269684 301476
rect 251772 300868 251836 300932
rect 91508 300188 91572 300252
rect 156644 300052 156708 300116
rect 258764 300732 258828 300796
rect 245700 300596 245764 300660
rect 188292 299780 188356 299844
rect 256740 298692 256804 298756
rect 258764 298012 258828 298076
rect 154436 297332 154500 297396
rect 168420 297392 168484 297396
rect 168420 297336 168470 297392
rect 168470 297336 168484 297392
rect 168420 297332 168484 297336
rect 255268 297332 255332 297396
rect 269804 296788 269868 296852
rect 258396 293932 258460 293996
rect 259684 293524 259748 293588
rect 81940 292572 82004 292636
rect 160692 291756 160756 291820
rect 166212 291756 166276 291820
rect 185348 291756 185412 291820
rect 258396 290804 258460 290868
rect 81020 289852 81084 289916
rect 259684 289716 259748 289780
rect 259500 288764 259564 288828
rect 91508 288492 91572 288556
rect 99972 287676 100036 287740
rect 79180 286996 79244 287060
rect 73292 285772 73356 285836
rect 87092 285772 87156 285836
rect 84700 285560 84764 285564
rect 84700 285504 84714 285560
rect 84714 285504 84764 285560
rect 84700 285500 84764 285504
rect 91140 285500 91204 285564
rect 72924 284276 72988 284340
rect 67404 284140 67468 284204
rect 69244 284140 69308 284204
rect 70164 284140 70228 284204
rect 71636 283732 71700 283796
rect 86724 283596 86788 283660
rect 89852 283520 89916 283524
rect 89852 283464 89866 283520
rect 89866 283464 89916 283520
rect 89852 283460 89916 283464
rect 93716 283460 93780 283524
rect 94268 283460 94332 283524
rect 269804 283460 269868 283524
rect 68692 283188 68756 283252
rect 71820 283188 71884 283252
rect 73108 283188 73172 283252
rect 98868 283188 98932 283252
rect 83412 283112 83476 283116
rect 83412 283056 83462 283112
rect 83462 283056 83476 283112
rect 83412 283052 83476 283056
rect 88748 283052 88812 283116
rect 95372 282976 95436 282980
rect 95372 282920 95386 282976
rect 95386 282920 95436 282976
rect 95372 282916 95436 282920
rect 159772 282916 159836 282980
rect 99972 280196 100036 280260
rect 267780 278836 267844 278900
rect 100708 278700 100772 278764
rect 184060 278020 184124 278084
rect 260972 278156 261036 278220
rect 100708 277748 100772 277812
rect 262444 277340 262508 277404
rect 67404 277204 67468 277268
rect 160692 276660 160756 276724
rect 166212 276660 166276 276724
rect 67404 275980 67468 276044
rect 193812 275300 193876 275364
rect 66300 275164 66364 275228
rect 262260 272716 262324 272780
rect 259316 272444 259380 272508
rect 258396 270812 258460 270876
rect 259132 270812 259196 270876
rect 266492 270132 266556 270196
rect 266492 269180 266556 269244
rect 162716 269044 162780 269108
rect 271092 269104 271156 269108
rect 271092 269048 271142 269104
rect 271142 269048 271156 269104
rect 271092 269044 271156 269048
rect 98868 268364 98932 268428
rect 269620 268364 269684 268428
rect 159956 267004 160020 267068
rect 61700 266460 61764 266524
rect 159956 266324 160020 266388
rect 287100 267140 287164 267204
rect 263364 267004 263428 267068
rect 168420 265508 168484 265572
rect 259132 265508 259196 265572
rect 166396 264828 166460 264892
rect 141372 264148 141436 264212
rect 175780 264148 175844 264212
rect 259132 263604 259196 263668
rect 265940 263468 266004 263532
rect 265940 263060 266004 263124
rect 266308 262924 266372 262988
rect 177988 262788 178052 262852
rect 281580 262108 281644 262172
rect 66300 260944 66364 260948
rect 105492 261428 105556 261492
rect 269068 261156 269132 261220
rect 258580 261020 258644 261084
rect 277900 261292 277964 261356
rect 66300 260888 66350 260944
rect 66350 260888 66364 260944
rect 66300 260884 66364 260888
rect 259132 260884 259196 260948
rect 168236 260808 168300 260812
rect 168236 260752 168250 260808
rect 168250 260752 168300 260808
rect 168236 260748 168300 260752
rect 66300 260068 66364 260132
rect 168236 259796 168300 259860
rect 284340 260068 284404 260132
rect 266492 259720 266556 259724
rect 266492 259664 266506 259720
rect 266506 259664 266556 259720
rect 266492 259660 266556 259664
rect 187556 258844 187620 258908
rect 173020 258708 173084 258772
rect 263548 259116 263612 259180
rect 187556 258028 187620 258092
rect 276428 258028 276492 258092
rect 270724 257892 270788 257956
rect 184796 257348 184860 257412
rect 177804 257212 177868 257276
rect 66668 256804 66732 256868
rect 184796 256668 184860 256732
rect 258580 257076 258644 257140
rect 267964 257076 268028 257140
rect 267964 256940 268028 257004
rect 285628 256668 285692 256732
rect 266308 255852 266372 255916
rect 280292 255852 280356 255916
rect 170812 254280 170876 254284
rect 170812 254224 170826 254280
rect 170826 254224 170876 254280
rect 170812 254220 170876 254224
rect 263548 254008 263612 254012
rect 263548 253952 263598 254008
rect 263598 253952 263612 254008
rect 263548 253948 263612 253952
rect 177620 253812 177684 253876
rect 262260 253268 262324 253332
rect 263364 253268 263428 253332
rect 262444 253132 262508 253196
rect 258396 252724 258460 252788
rect 191788 252588 191852 252652
rect 193996 252588 194060 252652
rect 163452 251908 163516 251972
rect 266308 251908 266372 251972
rect 179276 251772 179340 251836
rect 98316 251228 98380 251292
rect 101260 251092 101324 251156
rect 168420 251092 168484 251156
rect 155724 250412 155788 250476
rect 258396 250004 258460 250068
rect 259316 250004 259380 250068
rect 193444 249052 193508 249116
rect 166764 248372 166828 248436
rect 192340 247692 192404 247756
rect 191788 247420 191852 247484
rect 98132 247148 98196 247212
rect 274588 247012 274652 247076
rect 257292 246332 257356 246396
rect 65932 245380 65996 245444
rect 270540 243612 270604 243676
rect 277532 243672 277596 243676
rect 277532 243616 277546 243672
rect 277546 243616 277596 243672
rect 277532 243612 277596 243616
rect 252876 243204 252940 243268
rect 68692 241708 68756 241772
rect 70900 241768 70964 241772
rect 70900 241712 70950 241768
rect 70950 241712 70964 241768
rect 70900 241708 70964 241712
rect 91508 241708 91572 241772
rect 84700 241572 84764 241636
rect 197860 241980 197924 242044
rect 242940 242040 243004 242044
rect 242940 241984 242990 242040
rect 242990 241984 243004 242040
rect 242940 241980 243004 241984
rect 251036 241980 251100 242044
rect 68876 241496 68940 241500
rect 68876 241440 68890 241496
rect 68890 241440 68940 241496
rect 68876 241436 68940 241440
rect 84332 241300 84396 241364
rect 252876 241028 252940 241092
rect 258396 240892 258460 240956
rect 267780 240484 267844 240548
rect 86540 240076 86604 240140
rect 93532 240136 93596 240140
rect 93532 240080 93546 240136
rect 93546 240080 93596 240136
rect 93532 240076 93596 240080
rect 97764 240076 97828 240140
rect 191788 240076 191852 240140
rect 193996 240076 194060 240140
rect 66116 239940 66180 240004
rect 68876 239940 68940 240004
rect 73108 239940 73172 240004
rect 87460 239940 87524 240004
rect 273484 239940 273548 240004
rect 201540 239396 201604 239460
rect 263732 239396 263796 239460
rect 61884 238716 61948 238780
rect 91140 238580 91204 238644
rect 193812 238580 193876 238644
rect 96660 238444 96724 238508
rect 211660 237900 211724 237964
rect 91508 237356 91572 237420
rect 93900 237356 93964 237420
rect 73476 236676 73540 236740
rect 95188 236676 95252 236740
rect 94268 236540 94332 236604
rect 262444 236540 262508 236604
rect 257292 235996 257356 236060
rect 258396 234500 258460 234564
rect 160692 233140 160756 233204
rect 266492 231236 266556 231300
rect 269068 230284 269132 230348
rect 192340 228788 192404 228852
rect 61700 228244 61764 228308
rect 88748 227700 88812 227764
rect 94084 227700 94148 227764
rect 101260 227700 101324 227764
rect 71452 227564 71516 227628
rect 267964 227564 268028 227628
rect 270724 223484 270788 223548
rect 98132 220900 98196 220964
rect 215340 216684 215404 216748
rect 188476 215868 188540 215932
rect 205588 215868 205652 215932
rect 97948 214508 98012 214572
rect 92980 213148 93044 213212
rect 93532 213148 93596 213212
rect 267780 210292 267844 210356
rect 219572 208252 219636 208316
rect 262076 205668 262140 205732
rect 166212 205532 166276 205596
rect 97764 204308 97828 204372
rect 242940 200636 243004 200700
rect 66116 199276 66180 199340
rect 188844 199276 188908 199340
rect 262260 193836 262324 193900
rect 104020 192476 104084 192540
rect 263548 192476 263612 192540
rect 168420 188260 168484 188324
rect 86540 185540 86604 185604
rect 188292 185540 188356 185604
rect 188292 181324 188356 181388
rect 277900 181324 277964 181388
rect 200620 179964 200684 180028
rect 188292 179420 188356 179484
rect 93716 176760 93780 176764
rect 93716 176704 93730 176760
rect 93730 176704 93780 176760
rect 93716 176700 93780 176704
rect 86724 175748 86788 175812
rect 266308 166908 266372 166972
rect 95188 163372 95252 163436
rect 190316 153716 190380 153780
rect 66668 149092 66732 149156
rect 224908 148412 224972 148476
rect 193812 148276 193876 148340
rect 71636 146372 71700 146436
rect 72924 145072 72988 145076
rect 72924 145016 72938 145072
rect 72938 145016 72988 145072
rect 72924 145012 72988 145016
rect 89852 144740 89916 144804
rect 99972 144740 100036 144804
rect 197860 144800 197924 144804
rect 197860 144744 197910 144800
rect 197910 144744 197924 144800
rect 197860 144740 197924 144744
rect 223620 144740 223684 144804
rect 224356 142428 224420 142492
rect 196572 142292 196636 142356
rect 203196 142156 203260 142220
rect 83412 141340 83476 141404
rect 193076 141068 193140 141132
rect 226380 140660 226444 140724
rect 209820 140524 209884 140588
rect 195100 140388 195164 140452
rect 65932 139980 65996 140044
rect 68692 139572 68756 139636
rect 193076 139028 193140 139092
rect 72924 138348 72988 138412
rect 71820 137940 71884 138004
rect 87092 137592 87156 137596
rect 87092 137536 87106 137592
rect 87106 137536 87156 137592
rect 87092 137532 87156 137536
rect 70164 137396 70228 137460
rect 70164 137260 70228 137324
rect 69428 136580 69492 136644
rect 259500 136580 259564 136644
rect 72372 135084 72436 135148
rect 190316 134540 190380 134604
rect 224356 133452 224420 133516
rect 69428 133316 69492 133380
rect 190316 132500 190380 132564
rect 192708 131956 192772 132020
rect 192708 131412 192772 131476
rect 193444 131412 193508 131476
rect 188292 131140 188356 131204
rect 100708 129236 100772 129300
rect 224356 128964 224420 129028
rect 192340 123796 192404 123860
rect 224908 121348 224972 121412
rect 226380 119444 226444 119508
rect 106780 119308 106844 119372
rect 65932 116996 65996 117060
rect 66484 109380 66548 109444
rect 94084 109108 94148 109172
rect 188844 107748 188908 107812
rect 227668 108292 227732 108356
rect 270540 108292 270604 108356
rect 66668 106932 66732 106996
rect 94268 106116 94332 106180
rect 98500 105028 98564 105092
rect 104020 103532 104084 103596
rect 193812 102172 193876 102236
rect 224356 99452 224420 99516
rect 226380 97140 226444 97204
rect 189948 96868 190012 96932
rect 66116 96324 66180 96388
rect 97212 96052 97276 96116
rect 94820 95780 94884 95844
rect 273300 95780 273364 95844
rect 69428 94012 69492 94076
rect 200620 93332 200684 93396
rect 209820 93332 209884 93396
rect 68692 92652 68756 92716
rect 72372 92652 72436 92716
rect 68876 92516 68940 92580
rect 192340 92516 192404 92580
rect 71452 92380 71516 92444
rect 91692 92380 91756 92444
rect 92980 92380 93044 92444
rect 201540 92380 201604 92444
rect 211660 92380 211724 92444
rect 61884 92244 61948 92308
rect 72924 92244 72988 92308
rect 224356 92244 224420 92308
rect 251772 92108 251836 92172
rect 94820 91972 94884 92036
rect 251772 91700 251836 91764
rect 219204 91080 219268 91084
rect 219204 91024 219218 91080
rect 219218 91024 219268 91080
rect 219204 91020 219268 91024
rect 205588 90264 205652 90268
rect 205588 90208 205638 90264
rect 205638 90208 205652 90264
rect 205588 90204 205652 90208
rect 215340 90264 215404 90268
rect 215340 90208 215354 90264
rect 215354 90208 215404 90264
rect 215340 90204 215404 90208
rect 95188 89796 95252 89860
rect 70164 89524 70228 89588
rect 227668 87892 227732 87956
rect 189948 86668 190012 86732
rect 226380 86668 226444 86732
rect 192708 86124 192772 86188
rect 193812 85444 193876 85508
rect 194548 85444 194612 85508
rect 66484 85172 66548 85236
rect 194548 84764 194612 84828
rect 69612 83948 69676 84012
rect 195100 82044 195164 82108
rect 196572 79324 196636 79388
rect 97212 75788 97276 75852
rect 168236 72388 168300 72452
rect 105492 55796 105556 55860
rect 141372 44780 141436 44844
rect 144132 43420 144196 43484
rect 203196 40564 203260 40628
rect 166212 30908 166276 30972
rect 106780 28188 106844 28252
rect 175780 26828 175844 26892
rect 124812 15812 124876 15876
rect 186820 6156 186884 6220
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 72923 699820 72989 699821
rect 72923 699756 72924 699820
rect 72988 699756 72989 699820
rect 72923 699755 72989 699756
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 583166 67574 608058
rect 70899 580820 70965 580821
rect 70899 580756 70900 580820
rect 70964 580756 70965 580820
rect 70899 580755 70965 580756
rect 66667 578644 66733 578645
rect 66667 578580 66668 578644
rect 66732 578580 66733 578644
rect 66667 578579 66733 578580
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 66115 526420 66181 526421
rect 66115 526356 66116 526420
rect 66180 526356 66181 526420
rect 66115 526355 66181 526356
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 66118 466581 66178 526355
rect 66115 466580 66181 466581
rect 66115 466516 66116 466580
rect 66180 466516 66181 466580
rect 66115 466515 66181 466516
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66118 423333 66178 466515
rect 66115 423332 66181 423333
rect 66115 423268 66116 423332
rect 66180 423268 66181 423332
rect 66115 423267 66181 423268
rect 66670 402661 66730 578579
rect 67771 562052 67837 562053
rect 67771 561988 67772 562052
rect 67836 561988 67837 562052
rect 67771 561987 67837 561988
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 67774 465765 67834 561987
rect 69427 551172 69493 551173
rect 69427 551108 69428 551172
rect 69492 551170 69493 551172
rect 69492 551110 69674 551170
rect 69492 551108 69493 551110
rect 69427 551107 69493 551108
rect 69427 549540 69493 549541
rect 69427 549476 69428 549540
rect 69492 549476 69493 549540
rect 69427 549475 69493 549476
rect 67955 543420 68021 543421
rect 67955 543356 67956 543420
rect 68020 543356 68021 543420
rect 67955 543355 68021 543356
rect 67958 521661 68018 543355
rect 69430 536890 69490 549475
rect 69614 539069 69674 551110
rect 69611 539068 69677 539069
rect 69611 539004 69612 539068
rect 69676 539004 69677 539068
rect 69611 539003 69677 539004
rect 69430 536830 69858 536890
rect 69611 536212 69677 536213
rect 69611 536148 69612 536212
rect 69676 536148 69677 536212
rect 69611 536147 69677 536148
rect 67955 521660 68021 521661
rect 67955 521596 67956 521660
rect 68020 521596 68021 521660
rect 67955 521595 68021 521596
rect 68875 521660 68941 521661
rect 68875 521596 68876 521660
rect 68940 521596 68941 521660
rect 68875 521595 68941 521596
rect 68878 467941 68938 521595
rect 69614 516765 69674 536147
rect 69798 530637 69858 536830
rect 69795 530636 69861 530637
rect 69795 530572 69796 530636
rect 69860 530572 69861 530636
rect 69795 530571 69861 530572
rect 69611 516764 69677 516765
rect 69611 516700 69612 516764
rect 69676 516700 69677 516764
rect 69611 516699 69677 516700
rect 68875 467940 68941 467941
rect 68875 467876 68876 467940
rect 68940 467876 68941 467940
rect 68875 467875 68941 467876
rect 67771 465764 67837 465765
rect 67771 465700 67772 465764
rect 67836 465700 67837 465764
rect 67771 465699 67837 465700
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 436356 67574 464058
rect 70902 448629 70962 580755
rect 72926 539613 72986 699755
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 583166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 583166 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 583166 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 583166 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 583166 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 75683 580956 75749 580957
rect 75683 580892 75684 580956
rect 75748 580892 75749 580956
rect 75683 580891 75749 580892
rect 73679 543454 73999 543486
rect 73679 543218 73721 543454
rect 73957 543218 73999 543454
rect 73679 543134 73999 543218
rect 73679 542898 73721 543134
rect 73957 542898 73999 543134
rect 73679 542866 73999 542898
rect 72923 539612 72989 539613
rect 72923 539548 72924 539612
rect 72988 539548 72989 539612
rect 72923 539547 72989 539548
rect 72739 512684 72805 512685
rect 72739 512620 72740 512684
rect 72804 512620 72805 512684
rect 72739 512619 72805 512620
rect 70899 448628 70965 448629
rect 70899 448564 70900 448628
rect 70964 448564 70965 448628
rect 70899 448563 70965 448564
rect 69611 447812 69677 447813
rect 69611 447748 69612 447812
rect 69676 447748 69677 447812
rect 69611 447747 69677 447748
rect 69614 441630 69674 447747
rect 69430 441570 69674 441630
rect 69243 434348 69309 434349
rect 69243 434284 69244 434348
rect 69308 434284 69309 434348
rect 69243 434283 69309 434284
rect 67955 433940 68021 433941
rect 67955 433876 67956 433940
rect 68020 433876 68021 433940
rect 67955 433875 68021 433876
rect 67958 422245 68018 433875
rect 67955 422244 68021 422245
rect 67955 422180 67956 422244
rect 68020 422180 68021 422244
rect 67955 422179 68021 422180
rect 66667 402660 66733 402661
rect 66667 402596 66668 402660
rect 66732 402596 66733 402660
rect 66667 402595 66733 402596
rect 66299 397356 66365 397357
rect 66299 397292 66300 397356
rect 66364 397292 66365 397356
rect 66299 397291 66365 397292
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 66115 303652 66181 303653
rect 66115 303588 66116 303652
rect 66180 303588 66181 303652
rect 66115 303587 66181 303588
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 61699 266524 61765 266525
rect 61699 266460 61700 266524
rect 61764 266460 61765 266524
rect 61699 266459 61765 266460
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 61702 228309 61762 266459
rect 63234 244894 63854 280338
rect 65931 245444 65997 245445
rect 65931 245380 65932 245444
rect 65996 245380 65997 245444
rect 65931 245379 65997 245380
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 61883 238780 61949 238781
rect 61883 238716 61884 238780
rect 61948 238716 61949 238780
rect 61883 238715 61949 238716
rect 61699 228308 61765 228309
rect 61699 228244 61700 228308
rect 61764 228244 61765 228308
rect 61699 228243 61765 228244
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 61886 92309 61946 238715
rect 63234 208894 63854 244338
rect 65934 209790 65994 245379
rect 66118 240005 66178 303587
rect 66302 275229 66362 397291
rect 66954 356614 67574 388356
rect 68875 357372 68941 357373
rect 68875 357308 68876 357372
rect 68940 357308 68941 357372
rect 68875 357307 68941 357308
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 285592 67574 320058
rect 67403 284204 67469 284205
rect 67403 284140 67404 284204
rect 67468 284140 67469 284204
rect 67403 284139 67469 284140
rect 67406 277269 67466 284139
rect 68691 283252 68757 283253
rect 68691 283188 68692 283252
rect 68756 283188 68757 283252
rect 68691 283187 68757 283188
rect 67403 277268 67469 277269
rect 67403 277204 67404 277268
rect 67468 277204 67469 277268
rect 67403 277203 67469 277204
rect 67406 276045 67466 277203
rect 67403 276044 67469 276045
rect 67403 275980 67404 276044
rect 67468 275980 67469 276044
rect 67403 275979 67469 275980
rect 66299 275228 66365 275229
rect 66299 275164 66300 275228
rect 66364 275164 66365 275228
rect 66299 275163 66365 275164
rect 66299 260948 66365 260949
rect 66299 260884 66300 260948
rect 66364 260884 66365 260948
rect 66299 260883 66365 260884
rect 66302 260133 66362 260883
rect 66299 260132 66365 260133
rect 66299 260068 66300 260132
rect 66364 260068 66365 260132
rect 66299 260067 66365 260068
rect 66667 256868 66733 256869
rect 66667 256804 66668 256868
rect 66732 256804 66733 256868
rect 66667 256803 66733 256804
rect 66115 240004 66181 240005
rect 66115 239940 66116 240004
rect 66180 239940 66181 240004
rect 66115 239939 66181 239940
rect 65934 209730 66178 209790
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 66118 199341 66178 209730
rect 66115 199340 66181 199341
rect 66115 199276 66116 199340
rect 66180 199276 66181 199340
rect 66115 199275 66181 199276
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 65931 140044 65997 140045
rect 65931 139980 65932 140044
rect 65996 139980 65997 140044
rect 65931 139979 65997 139980
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 65934 117061 65994 139979
rect 65931 117060 65997 117061
rect 65931 116996 65932 117060
rect 65996 116996 65997 117060
rect 65931 116995 65997 116996
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 61883 92308 61949 92309
rect 61883 92244 61884 92308
rect 61948 92244 61949 92308
rect 61883 92243 61949 92244
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 64894 63854 100338
rect 66118 96389 66178 199275
rect 66670 149157 66730 256803
rect 68694 241773 68754 283187
rect 68691 241772 68757 241773
rect 68691 241708 68692 241772
rect 68756 241708 68757 241772
rect 68691 241707 68757 241708
rect 68878 241501 68938 357307
rect 69246 284205 69306 434283
rect 69430 433125 69490 441570
rect 71083 436116 71149 436117
rect 71083 436052 71084 436116
rect 71148 436052 71149 436116
rect 71083 436051 71149 436052
rect 69427 433124 69493 433125
rect 69427 433060 69428 433124
rect 69492 433060 69493 433124
rect 69427 433059 69493 433060
rect 70899 369068 70965 369069
rect 70899 369004 70900 369068
rect 70964 369004 70965 369068
rect 70899 369003 70965 369004
rect 69243 284204 69309 284205
rect 69243 284140 69244 284204
rect 69308 284140 69309 284204
rect 69243 284139 69309 284140
rect 70163 284204 70229 284205
rect 70163 284140 70164 284204
rect 70228 284140 70229 284204
rect 70163 284139 70229 284140
rect 68875 241500 68941 241501
rect 68875 241436 68876 241500
rect 68940 241436 68941 241500
rect 68875 241435 68941 241436
rect 68875 240004 68941 240005
rect 68875 239940 68876 240004
rect 68940 239940 68941 240004
rect 68875 239939 68941 239940
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66667 149156 66733 149157
rect 66667 149092 66668 149156
rect 66732 149092 66733 149156
rect 66667 149091 66733 149092
rect 66483 109444 66549 109445
rect 66483 109380 66484 109444
rect 66548 109380 66549 109444
rect 66483 109379 66549 109380
rect 66115 96388 66181 96389
rect 66115 96324 66116 96388
rect 66180 96324 66181 96388
rect 66115 96323 66181 96324
rect 66486 85237 66546 109379
rect 66670 106997 66730 149091
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 136782 67574 140058
rect 68691 139636 68757 139637
rect 68691 139572 68692 139636
rect 68756 139572 68757 139636
rect 68691 139571 68757 139572
rect 66667 106996 66733 106997
rect 66667 106932 66668 106996
rect 66732 106932 66733 106996
rect 66667 106931 66733 106932
rect 68694 92717 68754 139571
rect 68691 92716 68757 92717
rect 68691 92652 68692 92716
rect 68756 92652 68757 92716
rect 68691 92651 68757 92652
rect 68878 92581 68938 239939
rect 70166 137461 70226 284139
rect 70902 241773 70962 369003
rect 71086 307733 71146 436051
rect 72742 390965 72802 512619
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 75686 500173 75746 580891
rect 79915 580820 79981 580821
rect 79915 580756 79916 580820
rect 79980 580756 79981 580820
rect 79915 580755 79981 580756
rect 84699 580820 84765 580821
rect 84699 580756 84700 580820
rect 84764 580756 84765 580820
rect 84699 580755 84765 580756
rect 89299 580820 89365 580821
rect 89299 580756 89300 580820
rect 89364 580756 89365 580820
rect 89299 580755 89365 580756
rect 77644 561454 77964 561486
rect 77644 561218 77686 561454
rect 77922 561218 77964 561454
rect 77644 561134 77964 561218
rect 77644 560898 77686 561134
rect 77922 560898 77964 561134
rect 77644 560866 77964 560898
rect 77155 520980 77221 520981
rect 77155 520916 77156 520980
rect 77220 520916 77221 520980
rect 77155 520915 77221 520916
rect 75683 500172 75749 500173
rect 75683 500108 75684 500172
rect 75748 500108 75749 500172
rect 75683 500107 75749 500108
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73475 436524 73541 436525
rect 73475 436460 73476 436524
rect 73540 436460 73541 436524
rect 73475 436459 73541 436460
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 72739 390964 72805 390965
rect 72739 390900 72740 390964
rect 72804 390900 72805 390964
rect 72739 390899 72805 390900
rect 72742 388925 72802 390899
rect 72739 388924 72805 388925
rect 72739 388860 72740 388924
rect 72804 388860 72805 388924
rect 72739 388859 72805 388860
rect 71083 307732 71149 307733
rect 71083 307668 71084 307732
rect 71148 307668 71149 307732
rect 71083 307667 71149 307668
rect 73478 292590 73538 436459
rect 73794 436356 74414 470898
rect 75131 436252 75197 436253
rect 75131 436188 75132 436252
rect 75196 436188 75197 436252
rect 75131 436187 75197 436188
rect 74763 433668 74829 433669
rect 74763 433604 74764 433668
rect 74828 433604 74829 433668
rect 74763 433603 74829 433604
rect 73110 292530 73538 292590
rect 73794 363454 74414 388356
rect 74766 385117 74826 433603
rect 75134 387701 75194 436187
rect 75867 433668 75933 433669
rect 75867 433604 75868 433668
rect 75932 433604 75933 433668
rect 75867 433603 75933 433604
rect 75131 387700 75197 387701
rect 75131 387636 75132 387700
rect 75196 387636 75197 387700
rect 75131 387635 75197 387636
rect 74763 385116 74829 385117
rect 74763 385052 74764 385116
rect 74828 385052 74829 385116
rect 74763 385051 74829 385052
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 72923 284340 72989 284341
rect 72923 284276 72924 284340
rect 72988 284276 72989 284340
rect 72923 284275 72989 284276
rect 71635 283796 71701 283797
rect 71635 283732 71636 283796
rect 71700 283732 71701 283796
rect 71635 283731 71701 283732
rect 70899 241772 70965 241773
rect 70899 241708 70900 241772
rect 70964 241708 70965 241772
rect 70899 241707 70965 241708
rect 71451 227628 71517 227629
rect 71451 227564 71452 227628
rect 71516 227564 71517 227628
rect 71451 227563 71517 227564
rect 70163 137460 70229 137461
rect 70163 137396 70164 137460
rect 70228 137396 70229 137460
rect 70163 137395 70229 137396
rect 70163 137324 70229 137325
rect 70163 137260 70164 137324
rect 70228 137260 70229 137324
rect 70163 137259 70229 137260
rect 69427 136644 69493 136645
rect 69427 136580 69428 136644
rect 69492 136580 69493 136644
rect 69427 136579 69493 136580
rect 69430 133381 69490 136579
rect 69427 133380 69493 133381
rect 69427 133316 69428 133380
rect 69492 133316 69493 133380
rect 69427 133315 69493 133316
rect 69427 94076 69493 94077
rect 69427 94012 69428 94076
rect 69492 94012 69493 94076
rect 69427 94011 69493 94012
rect 69430 93870 69490 94011
rect 69430 93810 69674 93870
rect 68875 92580 68941 92581
rect 68875 92516 68876 92580
rect 68940 92516 68941 92580
rect 68875 92515 68941 92516
rect 66483 85236 66549 85237
rect 66483 85172 66484 85236
rect 66548 85172 66549 85236
rect 66483 85171 66549 85172
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 90782
rect 69614 84013 69674 93810
rect 70166 89589 70226 137259
rect 71454 92445 71514 227563
rect 71638 146437 71698 283731
rect 71819 283252 71885 283253
rect 71819 283188 71820 283252
rect 71884 283188 71885 283252
rect 71819 283187 71885 283188
rect 71635 146436 71701 146437
rect 71635 146372 71636 146436
rect 71700 146372 71701 146436
rect 71635 146371 71701 146372
rect 71822 138005 71882 283187
rect 72926 145077 72986 284275
rect 73110 283253 73170 292530
rect 73794 291454 74414 326898
rect 75870 304197 75930 433603
rect 77158 390421 77218 520915
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 436356 78134 438618
rect 79179 436388 79245 436389
rect 79179 436324 79180 436388
rect 79244 436324 79245 436388
rect 79179 436323 79245 436324
rect 78443 433804 78509 433805
rect 78443 433740 78444 433804
rect 78508 433740 78509 433804
rect 78443 433739 78509 433740
rect 78259 433668 78325 433669
rect 78259 433604 78260 433668
rect 78324 433604 78325 433668
rect 78259 433603 78325 433604
rect 77155 390420 77221 390421
rect 77155 390356 77156 390420
rect 77220 390356 77221 390420
rect 77155 390355 77221 390356
rect 78262 388517 78322 433603
rect 78259 388516 78325 388517
rect 78259 388452 78260 388516
rect 78324 388452 78325 388516
rect 78259 388451 78325 388452
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 75867 304196 75933 304197
rect 75867 304132 75868 304196
rect 75932 304132 75933 304196
rect 75867 304131 75933 304132
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73291 285836 73357 285837
rect 73291 285772 73292 285836
rect 73356 285772 73357 285836
rect 73291 285771 73357 285772
rect 73107 283252 73173 283253
rect 73107 283188 73108 283252
rect 73172 283188 73173 283252
rect 73107 283187 73173 283188
rect 73110 240005 73170 283187
rect 73294 277410 73354 285771
rect 73794 285592 74414 290898
rect 77514 295174 78134 330618
rect 78446 319429 78506 433739
rect 78443 319428 78509 319429
rect 78443 319364 78444 319428
rect 78508 319364 78509 319428
rect 78443 319363 78509 319364
rect 78446 316050 78506 319363
rect 78262 315990 78506 316050
rect 78262 313989 78322 315990
rect 78259 313988 78325 313989
rect 78259 313924 78260 313988
rect 78324 313924 78325 313988
rect 78259 313923 78325 313924
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285592 78134 294618
rect 79182 287061 79242 436323
rect 79918 390829 79978 580755
rect 81609 543454 81929 543486
rect 81609 543218 81651 543454
rect 81887 543218 81929 543454
rect 81609 543134 81929 543218
rect 81609 542898 81651 543134
rect 81887 542898 81929 543134
rect 81609 542866 81929 542898
rect 81234 514894 81854 537166
rect 82859 530636 82925 530637
rect 82859 530572 82860 530636
rect 82924 530572 82925 530636
rect 82859 530571 82925 530572
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 436356 81854 442338
rect 81019 436252 81085 436253
rect 81019 436188 81020 436252
rect 81084 436188 81085 436252
rect 81019 436187 81085 436188
rect 80651 434076 80717 434077
rect 80651 434012 80652 434076
rect 80716 434012 80717 434076
rect 80651 434011 80717 434012
rect 79915 390828 79981 390829
rect 79915 390764 79916 390828
rect 79980 390764 79981 390828
rect 79915 390763 79981 390764
rect 80654 388517 80714 434011
rect 80651 388516 80717 388517
rect 80651 388452 80652 388516
rect 80716 388452 80717 388516
rect 80651 388451 80717 388452
rect 81022 289917 81082 436187
rect 81939 433668 82005 433669
rect 81939 433604 81940 433668
rect 82004 433604 82005 433668
rect 81939 433603 82005 433604
rect 82491 433668 82557 433669
rect 82491 433604 82492 433668
rect 82556 433604 82557 433668
rect 82491 433603 82557 433604
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81942 339557 82002 433603
rect 82494 388517 82554 433603
rect 82862 390829 82922 530571
rect 83043 433668 83109 433669
rect 83043 433604 83044 433668
rect 83108 433604 83109 433668
rect 83043 433603 83109 433604
rect 84515 433668 84581 433669
rect 84515 433604 84516 433668
rect 84580 433604 84581 433668
rect 84515 433603 84581 433604
rect 82859 390828 82925 390829
rect 82859 390764 82860 390828
rect 82924 390764 82925 390828
rect 82859 390763 82925 390764
rect 82491 388516 82557 388517
rect 82491 388452 82492 388516
rect 82556 388452 82557 388516
rect 82491 388451 82557 388452
rect 81939 339556 82005 339557
rect 81939 339492 81940 339556
rect 82004 339492 82005 339556
rect 81939 339491 82005 339492
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81019 289916 81085 289917
rect 81019 289852 81020 289916
rect 81084 289852 81085 289916
rect 81019 289851 81085 289852
rect 79179 287060 79245 287061
rect 79179 286996 79180 287060
rect 79244 286996 79245 287060
rect 79179 286995 79245 286996
rect 81234 285592 81854 298338
rect 81942 292637 82002 339491
rect 83046 303653 83106 433603
rect 84518 390965 84578 433603
rect 84515 390964 84581 390965
rect 84515 390900 84516 390964
rect 84580 390900 84581 390964
rect 84515 390899 84581 390900
rect 84702 390557 84762 580755
rect 85575 561454 85895 561486
rect 85575 561218 85617 561454
rect 85853 561218 85895 561454
rect 85575 561134 85895 561218
rect 85575 560898 85617 561134
rect 85853 560898 85895 561134
rect 85575 560866 85895 560898
rect 84954 518614 85574 537166
rect 88195 535532 88261 535533
rect 88195 535468 88196 535532
rect 88260 535468 88261 535532
rect 88195 535467 88261 535468
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 436356 85574 446058
rect 86723 433804 86789 433805
rect 86723 433740 86724 433804
rect 86788 433740 86789 433804
rect 86723 433739 86789 433740
rect 85803 433668 85869 433669
rect 85803 433604 85804 433668
rect 85868 433604 85869 433668
rect 85803 433603 85869 433604
rect 84699 390556 84765 390557
rect 84699 390492 84700 390556
rect 84764 390492 84765 390556
rect 84699 390491 84765 390492
rect 83963 388380 84029 388381
rect 83963 388316 83964 388380
rect 84028 388316 84029 388380
rect 83963 388315 84029 388316
rect 83043 303652 83109 303653
rect 83043 303588 83044 303652
rect 83108 303588 83109 303652
rect 83043 303587 83109 303588
rect 81939 292636 82005 292637
rect 81939 292572 81940 292636
rect 82004 292572 82005 292636
rect 81939 292571 82005 292572
rect 83966 292590 84026 388315
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 85806 313989 85866 433603
rect 86726 318069 86786 433739
rect 87091 433668 87157 433669
rect 87091 433604 87092 433668
rect 87156 433604 87157 433668
rect 87091 433603 87157 433604
rect 86723 318068 86789 318069
rect 86723 318004 86724 318068
rect 86788 318004 86789 318068
rect 86723 318003 86789 318004
rect 86726 316050 86786 318003
rect 86174 315990 86786 316050
rect 85803 313988 85869 313989
rect 85803 313924 85804 313988
rect 85868 313924 85869 313988
rect 85803 313923 85869 313924
rect 86174 306645 86234 315990
rect 87094 311133 87154 433603
rect 88198 389333 88258 535467
rect 89302 482901 89362 580755
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 96659 553484 96725 553485
rect 96659 553420 96660 553484
rect 96724 553420 96725 553484
rect 96659 553419 96725 553420
rect 96662 551309 96722 553419
rect 96659 551308 96725 551309
rect 96659 551244 96660 551308
rect 96724 551244 96725 551308
rect 96659 551243 96725 551244
rect 96843 547092 96909 547093
rect 96843 547028 96844 547092
rect 96908 547028 96909 547092
rect 96843 547027 96909 547028
rect 89540 543454 89860 543486
rect 89540 543218 89582 543454
rect 89818 543218 89860 543454
rect 89540 543134 89860 543218
rect 89540 542898 89582 543134
rect 89818 542898 89860 543134
rect 89540 542866 89860 542898
rect 91794 525454 92414 537166
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 89299 482900 89365 482901
rect 89299 482836 89300 482900
rect 89364 482836 89365 482900
rect 89299 482835 89365 482836
rect 91323 465764 91389 465765
rect 91323 465700 91324 465764
rect 91388 465700 91389 465764
rect 91323 465699 91389 465700
rect 89667 433668 89733 433669
rect 89667 433604 89668 433668
rect 89732 433604 89733 433668
rect 89667 433603 89733 433604
rect 90219 433668 90285 433669
rect 90219 433604 90220 433668
rect 90284 433604 90285 433668
rect 90219 433603 90285 433604
rect 89670 433530 89730 433603
rect 89486 433470 89730 433530
rect 89486 427830 89546 433470
rect 89486 427770 89730 427830
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 89670 398850 89730 427770
rect 89486 398790 89730 398850
rect 88195 389332 88261 389333
rect 88195 389268 88196 389332
rect 88260 389268 88261 389332
rect 88195 389267 88261 389268
rect 89486 389190 89546 398790
rect 89486 389130 89730 389190
rect 89670 387293 89730 389130
rect 89667 387292 89733 387293
rect 89667 387228 89668 387292
rect 89732 387228 89733 387292
rect 89667 387227 89733 387228
rect 90222 316709 90282 433603
rect 91326 390421 91386 465699
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 436356 92414 452898
rect 95514 529174 96134 537166
rect 96659 529276 96725 529277
rect 96659 529212 96660 529276
rect 96724 529212 96725 529276
rect 96659 529211 96725 529212
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 436356 96134 456618
rect 94451 436116 94517 436117
rect 94451 436052 94452 436116
rect 94516 436052 94517 436116
rect 94451 436051 94517 436052
rect 92795 434212 92861 434213
rect 92795 434148 92796 434212
rect 92860 434148 92861 434212
rect 92795 434147 92861 434148
rect 91507 433668 91573 433669
rect 91507 433604 91508 433668
rect 91572 433604 91573 433668
rect 91507 433603 91573 433604
rect 91323 390420 91389 390421
rect 91323 390356 91324 390420
rect 91388 390356 91389 390420
rect 91323 390355 91389 390356
rect 90219 316708 90285 316709
rect 90219 316644 90220 316708
rect 90284 316644 90285 316708
rect 90219 316643 90285 316644
rect 87459 311268 87525 311269
rect 87459 311204 87460 311268
rect 87524 311204 87525 311268
rect 87459 311203 87525 311204
rect 87091 311132 87157 311133
rect 87091 311068 87092 311132
rect 87156 311068 87157 311132
rect 87091 311067 87157 311068
rect 86539 307732 86605 307733
rect 86539 307668 86540 307732
rect 86604 307668 86605 307732
rect 86539 307667 86605 307668
rect 86171 306644 86237 306645
rect 86171 306580 86172 306644
rect 86236 306580 86237 306644
rect 86171 306579 86237 306580
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 83966 292530 84210 292590
rect 83411 283116 83477 283117
rect 83411 283052 83412 283116
rect 83476 283052 83477 283116
rect 83411 283051 83477 283052
rect 73294 277350 73538 277410
rect 73107 240004 73173 240005
rect 73107 239940 73108 240004
rect 73172 239940 73173 240004
rect 73107 239939 73173 239940
rect 73478 236741 73538 277350
rect 78977 273454 79297 273486
rect 78977 273218 79019 273454
rect 79255 273218 79297 273454
rect 78977 273134 79297 273218
rect 78977 272898 79019 273134
rect 79255 272898 79297 273134
rect 78977 272866 79297 272898
rect 74345 255454 74665 255486
rect 74345 255218 74387 255454
rect 74623 255218 74665 255454
rect 74345 255134 74665 255218
rect 74345 254898 74387 255134
rect 74623 254898 74665 255134
rect 74345 254866 74665 254898
rect 73475 236740 73541 236741
rect 73475 236676 73476 236740
rect 73540 236676 73541 236740
rect 73475 236675 73541 236676
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 72923 145076 72989 145077
rect 72923 145012 72924 145076
rect 72988 145012 72989 145076
rect 72923 145011 72989 145012
rect 72923 138412 72989 138413
rect 72923 138348 72924 138412
rect 72988 138348 72989 138412
rect 72923 138347 72989 138348
rect 71819 138004 71885 138005
rect 71819 137940 71820 138004
rect 71884 137940 71885 138004
rect 71819 137939 71885 137940
rect 72371 135148 72437 135149
rect 72371 135084 72372 135148
rect 72436 135084 72437 135148
rect 72371 135083 72437 135084
rect 72374 92717 72434 135083
rect 72371 92716 72437 92717
rect 72371 92652 72372 92716
rect 72436 92652 72437 92716
rect 72371 92651 72437 92652
rect 71451 92444 71517 92445
rect 71451 92380 71452 92444
rect 71516 92380 71517 92444
rect 71451 92379 71517 92380
rect 72926 92309 72986 138347
rect 73794 136782 74414 146898
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 136782 78134 150618
rect 81234 226894 81854 239592
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 136782 81854 154338
rect 83414 141405 83474 283051
rect 84150 282930 84210 292530
rect 84954 285592 85574 302058
rect 84699 285564 84765 285565
rect 84699 285500 84700 285564
rect 84764 285500 84765 285564
rect 84699 285499 84765 285500
rect 83966 282870 84210 282930
rect 83966 281890 84026 282870
rect 83966 281830 84394 281890
rect 83609 255454 83929 255486
rect 83609 255218 83651 255454
rect 83887 255218 83929 255454
rect 83609 255134 83929 255218
rect 83609 254898 83651 255134
rect 83887 254898 83929 255134
rect 83609 254866 83929 254898
rect 84334 241365 84394 281830
rect 84702 241637 84762 285499
rect 84699 241636 84765 241637
rect 84699 241572 84700 241636
rect 84764 241572 84765 241636
rect 84699 241571 84765 241572
rect 84331 241364 84397 241365
rect 84331 241300 84332 241364
rect 84396 241300 84397 241364
rect 84331 241299 84397 241300
rect 86542 240141 86602 307667
rect 87091 285836 87157 285837
rect 87091 285772 87092 285836
rect 87156 285772 87157 285836
rect 87091 285771 87157 285772
rect 86723 283660 86789 283661
rect 86723 283596 86724 283660
rect 86788 283596 86789 283660
rect 86723 283595 86789 283596
rect 86539 240140 86605 240141
rect 86539 240076 86540 240140
rect 86604 240076 86605 240140
rect 86539 240075 86605 240076
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 86542 185605 86602 240075
rect 86539 185604 86605 185605
rect 86539 185540 86540 185604
rect 86604 185540 86605 185604
rect 86539 185539 86605 185540
rect 86726 175813 86786 283595
rect 86723 175812 86789 175813
rect 86723 175748 86724 175812
rect 86788 175748 86789 175812
rect 86723 175747 86789 175748
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 83411 141404 83477 141405
rect 83411 141340 83412 141404
rect 83476 141340 83477 141404
rect 83411 141339 83477 141340
rect 84954 136782 85574 158058
rect 87094 137597 87154 285771
rect 87462 240005 87522 311203
rect 91510 300253 91570 433603
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 92798 370565 92858 434147
rect 92979 433668 93045 433669
rect 92979 433604 92980 433668
rect 93044 433604 93045 433668
rect 92979 433603 93045 433604
rect 92795 370564 92861 370565
rect 92795 370500 92796 370564
rect 92860 370500 92861 370564
rect 92795 370499 92861 370500
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91507 300252 91573 300253
rect 91507 300188 91508 300252
rect 91572 300188 91573 300252
rect 91507 300187 91573 300188
rect 91507 288556 91573 288557
rect 91507 288492 91508 288556
rect 91572 288492 91573 288556
rect 91507 288491 91573 288492
rect 91139 285564 91205 285565
rect 91139 285500 91140 285564
rect 91204 285500 91205 285564
rect 91139 285499 91205 285500
rect 89851 283524 89917 283525
rect 89851 283460 89852 283524
rect 89916 283460 89917 283524
rect 89851 283459 89917 283460
rect 88747 283116 88813 283117
rect 88747 283052 88748 283116
rect 88812 283052 88813 283116
rect 88747 283051 88813 283052
rect 88241 273454 88561 273486
rect 88241 273218 88283 273454
rect 88519 273218 88561 273454
rect 88241 273134 88561 273218
rect 88241 272898 88283 273134
rect 88519 272898 88561 273134
rect 88241 272866 88561 272898
rect 87459 240004 87525 240005
rect 87459 239940 87460 240004
rect 87524 239940 87525 240004
rect 87459 239939 87525 239940
rect 88750 227765 88810 283051
rect 88747 227764 88813 227765
rect 88747 227700 88748 227764
rect 88812 227700 88813 227764
rect 88747 227699 88813 227700
rect 89854 144805 89914 283459
rect 91142 238645 91202 285499
rect 91510 241773 91570 288491
rect 91794 285592 92414 308898
rect 92982 304197 93042 433603
rect 94454 313989 94514 436051
rect 95187 434348 95253 434349
rect 95187 434284 95188 434348
rect 95252 434284 95253 434348
rect 95187 434283 95253 434284
rect 94451 313988 94517 313989
rect 94451 313924 94452 313988
rect 94516 313924 94517 313988
rect 94451 313923 94517 313924
rect 95190 304333 95250 434283
rect 96662 390421 96722 529211
rect 96846 519485 96906 547027
rect 99234 532894 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 101259 549404 101325 549405
rect 101259 549340 101260 549404
rect 101324 549340 101325 549404
rect 101259 549339 101325 549340
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 96843 519484 96909 519485
rect 96843 519420 96844 519484
rect 96908 519420 96909 519484
rect 96843 519419 96909 519420
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 436356 99854 460338
rect 100155 434348 100221 434349
rect 100155 434284 100156 434348
rect 100220 434284 100221 434348
rect 100155 434283 100221 434284
rect 98499 433804 98565 433805
rect 98499 433740 98500 433804
rect 98564 433740 98565 433804
rect 98499 433739 98565 433740
rect 97947 433668 98013 433669
rect 97947 433604 97948 433668
rect 98012 433604 98013 433668
rect 97947 433603 98013 433604
rect 96659 390420 96725 390421
rect 96659 390356 96660 390420
rect 96724 390356 96725 390420
rect 96659 390355 96725 390356
rect 95514 385174 96134 388356
rect 96659 387836 96725 387837
rect 96659 387772 96660 387836
rect 96724 387772 96725 387836
rect 96659 387771 96725 387772
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95187 304332 95253 304333
rect 95187 304268 95188 304332
rect 95252 304268 95253 304332
rect 95187 304267 95253 304268
rect 92979 304196 93045 304197
rect 92979 304132 92980 304196
rect 93044 304132 93045 304196
rect 92979 304131 93045 304132
rect 95514 285592 96134 312618
rect 93715 283524 93781 283525
rect 93715 283460 93716 283524
rect 93780 283460 93781 283524
rect 93715 283459 93781 283460
rect 94267 283524 94333 283525
rect 94267 283460 94268 283524
rect 94332 283460 94333 283524
rect 94267 283459 94333 283460
rect 92873 255454 93193 255486
rect 92873 255218 92915 255454
rect 93151 255218 93193 255454
rect 92873 255134 93193 255218
rect 92873 254898 92915 255134
rect 93151 254898 93193 255134
rect 92873 254866 93193 254898
rect 91507 241772 91573 241773
rect 91507 241708 91508 241772
rect 91572 241708 91573 241772
rect 91507 241707 91573 241708
rect 93531 240140 93597 240141
rect 93531 240076 93532 240140
rect 93596 240076 93597 240140
rect 93531 240075 93597 240076
rect 91139 238644 91205 238645
rect 91139 238580 91140 238644
rect 91204 238580 91205 238644
rect 91139 238579 91205 238580
rect 91794 237454 92414 239592
rect 91507 237420 91573 237421
rect 91507 237356 91508 237420
rect 91572 237356 91573 237420
rect 91507 237355 91573 237356
rect 89851 144804 89917 144805
rect 89851 144740 89852 144804
rect 89916 144740 89917 144804
rect 89851 144739 89917 144740
rect 87091 137596 87157 137597
rect 87091 137532 87092 137596
rect 87156 137532 87157 137596
rect 87091 137531 87157 137532
rect 91510 136370 91570 237355
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 93534 213213 93594 240075
rect 92979 213212 93045 213213
rect 92979 213148 92980 213212
rect 93044 213148 93045 213212
rect 92979 213147 93045 213148
rect 93531 213212 93597 213213
rect 93531 213148 93532 213212
rect 93596 213148 93597 213212
rect 93531 213147 93597 213148
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 136782 92414 164898
rect 91510 136310 91754 136370
rect 77644 129454 77964 129486
rect 77644 129218 77686 129454
rect 77922 129218 77964 129454
rect 77644 129134 77964 129218
rect 77644 128898 77686 129134
rect 77922 128898 77964 129134
rect 77644 128866 77964 128898
rect 85575 129454 85895 129486
rect 85575 129218 85617 129454
rect 85853 129218 85895 129454
rect 85575 129134 85895 129218
rect 85575 128898 85617 129134
rect 85853 128898 85895 129134
rect 85575 128866 85895 128898
rect 73679 111454 73999 111486
rect 73679 111218 73721 111454
rect 73957 111218 73999 111454
rect 73679 111134 73999 111218
rect 73679 110898 73721 111134
rect 73957 110898 73999 111134
rect 73679 110866 73999 110898
rect 81609 111454 81929 111486
rect 81609 111218 81651 111454
rect 81887 111218 81929 111454
rect 81609 111134 81929 111218
rect 81609 110898 81651 111134
rect 81887 110898 81929 111134
rect 81609 110866 81929 110898
rect 89540 111454 89860 111486
rect 89540 111218 89582 111454
rect 89818 111218 89860 111454
rect 89540 111134 89860 111218
rect 89540 110898 89582 111134
rect 89818 110898 89860 111134
rect 89540 110866 89860 110898
rect 91694 92445 91754 136310
rect 92982 92445 93042 213147
rect 93718 176765 93778 283459
rect 93899 237420 93965 237421
rect 93899 237356 93900 237420
rect 93964 237356 93965 237420
rect 93899 237355 93965 237356
rect 93715 176764 93781 176765
rect 93715 176700 93716 176764
rect 93780 176700 93781 176764
rect 93715 176699 93781 176700
rect 93902 113190 93962 237355
rect 94270 236605 94330 283459
rect 95371 282980 95437 282981
rect 95371 282916 95372 282980
rect 95436 282916 95437 282980
rect 95371 282915 95437 282916
rect 95374 238770 95434 282915
rect 95190 238710 95434 238770
rect 95190 236741 95250 238710
rect 95187 236740 95253 236741
rect 95187 236676 95188 236740
rect 95252 236676 95253 236740
rect 95187 236675 95253 236676
rect 94267 236604 94333 236605
rect 94267 236540 94268 236604
rect 94332 236540 94333 236604
rect 94267 236539 94333 236540
rect 94083 227764 94149 227765
rect 94083 227700 94084 227764
rect 94148 227700 94149 227764
rect 94083 227699 94149 227700
rect 94086 132510 94146 227699
rect 95514 205174 96134 239592
rect 96662 238509 96722 387771
rect 97950 308549 98010 433603
rect 98502 312493 98562 433739
rect 99971 433668 100037 433669
rect 99971 433604 99972 433668
rect 100036 433604 100037 433668
rect 99971 433603 100037 433604
rect 99234 352894 99854 388356
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 98499 312492 98565 312493
rect 98499 312428 98500 312492
rect 98564 312428 98565 312492
rect 98499 312427 98565 312428
rect 97947 308548 98013 308549
rect 97947 308484 97948 308548
rect 98012 308484 98013 308548
rect 97947 308483 98013 308484
rect 99234 285592 99854 316338
rect 99974 287741 100034 433603
rect 100158 390965 100218 434283
rect 100707 433668 100773 433669
rect 100707 433604 100708 433668
rect 100772 433604 100773 433668
rect 100707 433603 100773 433604
rect 100155 390964 100221 390965
rect 100155 390900 100156 390964
rect 100220 390900 100221 390964
rect 100155 390899 100221 390900
rect 100710 385797 100770 433603
rect 101262 388653 101322 549339
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 104939 551988 105005 551989
rect 104939 551924 104940 551988
rect 105004 551924 105005 551988
rect 104939 551923 105005 551924
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 436356 103574 464058
rect 104203 462908 104269 462909
rect 104203 462844 104204 462908
rect 104268 462844 104269 462908
rect 104203 462843 104269 462844
rect 102731 434620 102797 434621
rect 102731 434556 102732 434620
rect 102796 434556 102797 434620
rect 102731 434555 102797 434556
rect 101259 388652 101325 388653
rect 101259 388588 101260 388652
rect 101324 388588 101325 388652
rect 101259 388587 101325 388588
rect 100707 385796 100773 385797
rect 100707 385732 100708 385796
rect 100772 385732 100773 385796
rect 100707 385731 100773 385732
rect 102734 382941 102794 434555
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 104206 390965 104266 462843
rect 104942 390965 105002 551923
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 111747 530636 111813 530637
rect 111747 530572 111748 530636
rect 111812 530572 111813 530636
rect 111747 530571 111813 530572
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 436356 110414 470898
rect 106043 436116 106109 436117
rect 106043 436052 106044 436116
rect 106108 436052 106109 436116
rect 106043 436051 106109 436052
rect 104203 390964 104269 390965
rect 104203 390900 104204 390964
rect 104268 390900 104269 390964
rect 104203 390899 104269 390900
rect 104939 390964 105005 390965
rect 104939 390900 104940 390964
rect 105004 390900 105005 390964
rect 104939 390899 105005 390900
rect 102731 382940 102797 382941
rect 102731 382876 102732 382940
rect 102796 382876 102797 382940
rect 102731 382875 102797 382876
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 106046 320653 106106 436051
rect 106411 433668 106477 433669
rect 106411 433604 106412 433668
rect 106476 433604 106477 433668
rect 106411 433603 106477 433604
rect 109539 433668 109605 433669
rect 109539 433604 109540 433668
rect 109604 433604 109605 433668
rect 109539 433603 109605 433604
rect 111011 433668 111077 433669
rect 111011 433604 111012 433668
rect 111076 433604 111077 433668
rect 111011 433603 111077 433604
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 104939 320652 105005 320653
rect 104939 320588 104940 320652
rect 105004 320588 105005 320652
rect 104939 320587 105005 320588
rect 106043 320652 106109 320653
rect 106043 320588 106044 320652
rect 106108 320588 106109 320652
rect 106043 320587 106109 320588
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 99971 287740 100037 287741
rect 99971 287676 99972 287740
rect 100036 287676 100037 287740
rect 99971 287675 100037 287676
rect 102954 284614 103574 320058
rect 104942 313989 105002 320587
rect 104939 313988 105005 313989
rect 104939 313924 104940 313988
rect 105004 313924 105005 313988
rect 104939 313923 105005 313924
rect 106414 311133 106474 433603
rect 109542 315349 109602 433603
rect 109794 363454 110414 388356
rect 111014 370701 111074 433603
rect 111750 422310 111810 530571
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 112299 454748 112365 454749
rect 112299 454684 112300 454748
rect 112364 454684 112365 454748
rect 112299 454683 112365 454684
rect 112302 422310 112362 454683
rect 113514 439174 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 114323 457468 114389 457469
rect 114323 457404 114324 457468
rect 114388 457404 114389 457468
rect 114323 457403 114389 457404
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 436356 114134 438618
rect 113219 428228 113285 428229
rect 113219 428164 113220 428228
rect 113284 428164 113285 428228
rect 113219 428163 113285 428164
rect 111750 422250 112178 422310
rect 112302 422250 112914 422310
rect 112118 402661 112178 422250
rect 112854 402990 112914 422250
rect 112854 402930 113098 402990
rect 112115 402660 112181 402661
rect 112115 402596 112116 402660
rect 112180 402596 112181 402660
rect 112115 402595 112181 402596
rect 113038 400213 113098 402930
rect 113035 400212 113101 400213
rect 113035 400148 113036 400212
rect 113100 400148 113101 400212
rect 113035 400147 113101 400148
rect 112851 393956 112917 393957
rect 112851 393892 112852 393956
rect 112916 393892 112917 393956
rect 112851 393891 112917 393892
rect 111931 391644 111997 391645
rect 111931 391580 111932 391644
rect 111996 391580 111997 391644
rect 111931 391579 111997 391580
rect 111934 390965 111994 391579
rect 111931 390964 111997 390965
rect 111931 390900 111932 390964
rect 111996 390900 111997 390964
rect 111931 390899 111997 390900
rect 112854 390557 112914 393891
rect 113038 391645 113098 400147
rect 113035 391644 113101 391645
rect 113035 391580 113036 391644
rect 113100 391580 113101 391644
rect 113035 391579 113101 391580
rect 112851 390556 112917 390557
rect 112851 390492 112852 390556
rect 112916 390492 112917 390556
rect 112851 390491 112917 390492
rect 111011 370700 111077 370701
rect 111011 370636 111012 370700
rect 111076 370636 111077 370700
rect 111011 370635 111077 370636
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109539 315348 109605 315349
rect 109539 315284 109540 315348
rect 109604 315284 109605 315348
rect 109539 315283 109605 315284
rect 106411 311132 106477 311133
rect 106411 311068 106412 311132
rect 106476 311068 106477 311132
rect 106411 311067 106477 311068
rect 109542 307053 109602 315283
rect 109539 307052 109605 307053
rect 109539 306988 109540 307052
rect 109604 306988 109605 307052
rect 109539 306987 109605 306988
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 98867 283252 98933 283253
rect 98867 283188 98868 283252
rect 98932 283188 98933 283252
rect 98867 283187 98933 283188
rect 98870 268429 98930 283187
rect 99971 280260 100037 280261
rect 99971 280196 99972 280260
rect 100036 280196 100037 280260
rect 99971 280195 100037 280196
rect 98867 268428 98933 268429
rect 98867 268364 98868 268428
rect 98932 268364 98933 268428
rect 98867 268363 98933 268364
rect 98315 251292 98381 251293
rect 98315 251228 98316 251292
rect 98380 251228 98381 251292
rect 98315 251227 98381 251228
rect 98131 247212 98197 247213
rect 98131 247210 98132 247212
rect 97950 247150 98132 247210
rect 97763 240140 97829 240141
rect 97763 240076 97764 240140
rect 97828 240076 97829 240140
rect 97763 240075 97829 240076
rect 96659 238508 96725 238509
rect 96659 238444 96660 238508
rect 96724 238444 96725 238508
rect 96659 238443 96725 238444
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 97766 204373 97826 240075
rect 97950 214573 98010 247150
rect 98131 247148 98132 247150
rect 98196 247148 98197 247212
rect 98131 247147 98197 247148
rect 98318 238770 98378 251227
rect 98134 238710 98378 238770
rect 98134 220965 98194 238710
rect 98131 220964 98197 220965
rect 98131 220900 98132 220964
rect 98196 220900 98197 220964
rect 98131 220899 98197 220900
rect 98134 219450 98194 220899
rect 98134 219390 98562 219450
rect 97947 214572 98013 214573
rect 97947 214508 97948 214572
rect 98012 214508 98013 214572
rect 97947 214507 98013 214508
rect 97763 204372 97829 204373
rect 97763 204308 97764 204372
rect 97828 204308 97829 204372
rect 97763 204307 97829 204308
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95187 163436 95253 163437
rect 95187 163372 95188 163436
rect 95252 163372 95253 163436
rect 95187 163371 95253 163372
rect 94086 132450 94330 132510
rect 93902 113130 94146 113190
rect 94086 109173 94146 113130
rect 94083 109172 94149 109173
rect 94083 109108 94084 109172
rect 94148 109108 94149 109172
rect 94083 109107 94149 109108
rect 94270 106181 94330 132450
rect 94267 106180 94333 106181
rect 94267 106116 94268 106180
rect 94332 106116 94333 106180
rect 94267 106115 94333 106116
rect 94819 95844 94885 95845
rect 94819 95780 94820 95844
rect 94884 95780 94885 95844
rect 94819 95779 94885 95780
rect 91691 92444 91757 92445
rect 91691 92380 91692 92444
rect 91756 92380 91757 92444
rect 91691 92379 91757 92380
rect 92979 92444 93045 92445
rect 92979 92380 92980 92444
rect 93044 92380 93045 92444
rect 92979 92379 93045 92380
rect 72923 92308 72989 92309
rect 72923 92244 72924 92308
rect 72988 92244 72989 92308
rect 72923 92243 72989 92244
rect 94822 92037 94882 95779
rect 94819 92036 94885 92037
rect 94819 91972 94820 92036
rect 94884 91972 94885 92036
rect 94819 91971 94885 91972
rect 70163 89588 70229 89589
rect 70163 89524 70164 89588
rect 70228 89524 70229 89588
rect 70163 89523 70229 89524
rect 69611 84012 69677 84013
rect 69611 83948 69612 84012
rect 69676 83948 69677 84012
rect 69611 83947 69677 83948
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 90782
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 90782
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 90782
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 90782
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 90782
rect 95190 89861 95250 163371
rect 95514 136782 96134 168618
rect 98502 105093 98562 219390
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99974 144805 100034 280195
rect 100707 278764 100773 278765
rect 100707 278700 100708 278764
rect 100772 278700 100773 278764
rect 100707 278699 100773 278700
rect 100710 277813 100770 278699
rect 100707 277812 100773 277813
rect 100707 277748 100708 277812
rect 100772 277748 100773 277812
rect 100707 277747 100773 277748
rect 99971 144804 100037 144805
rect 99971 144740 99972 144804
rect 100036 144740 100037 144804
rect 99971 144739 100037 144740
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 98499 105092 98565 105093
rect 98499 105028 98500 105092
rect 98564 105028 98565 105092
rect 98499 105027 98565 105028
rect 99234 100894 99854 136338
rect 100710 129301 100770 277747
rect 101259 251156 101325 251157
rect 101259 251092 101260 251156
rect 101324 251092 101325 251156
rect 101259 251091 101325 251092
rect 101262 227765 101322 251091
rect 102954 248614 103574 284058
rect 109794 291454 110414 326898
rect 113222 304197 113282 428163
rect 114326 396405 114386 457403
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 114507 427140 114573 427141
rect 114507 427076 114508 427140
rect 114572 427076 114573 427140
rect 114507 427075 114573 427076
rect 114323 396404 114389 396405
rect 114323 396340 114324 396404
rect 114388 396340 114389 396404
rect 114323 396339 114389 396340
rect 114510 391509 114570 427075
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 114507 391508 114573 391509
rect 114507 391444 114508 391508
rect 114572 391444 114573 391508
rect 114507 391443 114573 391444
rect 113514 367174 114134 388356
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113219 304196 113285 304197
rect 113219 304132 113220 304196
rect 113284 304132 113285 304196
rect 113219 304131 113285 304132
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 105491 261492 105557 261493
rect 105491 261428 105492 261492
rect 105556 261428 105557 261492
rect 105491 261427 105557 261428
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 101259 227764 101325 227765
rect 101259 227700 101260 227764
rect 101324 227700 101325 227764
rect 101259 227699 101325 227700
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 104019 192540 104085 192541
rect 104019 192476 104020 192540
rect 104084 192476 104085 192540
rect 104019 192475 104085 192476
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 100707 129300 100773 129301
rect 100707 129236 100708 129300
rect 100772 129236 100773 129300
rect 100707 129235 100773 129236
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 97211 96116 97277 96117
rect 97211 96052 97212 96116
rect 97276 96052 97277 96116
rect 97211 96051 97277 96052
rect 95187 89860 95253 89861
rect 95187 89796 95188 89860
rect 95252 89796 95253 89860
rect 95187 89795 95253 89796
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 90782
rect 97214 75853 97274 96051
rect 97211 75852 97277 75853
rect 97211 75788 97212 75852
rect 97276 75788 97277 75852
rect 97211 75787 97277 75788
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 104022 103597 104082 192475
rect 104019 103596 104085 103597
rect 104019 103532 104020 103596
rect 104084 103532 104085 103596
rect 104019 103531 104085 103532
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 105494 55861 105554 261427
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 106779 119372 106845 119373
rect 106779 119308 106780 119372
rect 106844 119308 106845 119372
rect 106779 119307 106845 119308
rect 105491 55860 105557 55861
rect 105491 55796 105492 55860
rect 105556 55796 105557 55860
rect 105491 55795 105557 55796
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 106782 28253 106842 119307
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 106779 28252 106845 28253
rect 106779 28188 106780 28252
rect 106844 28188 106845 28252
rect 106779 28187 106845 28188
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 124811 349756 124877 349757
rect 124811 349692 124812 349756
rect 124876 349692 124877 349756
rect 124811 349691 124877 349692
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 124814 15877 124874 349691
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 124811 15876 124877 15877
rect 124811 15812 124812 15876
rect 124876 15812 124877 15876
rect 124811 15811 124877 15812
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 148179 554844 148245 554845
rect 148179 554780 148180 554844
rect 148244 554780 148245 554844
rect 148179 554779 148245 554780
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 148182 433261 148242 554779
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 154435 600948 154501 600949
rect 154435 600884 154436 600948
rect 154500 600884 154501 600948
rect 154435 600883 154501 600884
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 150939 503028 151005 503029
rect 150939 502964 150940 503028
rect 151004 502964 151005 503028
rect 150939 502963 151005 502964
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 148179 433260 148245 433261
rect 148179 433196 148180 433260
rect 148244 433196 148245 433260
rect 148179 433195 148245 433196
rect 148179 429316 148245 429317
rect 148179 429252 148180 429316
rect 148244 429252 148245 429316
rect 148179 429251 148245 429252
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 144131 336836 144197 336837
rect 144131 336772 144132 336836
rect 144196 336772 144197 336836
rect 144131 336771 144197 336772
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 141371 264212 141437 264213
rect 141371 264148 141372 264212
rect 141436 264148 141437 264212
rect 141371 264147 141437 264148
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 141374 44845 141434 264147
rect 141371 44844 141437 44845
rect 141371 44780 141372 44844
rect 141436 44780 141437 44844
rect 141371 44779 141437 44780
rect 144134 43485 144194 336771
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 148182 310453 148242 429251
rect 149514 403174 150134 438618
rect 150942 413949 151002 502963
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 150939 413948 151005 413949
rect 150939 413884 150940 413948
rect 151004 413884 151005 413948
rect 150939 413883 151005 413884
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 148179 310452 148245 310453
rect 148179 310388 148180 310452
rect 148244 310388 148245 310452
rect 148179 310387 148245 310388
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 144131 43484 144197 43485
rect 144131 43420 144132 43484
rect 144196 43420 144197 43484
rect 144131 43419 144197 43420
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 154438 297397 154498 600883
rect 156954 590614 157574 626058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 162715 619716 162781 619717
rect 162715 619652 162716 619716
rect 162780 619652 162781 619716
rect 162715 619651 162781 619652
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156643 578916 156709 578917
rect 156643 578852 156644 578916
rect 156708 578852 156709 578916
rect 156643 578851 156709 578852
rect 155723 419660 155789 419661
rect 155723 419596 155724 419660
rect 155788 419596 155789 419660
rect 155723 419595 155789 419596
rect 154435 297396 154501 297397
rect 154435 297332 154436 297396
rect 154500 297332 154501 297396
rect 154435 297331 154501 297332
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 155726 250477 155786 419595
rect 156646 306373 156706 578851
rect 156954 554614 157574 590058
rect 159771 588028 159837 588029
rect 159771 587964 159772 588028
rect 159836 587964 159837 588028
rect 159771 587963 159837 587964
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 158483 552260 158549 552261
rect 158483 552196 158484 552260
rect 158548 552196 158549 552260
rect 158483 552195 158549 552196
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 158486 338061 158546 552195
rect 159774 349893 159834 587963
rect 161243 539612 161309 539613
rect 161243 539548 161244 539612
rect 161308 539548 161309 539612
rect 161243 539547 161309 539548
rect 159955 523700 160021 523701
rect 159955 523636 159956 523700
rect 160020 523636 160021 523700
rect 159955 523635 160021 523636
rect 159771 349892 159837 349893
rect 159771 349828 159772 349892
rect 159836 349828 159837 349892
rect 159771 349827 159837 349828
rect 156643 306372 156709 306373
rect 156643 306308 156644 306372
rect 156708 306308 156709 306372
rect 156643 306307 156709 306308
rect 156646 300117 156706 306307
rect 156954 302614 157574 338058
rect 158483 338060 158549 338061
rect 158483 337996 158484 338060
rect 158548 337996 158549 338060
rect 158483 337995 158549 337996
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156643 300116 156709 300117
rect 156643 300052 156644 300116
rect 156708 300052 156709 300116
rect 156643 300051 156709 300052
rect 156954 266614 157574 302058
rect 159771 301612 159837 301613
rect 159771 301548 159772 301612
rect 159836 301548 159837 301612
rect 159771 301547 159837 301548
rect 159774 282981 159834 301547
rect 159771 282980 159837 282981
rect 159771 282916 159772 282980
rect 159836 282916 159837 282980
rect 159771 282915 159837 282916
rect 159958 267069 160018 523635
rect 161059 497452 161125 497453
rect 161059 497388 161060 497452
rect 161124 497388 161125 497452
rect 161059 497387 161125 497388
rect 161062 371925 161122 497387
rect 161059 371924 161125 371925
rect 161059 371860 161060 371924
rect 161124 371860 161125 371924
rect 161059 371859 161125 371860
rect 161246 317661 161306 539547
rect 162531 468484 162597 468485
rect 162531 468420 162532 468484
rect 162596 468420 162597 468484
rect 162531 468419 162597 468420
rect 162534 321605 162594 468419
rect 162718 401709 162778 619651
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 166763 565860 166829 565861
rect 166763 565796 166764 565860
rect 166828 565796 166829 565860
rect 166763 565795 166829 565796
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 166211 512684 166277 512685
rect 166211 512620 166212 512684
rect 166276 512620 166277 512684
rect 166211 512619 166277 512620
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163451 438156 163517 438157
rect 163451 438092 163452 438156
rect 163516 438092 163517 438156
rect 163451 438091 163517 438092
rect 162715 401708 162781 401709
rect 162715 401644 162716 401708
rect 162780 401644 162781 401708
rect 162715 401643 162781 401644
rect 162715 401572 162781 401573
rect 162715 401508 162716 401572
rect 162780 401508 162781 401572
rect 162715 401507 162781 401508
rect 162531 321604 162597 321605
rect 162531 321540 162532 321604
rect 162596 321540 162597 321604
rect 162531 321539 162597 321540
rect 160691 317660 160757 317661
rect 160691 317596 160692 317660
rect 160756 317596 160757 317660
rect 160691 317595 160757 317596
rect 161243 317660 161309 317661
rect 161243 317596 161244 317660
rect 161308 317596 161309 317660
rect 161243 317595 161309 317596
rect 160694 291821 160754 317595
rect 160691 291820 160757 291821
rect 160691 291756 160692 291820
rect 160756 291756 160757 291820
rect 160691 291755 160757 291756
rect 160691 276724 160757 276725
rect 160691 276660 160692 276724
rect 160756 276660 160757 276724
rect 160691 276659 160757 276660
rect 159955 267068 160021 267069
rect 159955 267004 159956 267068
rect 160020 267004 160021 267068
rect 159955 267003 160021 267004
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 159958 266389 160018 267003
rect 156954 266294 157574 266378
rect 159955 266388 160021 266389
rect 159955 266324 159956 266388
rect 160020 266324 160021 266388
rect 159955 266323 160021 266324
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 155723 250476 155789 250477
rect 155723 250412 155724 250476
rect 155788 250412 155789 250476
rect 155723 250411 155789 250412
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 230614 157574 266058
rect 160694 233205 160754 276659
rect 162718 269109 162778 401507
rect 162715 269108 162781 269109
rect 162715 269044 162716 269108
rect 162780 269044 162781 269108
rect 162715 269043 162781 269044
rect 163454 251973 163514 438091
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 166214 301749 166274 512619
rect 166766 346493 166826 565795
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 180011 610060 180077 610061
rect 180011 609996 180012 610060
rect 180076 609996 180077 610060
rect 180011 609995 180077 609996
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 178539 572796 178605 572797
rect 178539 572732 178540 572796
rect 178604 572732 178605 572796
rect 178539 572731 178605 572732
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 171234 568574 171854 568658
rect 172099 568716 172165 568717
rect 172099 568652 172100 568716
rect 172164 568652 172165 568716
rect 172099 568651 172165 568652
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 170811 560420 170877 560421
rect 170811 560356 170812 560420
rect 170876 560356 170877 560420
rect 170811 560355 170877 560356
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 168971 486572 169037 486573
rect 168971 486508 168972 486572
rect 169036 486508 169037 486572
rect 168971 486507 169037 486508
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 166763 346492 166829 346493
rect 166763 346428 166764 346492
rect 166828 346428 166829 346492
rect 166763 346427 166829 346428
rect 166395 321604 166461 321605
rect 166395 321540 166396 321604
rect 166460 321540 166461 321604
rect 166395 321539 166461 321540
rect 166211 301748 166277 301749
rect 166211 301684 166212 301748
rect 166276 301684 166277 301748
rect 166211 301683 166277 301684
rect 166211 291820 166277 291821
rect 166211 291756 166212 291820
rect 166276 291756 166277 291820
rect 166211 291755 166277 291756
rect 166214 276725 166274 291755
rect 166211 276724 166277 276725
rect 166211 276660 166212 276724
rect 166276 276660 166277 276724
rect 166211 276659 166277 276660
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163451 251972 163517 251973
rect 163451 251908 163452 251972
rect 163516 251908 163517 251972
rect 163451 251907 163517 251908
rect 163794 237454 164414 272898
rect 166398 264893 166458 321539
rect 167514 313174 168134 348618
rect 168974 333301 169034 486507
rect 170814 427141 170874 560355
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 170995 465900 171061 465901
rect 170995 465836 170996 465900
rect 171060 465836 171061 465900
rect 170995 465835 171061 465836
rect 170811 427140 170877 427141
rect 170811 427076 170812 427140
rect 170876 427076 170877 427140
rect 170811 427075 170877 427076
rect 169707 388788 169773 388789
rect 169707 388724 169708 388788
rect 169772 388724 169773 388788
rect 169707 388723 169773 388724
rect 169710 386341 169770 388723
rect 169707 386340 169773 386341
rect 169707 386276 169708 386340
rect 169772 386276 169773 386340
rect 169707 386275 169773 386276
rect 170811 386340 170877 386341
rect 170811 386276 170812 386340
rect 170876 386276 170877 386340
rect 170811 386275 170877 386276
rect 168971 333300 169037 333301
rect 168971 333236 168972 333300
rect 169036 333236 169037 333300
rect 168971 333235 169037 333236
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 168419 297396 168485 297397
rect 168419 297332 168420 297396
rect 168484 297332 168485 297396
rect 168419 297331 168485 297332
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 166395 264892 166461 264893
rect 166395 264828 166396 264892
rect 166460 264828 166461 264892
rect 166395 264827 166461 264828
rect 166763 248436 166829 248437
rect 166763 248372 166764 248436
rect 166828 248372 166829 248436
rect 166763 248371 166829 248372
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 160691 233204 160757 233205
rect 160691 233140 160692 233204
rect 160756 233140 160757 233204
rect 160691 233139 160757 233140
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 201454 164414 236898
rect 166766 209790 166826 248371
rect 166214 209730 166826 209790
rect 167514 241174 168134 276618
rect 168422 265573 168482 297331
rect 168419 265572 168485 265573
rect 168419 265508 168420 265572
rect 168484 265508 168485 265572
rect 168419 265507 168485 265508
rect 168235 260812 168301 260813
rect 168235 260748 168236 260812
rect 168300 260748 168301 260812
rect 168235 260747 168301 260748
rect 168238 259861 168298 260747
rect 168235 259860 168301 259861
rect 168235 259796 168236 259860
rect 168300 259796 168301 259860
rect 168235 259795 168301 259796
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 166214 205597 166274 209730
rect 166211 205596 166277 205597
rect 166211 205532 166212 205596
rect 166276 205532 166277 205596
rect 166211 205531 166277 205532
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 166214 30973 166274 205531
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 168238 72453 168298 259795
rect 170814 254285 170874 386275
rect 170998 327861 171058 465835
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 172102 423741 172162 568651
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 173571 471340 173637 471341
rect 173571 471276 173572 471340
rect 173636 471276 173637 471340
rect 173571 471275 173637 471276
rect 173574 453933 173634 471275
rect 173755 469300 173821 469301
rect 173755 469236 173756 469300
rect 173820 469236 173821 469300
rect 173755 469235 173821 469236
rect 173571 453932 173637 453933
rect 173571 453868 173572 453932
rect 173636 453868 173637 453932
rect 173571 453867 173637 453868
rect 173571 453796 173637 453797
rect 173571 453732 173572 453796
rect 173636 453732 173637 453796
rect 173571 453731 173637 453732
rect 172099 423740 172165 423741
rect 172099 423676 172100 423740
rect 172164 423676 172165 423740
rect 172099 423675 172165 423676
rect 172283 419660 172349 419661
rect 172283 419596 172284 419660
rect 172348 419596 172349 419660
rect 172283 419595 172349 419596
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 170995 327860 171061 327861
rect 170995 327796 170996 327860
rect 171060 327796 171061 327860
rect 170995 327795 171061 327796
rect 171234 316894 171854 352338
rect 172286 334797 172346 419595
rect 172283 334796 172349 334797
rect 172283 334732 172284 334796
rect 172348 334732 172349 334796
rect 172283 334731 172349 334732
rect 173574 327725 173634 453731
rect 173758 331941 173818 469235
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 176515 464404 176581 464405
rect 176515 464340 176516 464404
rect 176580 464340 176581 464404
rect 176515 464339 176581 464340
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 176518 444277 176578 464339
rect 177619 462908 177685 462909
rect 177619 462844 177620 462908
rect 177684 462844 177685 462908
rect 177619 462843 177685 462844
rect 176515 444276 176581 444277
rect 176515 444212 176516 444276
rect 176580 444212 176581 444276
rect 176515 444211 176581 444212
rect 176331 443596 176397 443597
rect 176331 443532 176332 443596
rect 176396 443532 176397 443596
rect 176331 443531 176397 443532
rect 176334 441630 176394 443531
rect 176334 441570 176578 441630
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 173755 331940 173821 331941
rect 173755 331876 173756 331940
rect 173820 331876 173821 331940
rect 173755 331875 173821 331876
rect 173571 327724 173637 327725
rect 173571 327660 173572 327724
rect 173636 327660 173637 327724
rect 173571 327659 173637 327660
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 173019 309364 173085 309365
rect 173019 309300 173020 309364
rect 173084 309300 173085 309364
rect 173019 309299 173085 309300
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 170811 254284 170877 254285
rect 170811 254220 170812 254284
rect 170876 254220 170877 254284
rect 170811 254219 170877 254220
rect 168419 251156 168485 251157
rect 168419 251092 168420 251156
rect 168484 251092 168485 251156
rect 168419 251091 168485 251092
rect 168422 188325 168482 251091
rect 171234 244894 171854 280338
rect 173022 258773 173082 309299
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 173019 258772 173085 258773
rect 173019 258708 173020 258772
rect 173084 258708 173085 258772
rect 173019 258707 173085 258708
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 168419 188324 168485 188325
rect 168419 188260 168420 188324
rect 168484 188260 168485 188324
rect 168419 188259 168485 188260
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 168235 72452 168301 72453
rect 168235 72388 168236 72452
rect 168300 72388 168301 72452
rect 168235 72387 168301 72388
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 166211 30972 166277 30973
rect 166211 30908 166212 30972
rect 166276 30908 166277 30972
rect 166211 30907 166277 30908
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 248614 175574 284058
rect 176518 267750 176578 441570
rect 177622 340917 177682 462843
rect 177803 449444 177869 449445
rect 177803 449380 177804 449444
rect 177868 449380 177869 449444
rect 177803 449379 177869 449380
rect 177619 340916 177685 340917
rect 177619 340852 177620 340916
rect 177684 340852 177685 340916
rect 177619 340851 177685 340852
rect 177619 340236 177685 340237
rect 177619 340172 177620 340236
rect 177684 340172 177685 340236
rect 177619 340171 177685 340172
rect 175782 267690 176578 267750
rect 175782 264213 175842 267690
rect 175779 264212 175845 264213
rect 175779 264148 175780 264212
rect 175844 264148 175845 264212
rect 175779 264147 175845 264148
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 175782 26893 175842 264147
rect 177622 253877 177682 340171
rect 177806 257277 177866 449379
rect 177987 337924 178053 337925
rect 177987 337860 177988 337924
rect 178052 337860 178053 337924
rect 177987 337859 178053 337860
rect 177990 262853 178050 337859
rect 178542 334661 178602 572731
rect 178723 476780 178789 476781
rect 178723 476716 178724 476780
rect 178788 476716 178789 476780
rect 178723 476715 178789 476716
rect 178726 337245 178786 476715
rect 180014 469301 180074 609995
rect 181794 579454 182414 614898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 184059 608836 184125 608837
rect 184059 608772 184060 608836
rect 184124 608772 184125 608836
rect 184059 608771 184125 608772
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 184062 515405 184122 608771
rect 185514 583174 186134 618618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 188291 596324 188357 596325
rect 188291 596260 188292 596324
rect 188356 596260 188357 596324
rect 188291 596259 188357 596260
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 186819 558244 186885 558245
rect 186819 558180 186820 558244
rect 186884 558180 186885 558244
rect 186819 558179 186885 558180
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 184059 515404 184125 515405
rect 184059 515340 184060 515404
rect 184124 515340 184125 515404
rect 184059 515339 184125 515340
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181483 471884 181549 471885
rect 181483 471820 181484 471884
rect 181548 471820 181549 471884
rect 181483 471819 181549 471820
rect 180011 469300 180077 469301
rect 180011 469236 180012 469300
rect 180076 469236 180077 469300
rect 180011 469235 180077 469236
rect 180563 456380 180629 456381
rect 180563 456316 180564 456380
rect 180628 456316 180629 456380
rect 180563 456315 180629 456316
rect 178723 337244 178789 337245
rect 178723 337180 178724 337244
rect 178788 337180 178789 337244
rect 178723 337179 178789 337180
rect 178539 334660 178605 334661
rect 178539 334596 178540 334660
rect 178604 334596 178605 334660
rect 178539 334595 178605 334596
rect 180566 304197 180626 456315
rect 181486 406333 181546 471819
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 184795 458828 184861 458829
rect 184795 458764 184796 458828
rect 184860 458764 184861 458828
rect 184795 458763 184861 458764
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181483 406332 181549 406333
rect 181483 406268 181484 406332
rect 181548 406268 181549 406332
rect 181483 406267 181549 406268
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 180747 393412 180813 393413
rect 180747 393348 180748 393412
rect 180812 393348 180813 393412
rect 180747 393347 180813 393348
rect 180750 393141 180810 393347
rect 180747 393140 180813 393141
rect 180747 393076 180748 393140
rect 180812 393076 180813 393140
rect 180747 393075 180813 393076
rect 180747 383892 180813 383893
rect 180747 383828 180748 383892
rect 180812 383828 180813 383892
rect 180747 383827 180813 383828
rect 180750 383670 180810 383827
rect 180750 383621 180994 383670
rect 180750 383620 180997 383621
rect 180750 383610 180932 383620
rect 180931 383556 180932 383610
rect 180996 383556 180997 383620
rect 180931 383555 180997 383556
rect 180747 374100 180813 374101
rect 180747 374036 180748 374100
rect 180812 374036 180813 374100
rect 180747 374035 180813 374036
rect 180750 373829 180810 374035
rect 180747 373828 180813 373829
rect 180747 373764 180748 373828
rect 180812 373764 180813 373828
rect 180747 373763 180813 373764
rect 180747 364444 180813 364445
rect 180747 364380 180748 364444
rect 180812 364380 180813 364444
rect 180747 364379 180813 364380
rect 180750 364173 180810 364379
rect 180747 364172 180813 364173
rect 180747 364108 180748 364172
rect 180812 364108 180813 364172
rect 180747 364107 180813 364108
rect 181794 363454 182414 398898
rect 184798 398037 184858 458763
rect 185514 439174 186134 474618
rect 186822 474197 186882 558179
rect 187555 475420 187621 475421
rect 187555 475356 187556 475420
rect 187620 475356 187621 475420
rect 187555 475355 187621 475356
rect 186819 474196 186885 474197
rect 186819 474132 186820 474196
rect 186884 474132 186885 474196
rect 186819 474131 186885 474132
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 184795 398036 184861 398037
rect 184795 397972 184796 398036
rect 184860 397972 184861 398036
rect 184795 397971 184861 397972
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 180747 354924 180813 354925
rect 180747 354860 180748 354924
rect 180812 354860 180813 354924
rect 180747 354859 180813 354860
rect 180750 354653 180810 354859
rect 180747 354652 180813 354653
rect 180747 354588 180748 354652
rect 180812 354588 180813 354652
rect 180747 354587 180813 354588
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 180563 304196 180629 304197
rect 180563 304132 180564 304196
rect 180628 304132 180629 304196
rect 180563 304131 180629 304132
rect 179275 302292 179341 302293
rect 179275 302228 179276 302292
rect 179340 302228 179341 302292
rect 179275 302227 179341 302228
rect 177987 262852 178053 262853
rect 177987 262788 177988 262852
rect 178052 262788 178053 262852
rect 177987 262787 178053 262788
rect 177803 257276 177869 257277
rect 177803 257212 177804 257276
rect 177868 257212 177869 257276
rect 177803 257211 177869 257212
rect 177619 253876 177685 253877
rect 177619 253812 177620 253876
rect 177684 253812 177685 253876
rect 177619 253811 177685 253812
rect 179278 251837 179338 302227
rect 181794 291454 182414 326898
rect 185514 367174 186134 402618
rect 187558 372741 187618 475355
rect 188294 417485 188354 596259
rect 189234 586894 189854 622338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192339 607340 192405 607341
rect 192339 607276 192340 607340
rect 192404 607276 192405 607340
rect 192339 607275 192405 607276
rect 192342 598229 192402 607275
rect 192954 601166 193574 626058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 601166 200414 632898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601166 204134 636618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 601166 207854 604338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 601166 211574 608058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 601166 218414 614898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 601166 222134 618618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 601166 225854 622338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 601166 229574 626058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 601166 236414 632898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601166 240134 636618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 601166 243854 604338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 244595 601900 244661 601901
rect 244595 601836 244596 601900
rect 244660 601836 244661 601900
rect 244595 601835 244661 601836
rect 219939 600812 220005 600813
rect 219939 600748 219940 600812
rect 220004 600748 220005 600812
rect 219939 600747 220005 600748
rect 193443 600540 193509 600541
rect 193443 600476 193444 600540
rect 193508 600476 193509 600540
rect 193443 600475 193509 600476
rect 193259 598500 193325 598501
rect 193259 598436 193260 598500
rect 193324 598436 193325 598500
rect 193259 598435 193325 598436
rect 192339 598228 192405 598229
rect 192339 598164 192340 598228
rect 192404 598164 192405 598228
rect 192339 598163 192405 598164
rect 193262 595509 193322 598435
rect 193446 596869 193506 600475
rect 215339 600404 215405 600405
rect 215339 600340 215340 600404
rect 215404 600340 215405 600404
rect 215339 600339 215405 600340
rect 218651 600404 218717 600405
rect 218651 600340 218652 600404
rect 218716 600340 218717 600404
rect 218651 600339 218717 600340
rect 212395 599452 212461 599453
rect 212395 599388 212396 599452
rect 212460 599388 212461 599452
rect 212395 599387 212461 599388
rect 204851 599180 204917 599181
rect 204851 599116 204852 599180
rect 204916 599116 204917 599180
rect 204851 599115 204917 599116
rect 194547 599044 194613 599045
rect 194547 598980 194548 599044
rect 194612 598980 194613 599044
rect 194547 598979 194613 598980
rect 197123 599044 197189 599045
rect 197123 598980 197124 599044
rect 197188 598980 197189 599044
rect 197123 598979 197189 598980
rect 201539 599044 201605 599045
rect 201539 598980 201540 599044
rect 201604 598980 201605 599044
rect 201539 598979 201605 598980
rect 203011 599044 203077 599045
rect 203011 598980 203012 599044
rect 203076 598980 203077 599044
rect 203011 598979 203077 598980
rect 193443 596868 193509 596869
rect 193443 596804 193444 596868
rect 193508 596804 193509 596868
rect 193443 596803 193509 596804
rect 193259 595508 193325 595509
rect 193259 595444 193260 595508
rect 193324 595444 193325 595508
rect 193259 595443 193325 595444
rect 193811 590204 193877 590205
rect 193811 590140 193812 590204
rect 193876 590140 193877 590204
rect 193811 590139 193877 590140
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 188475 542468 188541 542469
rect 188475 542404 188476 542468
rect 188540 542404 188541 542468
rect 188475 542403 188541 542404
rect 188478 498813 188538 542403
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 188475 498812 188541 498813
rect 188475 498748 188476 498812
rect 188540 498748 188541 498812
rect 188475 498747 188541 498748
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 188843 459100 188909 459101
rect 188843 459036 188844 459100
rect 188908 459036 188909 459100
rect 188843 459035 188909 459036
rect 188291 417484 188357 417485
rect 188291 417420 188292 417484
rect 188356 417420 188357 417484
rect 188291 417419 188357 417420
rect 188846 375461 188906 459035
rect 189234 442894 189854 478338
rect 192954 518614 193574 537166
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 190315 467124 190381 467125
rect 190315 467060 190316 467124
rect 190380 467060 190381 467124
rect 190315 467059 190381 467060
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 188843 375460 188909 375461
rect 188843 375396 188844 375460
rect 188908 375396 188909 375460
rect 188843 375395 188909 375396
rect 187555 372740 187621 372741
rect 187555 372676 187556 372740
rect 187620 372676 187621 372740
rect 187555 372675 187621 372676
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 184795 323644 184861 323645
rect 184795 323580 184796 323644
rect 184860 323580 184861 323644
rect 184795 323579 184861 323580
rect 184059 302564 184125 302565
rect 184059 302500 184060 302564
rect 184124 302500 184125 302564
rect 184059 302499 184125 302500
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 184062 278085 184122 302499
rect 184059 278084 184125 278085
rect 184059 278020 184060 278084
rect 184124 278020 184125 278084
rect 184059 278019 184125 278020
rect 184798 257413 184858 323579
rect 185347 306780 185413 306781
rect 185347 306716 185348 306780
rect 185412 306716 185413 306780
rect 185347 306715 185413 306716
rect 185350 291821 185410 306715
rect 185514 295174 186134 330618
rect 189234 370894 189854 406338
rect 190318 389877 190378 467059
rect 192954 452356 193574 482058
rect 193075 450396 193141 450397
rect 193075 450332 193076 450396
rect 193140 450332 193141 450396
rect 193075 450331 193141 450332
rect 191787 448492 191853 448493
rect 191787 448428 191788 448492
rect 191852 448428 191853 448492
rect 191787 448427 191853 448428
rect 190315 389876 190381 389877
rect 190315 389812 190316 389876
rect 190380 389812 190381 389876
rect 190315 389811 190381 389812
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 187555 314124 187621 314125
rect 187555 314060 187556 314124
rect 187620 314060 187621 314124
rect 187555 314059 187621 314060
rect 186819 303652 186885 303653
rect 186819 303588 186820 303652
rect 186884 303588 186885 303652
rect 186819 303587 186885 303588
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185347 291820 185413 291821
rect 185347 291756 185348 291820
rect 185412 291756 185413 291820
rect 185347 291755 185413 291756
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 184795 257412 184861 257413
rect 184795 257348 184796 257412
rect 184860 257348 184861 257412
rect 184795 257347 184861 257348
rect 184798 256733 184858 257347
rect 184795 256732 184861 256733
rect 184795 256668 184796 256732
rect 184860 256668 184861 256732
rect 184795 256667 184861 256668
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 179275 251836 179341 251837
rect 179275 251772 179276 251836
rect 179340 251772 179341 251836
rect 179275 251771 179341 251772
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 175779 26892 175845 26893
rect 175779 26828 175780 26892
rect 175844 26828 175845 26892
rect 175779 26827 175845 26828
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 186822 6221 186882 303587
rect 187558 258909 187618 314059
rect 188475 303788 188541 303789
rect 188475 303724 188476 303788
rect 188540 303724 188541 303788
rect 188475 303723 188541 303724
rect 188291 299844 188357 299845
rect 188291 299780 188292 299844
rect 188356 299780 188357 299844
rect 188291 299779 188357 299780
rect 187555 258908 187621 258909
rect 187555 258844 187556 258908
rect 187620 258844 187621 258908
rect 187555 258843 187621 258844
rect 187558 258093 187618 258843
rect 187555 258092 187621 258093
rect 187555 258028 187556 258092
rect 187620 258028 187621 258092
rect 187555 258027 187621 258028
rect 188294 185605 188354 299779
rect 188478 215933 188538 303723
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 191790 252653 191850 448427
rect 193078 446589 193138 450331
rect 193075 446588 193141 446589
rect 193075 446524 193076 446588
rect 193140 446524 193141 446588
rect 193075 446523 193141 446524
rect 191971 406332 192037 406333
rect 191971 406268 191972 406332
rect 192036 406268 192037 406332
rect 191971 406267 192037 406268
rect 191974 390693 192034 406267
rect 191971 390692 192037 390693
rect 191971 390628 191972 390692
rect 192036 390628 192037 390692
rect 191971 390627 192037 390628
rect 192954 374614 193574 388356
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 303592 193574 338058
rect 193814 275365 193874 590139
rect 194550 309093 194610 598979
rect 196019 535532 196085 535533
rect 196019 535468 196020 535532
rect 196084 535468 196085 535532
rect 196019 535467 196085 535468
rect 196022 314941 196082 535467
rect 197126 486437 197186 598979
rect 197776 579454 198096 579486
rect 197776 579218 197818 579454
rect 198054 579218 198096 579454
rect 197776 579134 198096 579218
rect 197776 578898 197818 579134
rect 198054 578898 198096 579134
rect 197776 578866 198096 578898
rect 197776 543454 198096 543486
rect 197776 543218 197818 543454
rect 198054 543218 198096 543454
rect 197776 543134 198096 543218
rect 197776 542898 197818 543134
rect 198054 542898 198096 543134
rect 197776 542866 198096 542898
rect 199794 525454 200414 537166
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 197123 486436 197189 486437
rect 197123 486372 197124 486436
rect 197188 486372 197189 486436
rect 197123 486371 197189 486372
rect 199794 453454 200414 488898
rect 201542 465901 201602 598979
rect 203014 467125 203074 598979
rect 203514 529174 204134 537166
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 204854 498813 204914 599115
rect 207059 599044 207125 599045
rect 207059 598980 207060 599044
rect 207124 598980 207125 599044
rect 207059 598979 207125 598980
rect 210739 599044 210805 599045
rect 210739 598980 210740 599044
rect 210804 598980 210805 599044
rect 210739 598979 210805 598980
rect 204851 498812 204917 498813
rect 204851 498748 204852 498812
rect 204916 498748 204917 498812
rect 204851 498747 204917 498748
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203011 467124 203077 467125
rect 203011 467060 203012 467124
rect 203076 467060 203077 467124
rect 203011 467059 203077 467060
rect 201539 465900 201605 465901
rect 201539 465836 201540 465900
rect 201604 465836 201605 465900
rect 201539 465835 201605 465836
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 452356 200414 452898
rect 203514 457174 204134 492618
rect 207062 462909 207122 598979
rect 207234 532894 207854 537166
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 210742 511325 210802 598979
rect 212398 586530 212458 599387
rect 211662 586470 212458 586530
rect 210954 536614 211574 537166
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210739 511324 210805 511325
rect 210739 511260 210740 511324
rect 210804 511260 210805 511324
rect 210739 511259 210805 511260
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207059 462908 207125 462909
rect 207059 462844 207060 462908
rect 207124 462844 207125 462908
rect 207059 462843 207125 462844
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 452356 204134 456618
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 452356 207854 460338
rect 210954 500614 211574 536058
rect 211662 511461 211722 586470
rect 213136 561454 213456 561486
rect 213136 561218 213178 561454
rect 213414 561218 213456 561454
rect 213136 561134 213456 561218
rect 213136 560898 213178 561134
rect 213414 560898 213456 561134
rect 213136 560866 213456 560898
rect 211659 511460 211725 511461
rect 211659 511396 211660 511460
rect 211724 511396 211725 511460
rect 211659 511395 211725 511396
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 215342 464541 215402 600339
rect 217794 507454 218414 537166
rect 218654 530773 218714 600339
rect 219571 599044 219637 599045
rect 219571 598980 219572 599044
rect 219636 598980 219637 599044
rect 219571 598979 219637 598980
rect 218651 530772 218717 530773
rect 218651 530708 218652 530772
rect 218716 530708 218717 530772
rect 218651 530707 218717 530708
rect 219574 522477 219634 598979
rect 219942 526421 220002 600747
rect 232451 600676 232517 600677
rect 232451 600612 232452 600676
rect 232516 600612 232517 600676
rect 232451 600611 232517 600612
rect 230979 600404 231045 600405
rect 230979 600340 230980 600404
rect 231044 600340 231045 600404
rect 230979 600339 231045 600340
rect 226379 599452 226445 599453
rect 226379 599388 226380 599452
rect 226444 599388 226445 599452
rect 226379 599387 226445 599388
rect 222699 599180 222765 599181
rect 222699 599116 222700 599180
rect 222764 599116 222765 599180
rect 222699 599115 222765 599116
rect 220859 599044 220925 599045
rect 220859 598980 220860 599044
rect 220924 598980 220925 599044
rect 220859 598979 220925 598980
rect 219939 526420 220005 526421
rect 219939 526356 219940 526420
rect 220004 526356 220005 526420
rect 219939 526355 220005 526356
rect 219571 522476 219637 522477
rect 219571 522412 219572 522476
rect 219636 522412 219637 522476
rect 219571 522411 219637 522412
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 220862 482221 220922 598979
rect 221514 511174 222134 537166
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 220859 482220 220925 482221
rect 220859 482156 220860 482220
rect 220924 482156 220925 482220
rect 220859 482155 220925 482156
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 215339 464540 215405 464541
rect 215339 464476 215340 464540
rect 215404 464476 215405 464540
rect 215339 464475 215405 464476
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 452356 211574 464058
rect 217794 452356 218414 470898
rect 221514 475174 222134 510618
rect 222702 505749 222762 599115
rect 223803 599044 223869 599045
rect 223803 598980 223804 599044
rect 223868 598980 223869 599044
rect 223803 598979 223869 598980
rect 223987 599044 224053 599045
rect 223987 598980 223988 599044
rect 224052 598980 224053 599044
rect 223987 598979 224053 598980
rect 222699 505748 222765 505749
rect 222699 505684 222700 505748
rect 222764 505684 222765 505748
rect 222699 505683 222765 505684
rect 223806 489973 223866 598979
rect 223803 489972 223869 489973
rect 223803 489908 223804 489972
rect 223868 489908 223869 489972
rect 223803 489907 223869 489908
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 452356 222134 474618
rect 223806 464405 223866 489907
rect 223990 465765 224050 598979
rect 225234 514894 225854 537166
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 226382 509829 226442 599387
rect 229691 599180 229757 599181
rect 229691 599116 229692 599180
rect 229756 599116 229757 599180
rect 229691 599115 229757 599116
rect 228219 599044 228285 599045
rect 228219 598980 228220 599044
rect 228284 598980 228285 599044
rect 228219 598979 228285 598980
rect 226379 509828 226445 509829
rect 226379 509764 226380 509828
rect 226444 509764 226445 509828
rect 226379 509763 226445 509764
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 223987 465764 224053 465765
rect 223987 465700 223988 465764
rect 224052 465700 224053 465764
rect 223987 465699 224053 465700
rect 223803 464404 223869 464405
rect 223803 464340 223804 464404
rect 223868 464340 223869 464404
rect 223803 464339 223869 464340
rect 225234 452356 225854 478338
rect 228222 456245 228282 598979
rect 228496 579454 228816 579486
rect 228496 579218 228538 579454
rect 228774 579218 228816 579454
rect 228496 579134 228816 579218
rect 228496 578898 228538 579134
rect 228774 578898 228816 579134
rect 228496 578866 228816 578898
rect 228496 543454 228816 543486
rect 228496 543218 228538 543454
rect 228774 543218 228816 543454
rect 228496 543134 228816 543218
rect 228496 542898 228538 543134
rect 228774 542898 228816 543134
rect 228496 542866 228816 542898
rect 228954 518614 229574 537166
rect 229694 522341 229754 599115
rect 230611 599044 230677 599045
rect 230611 598980 230612 599044
rect 230676 598980 230677 599044
rect 230611 598979 230677 598980
rect 230614 530773 230674 598979
rect 230611 530772 230677 530773
rect 230611 530708 230612 530772
rect 230676 530708 230677 530772
rect 230611 530707 230677 530708
rect 229691 522340 229757 522341
rect 229691 522276 229692 522340
rect 229756 522276 229757 522340
rect 229691 522275 229757 522276
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 230982 511461 231042 600339
rect 232454 518941 232514 600611
rect 238523 599452 238589 599453
rect 238523 599388 238524 599452
rect 238588 599388 238589 599452
rect 238523 599387 238589 599388
rect 237419 599180 237485 599181
rect 237419 599116 237420 599180
rect 237484 599116 237485 599180
rect 237419 599115 237485 599116
rect 233187 599044 233253 599045
rect 233187 598980 233188 599044
rect 233252 598980 233253 599044
rect 233187 598979 233253 598980
rect 234659 599044 234725 599045
rect 234659 598980 234660 599044
rect 234724 598980 234725 599044
rect 234659 598979 234725 598980
rect 236499 599044 236565 599045
rect 236499 598980 236500 599044
rect 236564 598980 236565 599044
rect 236499 598979 236565 598980
rect 232451 518940 232517 518941
rect 232451 518876 232452 518940
rect 232516 518876 232517 518940
rect 232451 518875 232517 518876
rect 230979 511460 231045 511461
rect 230979 511396 230980 511460
rect 231044 511396 231045 511460
rect 230979 511395 231045 511396
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228219 456244 228285 456245
rect 228219 456180 228220 456244
rect 228284 456180 228285 456244
rect 228219 456179 228285 456180
rect 228954 452356 229574 482058
rect 233190 459101 233250 598979
rect 233187 459100 233253 459101
rect 233187 459036 233188 459100
rect 233252 459036 233253 459100
rect 233187 459035 233253 459036
rect 234662 458965 234722 598979
rect 235794 525454 236414 537166
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 234659 458964 234725 458965
rect 234659 458900 234660 458964
rect 234724 458900 234725 458964
rect 234659 458899 234725 458900
rect 235794 453454 236414 488898
rect 236502 465901 236562 598979
rect 237422 483717 237482 599115
rect 238526 531997 238586 599387
rect 241651 599180 241717 599181
rect 241651 599116 241652 599180
rect 241716 599116 241717 599180
rect 241651 599115 241717 599116
rect 240731 599044 240797 599045
rect 240731 598980 240732 599044
rect 240796 598980 240797 599044
rect 240731 598979 240797 598980
rect 238523 531996 238589 531997
rect 238523 531932 238524 531996
rect 238588 531932 238589 531996
rect 238523 531931 238589 531932
rect 239514 529174 240134 537166
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 237419 483716 237485 483717
rect 237419 483652 237420 483716
rect 237484 483652 237485 483716
rect 237419 483651 237485 483652
rect 236499 465900 236565 465901
rect 236499 465836 236500 465900
rect 236564 465836 236565 465900
rect 236499 465835 236565 465836
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 452356 236414 452898
rect 239514 457174 240134 492618
rect 240734 481541 240794 598979
rect 240731 481540 240797 481541
rect 240731 481476 240732 481540
rect 240796 481476 240797 481540
rect 240731 481475 240797 481476
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 452356 240134 456618
rect 197776 435454 198096 435486
rect 197776 435218 197818 435454
rect 198054 435218 198096 435454
rect 197776 435134 198096 435218
rect 197776 434898 197818 435134
rect 198054 434898 198096 435134
rect 197776 434866 198096 434898
rect 228496 435454 228816 435486
rect 228496 435218 228538 435454
rect 228774 435218 228816 435454
rect 228496 435134 228816 435218
rect 228496 434898 228538 435134
rect 228774 434898 228816 435134
rect 228496 434866 228816 434898
rect 213136 417454 213456 417486
rect 213136 417218 213178 417454
rect 213414 417218 213456 417454
rect 213136 417134 213456 417218
rect 213136 416898 213178 417134
rect 213414 416898 213456 417134
rect 213136 416866 213456 416898
rect 197776 399454 198096 399486
rect 197776 399218 197818 399454
rect 198054 399218 198096 399454
rect 197776 399134 198096 399218
rect 197776 398898 197818 399134
rect 198054 398898 198096 399134
rect 197776 398866 198096 398898
rect 228496 399454 228816 399486
rect 228496 399218 228538 399454
rect 228774 399218 228816 399454
rect 228496 399134 228816 399218
rect 228496 398898 228538 399134
rect 228774 398898 228816 399134
rect 228496 398866 228816 398898
rect 199794 381454 200414 388356
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 196019 314940 196085 314941
rect 196019 314876 196020 314940
rect 196084 314876 196085 314940
rect 196019 314875 196085 314876
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 194547 309092 194613 309093
rect 194547 309028 194548 309092
rect 194612 309028 194613 309092
rect 194547 309027 194613 309028
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 303592 200414 308898
rect 203514 385174 204134 388356
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 303592 204134 312618
rect 207234 352894 207854 388356
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 303592 207854 316338
rect 210954 356614 211574 388356
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 303592 211574 320058
rect 217794 363454 218414 388356
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 303592 218414 326898
rect 221514 367174 222134 388356
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 303592 222134 330618
rect 225234 370894 225854 388356
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 303592 225854 334338
rect 228954 374614 229574 388356
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 303592 229574 338058
rect 235794 381454 236414 388356
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 303592 236414 308898
rect 239514 385174 240134 388356
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 241654 373421 241714 599115
rect 242939 599044 243005 599045
rect 242939 598980 242940 599044
rect 243004 598980 243005 599044
rect 242939 598979 243005 598980
rect 242942 382941 243002 598979
rect 243856 561454 244176 561486
rect 243856 561218 243898 561454
rect 244134 561218 244176 561454
rect 243856 561134 244176 561218
rect 243856 560898 243898 561134
rect 244134 560898 244176 561134
rect 243856 560866 244176 560898
rect 243234 532894 243854 537166
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 244411 515404 244477 515405
rect 244411 515340 244412 515404
rect 244476 515340 244477 515404
rect 244411 515339 244477 515340
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 452356 243854 460338
rect 243856 417454 244176 417486
rect 243856 417218 243898 417454
rect 244134 417218 244176 417454
rect 243856 417134 244176 417218
rect 243856 416898 243898 417134
rect 244134 416898 244176 417134
rect 243856 416866 244176 416898
rect 244227 389060 244293 389061
rect 244227 388996 244228 389060
rect 244292 389058 244293 389060
rect 244414 389058 244474 515339
rect 244598 496637 244658 601835
rect 246954 601166 247574 608058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 601166 254414 614898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 247723 599044 247789 599045
rect 247723 598980 247724 599044
rect 247788 598980 247789 599044
rect 247723 598979 247789 598980
rect 249931 599044 249997 599045
rect 249931 598980 249932 599044
rect 249996 598980 249997 599044
rect 249931 598979 249997 598980
rect 252507 599044 252573 599045
rect 252507 598980 252508 599044
rect 252572 598980 252573 599044
rect 252507 598979 252573 598980
rect 246954 536614 247574 537166
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 245699 511460 245765 511461
rect 245699 511396 245700 511460
rect 245764 511396 245765 511460
rect 245699 511395 245765 511396
rect 244595 496636 244661 496637
rect 244595 496572 244596 496636
rect 244660 496572 244661 496636
rect 244595 496571 244661 496572
rect 245702 449989 245762 511395
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 452356 247574 464058
rect 247726 456109 247786 598979
rect 248459 528596 248525 528597
rect 248459 528532 248460 528596
rect 248524 528532 248525 528596
rect 248459 528531 248525 528532
rect 247723 456108 247789 456109
rect 247723 456044 247724 456108
rect 247788 456044 247789 456108
rect 247723 456043 247789 456044
rect 247171 450668 247237 450669
rect 247171 450604 247172 450668
rect 247236 450604 247237 450668
rect 247171 450603 247237 450604
rect 245699 449988 245765 449989
rect 245699 449924 245700 449988
rect 245764 449924 245765 449988
rect 245699 449923 245765 449924
rect 244292 388998 244474 389058
rect 244292 388996 244293 388998
rect 244227 388995 244293 388996
rect 242939 382940 243005 382941
rect 242939 382876 242940 382940
rect 243004 382876 243005 382940
rect 242939 382875 243005 382876
rect 241651 373420 241717 373421
rect 241651 373356 241652 373420
rect 241716 373356 241717 373420
rect 241651 373355 241717 373356
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 303592 240134 312618
rect 243234 352894 243854 388356
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 244230 344317 244290 388995
rect 244227 344316 244293 344317
rect 244227 344252 244228 344316
rect 244292 344252 244293 344316
rect 244227 344251 244293 344252
rect 245702 339829 245762 449923
rect 247174 388517 247234 450603
rect 247723 449716 247789 449717
rect 247723 449652 247724 449716
rect 247788 449652 247789 449716
rect 247723 449651 247789 449652
rect 247171 388516 247237 388517
rect 247171 388452 247172 388516
rect 247236 388452 247237 388516
rect 247171 388451 247237 388452
rect 246954 356614 247574 388356
rect 247726 387021 247786 449651
rect 247723 387020 247789 387021
rect 247723 386956 247724 387020
rect 247788 386956 247789 387020
rect 247723 386955 247789 386956
rect 248462 370565 248522 528531
rect 249747 523700 249813 523701
rect 249747 523636 249748 523700
rect 249812 523636 249813 523700
rect 249747 523635 249813 523636
rect 249379 476236 249445 476237
rect 249379 476172 249380 476236
rect 249444 476172 249445 476236
rect 249379 476171 249445 476172
rect 249382 389061 249442 476171
rect 249750 389333 249810 523635
rect 249934 481813 249994 598979
rect 251219 539068 251285 539069
rect 251219 539004 251220 539068
rect 251284 539004 251285 539068
rect 251219 539003 251285 539004
rect 251222 489157 251282 539003
rect 252510 499590 252570 598979
rect 257514 583174 258134 618618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 258395 603124 258461 603125
rect 258395 603060 258396 603124
rect 258460 603060 258461 603124
rect 258395 603059 258461 603060
rect 258398 596190 258458 603059
rect 259499 601764 259565 601765
rect 259499 601700 259500 601764
rect 259564 601700 259565 601764
rect 259499 601699 259565 601700
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 255267 570620 255333 570621
rect 255267 570556 255268 570620
rect 255332 570556 255333 570620
rect 255267 570555 255333 570556
rect 253979 551784 254045 551785
rect 253979 551720 253980 551784
rect 254044 551720 254045 551784
rect 253979 551719 254045 551720
rect 253982 537437 254042 551719
rect 255270 539341 255330 570555
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 255267 539340 255333 539341
rect 255267 539276 255268 539340
rect 255332 539276 255333 539340
rect 255267 539275 255333 539276
rect 253979 537436 254045 537437
rect 253979 537372 253980 537436
rect 254044 537372 254045 537436
rect 253979 537371 254045 537372
rect 253059 509828 253125 509829
rect 253059 509764 253060 509828
rect 253124 509764 253125 509828
rect 253059 509763 253125 509764
rect 252510 499530 252754 499590
rect 251219 489156 251285 489157
rect 251219 489092 251220 489156
rect 251284 489092 251285 489156
rect 251219 489091 251285 489092
rect 252507 484396 252573 484397
rect 252507 484332 252508 484396
rect 252572 484332 252573 484396
rect 252507 484331 252573 484332
rect 249931 481812 249997 481813
rect 249931 481748 249932 481812
rect 249996 481748 249997 481812
rect 249931 481747 249997 481748
rect 249934 480270 249994 481747
rect 249934 480210 250362 480270
rect 250302 455429 250362 480210
rect 252510 460950 252570 484331
rect 252694 483853 252754 499530
rect 252691 483852 252757 483853
rect 252691 483788 252692 483852
rect 252756 483788 252757 483852
rect 252691 483787 252757 483788
rect 252510 460890 252938 460950
rect 250299 455428 250365 455429
rect 250299 455364 250300 455428
rect 250364 455364 250365 455428
rect 250299 455363 250365 455364
rect 252878 441013 252938 460890
rect 253062 446861 253122 509763
rect 253794 507454 254414 537166
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 254531 486436 254597 486437
rect 254531 486372 254532 486436
rect 254596 486372 254597 486436
rect 254531 486371 254597 486372
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 452356 254414 470898
rect 253979 448764 254045 448765
rect 253979 448700 253980 448764
rect 254044 448700 254045 448764
rect 253979 448699 254045 448700
rect 253059 446860 253125 446861
rect 253059 446796 253060 446860
rect 253124 446796 253125 446860
rect 253059 446795 253125 446796
rect 252875 441012 252941 441013
rect 252875 440948 252876 441012
rect 252940 440948 252941 441012
rect 252875 440947 252941 440948
rect 253982 430949 254042 448699
rect 254534 448629 254594 486371
rect 255270 466581 255330 539275
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 255267 466580 255333 466581
rect 255267 466516 255268 466580
rect 255332 466516 255333 466580
rect 255267 466515 255333 466516
rect 254531 448628 254597 448629
rect 254531 448564 254532 448628
rect 254596 448564 254597 448628
rect 254531 448563 254597 448564
rect 255270 437613 255330 466515
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 255267 437612 255333 437613
rect 255267 437548 255268 437612
rect 255332 437548 255333 437612
rect 255267 437547 255333 437548
rect 253059 430948 253125 430949
rect 253059 430884 253060 430948
rect 253124 430884 253125 430948
rect 253059 430883 253125 430884
rect 253979 430948 254045 430949
rect 253979 430884 253980 430948
rect 254044 430884 254045 430948
rect 253979 430883 254045 430884
rect 252875 396812 252941 396813
rect 252875 396748 252876 396812
rect 252940 396748 252941 396812
rect 252875 396747 252941 396748
rect 252878 393330 252938 396747
rect 252510 393270 252938 393330
rect 249747 389332 249813 389333
rect 249747 389268 249748 389332
rect 249812 389268 249813 389332
rect 249747 389267 249813 389268
rect 251035 389332 251101 389333
rect 251035 389268 251036 389332
rect 251100 389268 251101 389332
rect 251035 389267 251101 389268
rect 248643 389060 248709 389061
rect 248643 388996 248644 389060
rect 248708 388996 248709 389060
rect 248643 388995 248709 388996
rect 249379 389060 249445 389061
rect 249379 388996 249380 389060
rect 249444 388996 249445 389060
rect 249379 388995 249445 388996
rect 248459 370564 248525 370565
rect 248459 370500 248460 370564
rect 248524 370500 248525 370564
rect 248459 370499 248525 370500
rect 248646 369069 248706 388995
rect 248643 369068 248709 369069
rect 248643 369004 248644 369068
rect 248708 369004 248709 369068
rect 248643 369003 248709 369004
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 245699 339828 245765 339829
rect 245699 339764 245700 339828
rect 245764 339764 245765 339828
rect 245699 339763 245765 339764
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 303592 243854 316338
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 245699 305692 245765 305693
rect 245699 305628 245700 305692
rect 245764 305628 245765 305692
rect 245699 305627 245765 305628
rect 245702 300661 245762 305627
rect 246954 303592 247574 320058
rect 245699 300660 245765 300661
rect 245699 300596 245700 300660
rect 245764 300596 245765 300660
rect 245699 300595 245765 300596
rect 197776 291454 198096 291486
rect 197776 291218 197818 291454
rect 198054 291218 198096 291454
rect 197776 291134 198096 291218
rect 197776 290898 197818 291134
rect 198054 290898 198096 291134
rect 197776 290866 198096 290898
rect 228496 291454 228816 291486
rect 228496 291218 228538 291454
rect 228774 291218 228816 291454
rect 228496 291134 228816 291218
rect 228496 290898 228538 291134
rect 228774 290898 228816 291134
rect 228496 290866 228816 290898
rect 193811 275364 193877 275365
rect 193811 275300 193812 275364
rect 193876 275300 193877 275364
rect 193811 275299 193877 275300
rect 213136 273454 213456 273486
rect 213136 273218 213178 273454
rect 213414 273218 213456 273454
rect 213136 273134 213456 273218
rect 213136 272898 213178 273134
rect 213414 272898 213456 273134
rect 213136 272866 213456 272898
rect 243856 273454 244176 273486
rect 243856 273218 243898 273454
rect 244134 273218 244176 273454
rect 243856 273134 244176 273218
rect 243856 272898 243898 273134
rect 244134 272898 244176 273134
rect 243856 272866 244176 272898
rect 197776 255454 198096 255486
rect 197776 255218 197818 255454
rect 198054 255218 198096 255454
rect 197776 255134 198096 255218
rect 197776 254898 197818 255134
rect 198054 254898 198096 255134
rect 197776 254866 198096 254898
rect 228496 255454 228816 255486
rect 228496 255218 228538 255454
rect 228774 255218 228816 255454
rect 228496 255134 228816 255218
rect 228496 254898 228538 255134
rect 228774 254898 228816 255134
rect 228496 254866 228816 254898
rect 191787 252652 191853 252653
rect 191787 252588 191788 252652
rect 191852 252588 191853 252652
rect 191787 252587 191853 252588
rect 193995 252652 194061 252653
rect 193995 252588 193996 252652
rect 194060 252588 194061 252652
rect 193995 252587 194061 252588
rect 193443 249116 193509 249117
rect 193443 249052 193444 249116
rect 193508 249052 193509 249116
rect 193443 249051 193509 249052
rect 193446 248430 193506 249051
rect 193446 248370 193874 248430
rect 192339 247756 192405 247757
rect 192339 247692 192340 247756
rect 192404 247692 192405 247756
rect 192339 247691 192405 247692
rect 191787 247484 191853 247485
rect 191787 247420 191788 247484
rect 191852 247420 191853 247484
rect 191787 247419 191853 247420
rect 191790 240141 191850 247419
rect 191787 240140 191853 240141
rect 191787 240076 191788 240140
rect 191852 240076 191853 240140
rect 191787 240075 191853 240076
rect 192342 228853 192402 247691
rect 192954 230614 193574 239592
rect 193814 238645 193874 248370
rect 193998 240141 194058 252587
rect 251038 242045 251098 389267
rect 252510 360093 252570 393270
rect 252507 360092 252573 360093
rect 252507 360028 252508 360092
rect 252572 360028 252573 360092
rect 252507 360027 252573 360028
rect 253062 346357 253122 430883
rect 254531 415172 254597 415173
rect 254531 415108 254532 415172
rect 254596 415108 254597 415172
rect 254531 415107 254597 415108
rect 253794 363454 254414 388356
rect 254534 378725 254594 415107
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 254715 402660 254781 402661
rect 254715 402596 254716 402660
rect 254780 402596 254781 402660
rect 254715 402595 254781 402596
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 254718 392053 254778 402595
rect 254715 392052 254781 392053
rect 254715 391988 254716 392052
rect 254780 391988 254781 392052
rect 254715 391987 254781 391988
rect 254531 378724 254597 378725
rect 254531 378660 254532 378724
rect 254596 378660 254597 378724
rect 254531 378659 254597 378660
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253059 346356 253125 346357
rect 253059 346292 253060 346356
rect 253124 346292 253125 346356
rect 253059 346291 253125 346292
rect 253794 327454 254414 362898
rect 257514 367174 258134 402618
rect 258214 596130 258458 596190
rect 258214 377770 258274 596130
rect 258395 594828 258461 594829
rect 258395 594764 258396 594828
rect 258460 594764 258461 594828
rect 258395 594763 258461 594764
rect 258398 381717 258458 594763
rect 258395 381716 258461 381717
rect 258395 381652 258396 381716
rect 258460 381652 258461 381716
rect 258395 381651 258461 381652
rect 258214 377710 258458 377770
rect 258398 377365 258458 377710
rect 258395 377364 258461 377365
rect 258395 377300 258396 377364
rect 258460 377300 258461 377364
rect 258395 377299 258461 377300
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 259502 352613 259562 601699
rect 261234 586894 261854 622338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 263547 600540 263613 600541
rect 263547 600476 263548 600540
rect 263612 600476 263613 600540
rect 263547 600475 263613 600476
rect 262259 599180 262325 599181
rect 262259 599116 262260 599180
rect 262324 599116 262325 599180
rect 262259 599115 262325 599116
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 260971 563412 261037 563413
rect 260971 563348 260972 563412
rect 261036 563348 261037 563412
rect 260971 563347 261037 563348
rect 260974 373285 261034 563347
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 260971 373284 261037 373285
rect 260971 373220 260972 373284
rect 261036 373220 261037 373284
rect 260971 373219 261037 373220
rect 261234 370894 261854 406338
rect 262262 371925 262322 599115
rect 262443 478140 262509 478141
rect 262443 478076 262444 478140
rect 262508 478076 262509 478140
rect 262443 478075 262509 478076
rect 262259 371924 262325 371925
rect 262259 371860 262260 371924
rect 262324 371860 262325 371924
rect 262259 371859 262325 371860
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 259499 352612 259565 352613
rect 259499 352548 259500 352612
rect 259564 352548 259565 352612
rect 259499 352547 259565 352548
rect 261234 334894 261854 370338
rect 262259 349892 262325 349893
rect 262259 349828 262260 349892
rect 262324 349828 262325 349892
rect 262259 349827 262325 349828
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 258395 333300 258461 333301
rect 258395 333236 258396 333300
rect 258460 333236 258461 333300
rect 258395 333235 258461 333236
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 255267 329084 255333 329085
rect 255267 329020 255268 329084
rect 255332 329020 255333 329084
rect 255267 329019 255333 329020
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 303592 254414 326898
rect 251771 300932 251837 300933
rect 251771 300868 251772 300932
rect 251836 300868 251837 300932
rect 251771 300867 251837 300868
rect 197859 242044 197925 242045
rect 197859 241980 197860 242044
rect 197924 241980 197925 242044
rect 197859 241979 197925 241980
rect 242939 242044 243005 242045
rect 242939 241980 242940 242044
rect 243004 241980 243005 242044
rect 242939 241979 243005 241980
rect 251035 242044 251101 242045
rect 251035 241980 251036 242044
rect 251100 241980 251101 242044
rect 251035 241979 251101 241980
rect 193995 240140 194061 240141
rect 193995 240076 193996 240140
rect 194060 240076 194061 240140
rect 193995 240075 194061 240076
rect 193811 238644 193877 238645
rect 193811 238580 193812 238644
rect 193876 238580 193877 238644
rect 193811 238579 193877 238580
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192339 228852 192405 228853
rect 192339 228788 192340 228852
rect 192404 228788 192405 228852
rect 192339 228787 192405 228788
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188475 215932 188541 215933
rect 188475 215868 188476 215932
rect 188540 215868 188541 215932
rect 188475 215867 188541 215868
rect 188843 199340 188909 199341
rect 188843 199276 188844 199340
rect 188908 199276 188909 199340
rect 188843 199275 188909 199276
rect 188291 185604 188357 185605
rect 188291 185540 188292 185604
rect 188356 185540 188357 185604
rect 188291 185539 188357 185540
rect 188291 181388 188357 181389
rect 188291 181324 188292 181388
rect 188356 181324 188357 181388
rect 188291 181323 188357 181324
rect 188294 179485 188354 181323
rect 188291 179484 188357 179485
rect 188291 179420 188292 179484
rect 188356 179420 188357 179484
rect 188291 179419 188357 179420
rect 188294 131205 188354 179419
rect 188291 131204 188357 131205
rect 188291 131140 188292 131204
rect 188356 131140 188357 131204
rect 188291 131139 188357 131140
rect 188846 107813 188906 199275
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 190315 153780 190381 153781
rect 190315 153716 190316 153780
rect 190380 153716 190381 153780
rect 190315 153715 190381 153716
rect 190318 134605 190378 153715
rect 192954 143035 193574 158058
rect 193811 148340 193877 148341
rect 193811 148276 193812 148340
rect 193876 148276 193877 148340
rect 193811 148275 193877 148276
rect 193075 141132 193141 141133
rect 193075 141068 193076 141132
rect 193140 141068 193141 141132
rect 193075 141067 193141 141068
rect 193078 139093 193138 141067
rect 193075 139092 193141 139093
rect 193075 139028 193076 139092
rect 193140 139028 193141 139092
rect 193075 139027 193141 139028
rect 190315 134604 190381 134605
rect 190315 134540 190316 134604
rect 190380 134540 190381 134604
rect 190315 134539 190381 134540
rect 190318 132565 190378 134539
rect 190315 132564 190381 132565
rect 190315 132500 190316 132564
rect 190380 132500 190381 132564
rect 193814 132510 193874 148275
rect 197862 144805 197922 241979
rect 199794 237454 200414 239592
rect 201539 239460 201605 239461
rect 201539 239396 201540 239460
rect 201604 239396 201605 239460
rect 201539 239395 201605 239396
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 200619 180028 200685 180029
rect 200619 179964 200620 180028
rect 200684 179964 200685 180028
rect 200619 179963 200685 179964
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 197859 144804 197925 144805
rect 197859 144740 197860 144804
rect 197924 144740 197925 144804
rect 197859 144739 197925 144740
rect 199794 143035 200414 164898
rect 196571 142356 196637 142357
rect 196571 142292 196572 142356
rect 196636 142292 196637 142356
rect 196571 142291 196637 142292
rect 195099 140452 195165 140453
rect 195099 140388 195100 140452
rect 195164 140388 195165 140452
rect 195099 140387 195165 140388
rect 190315 132499 190381 132500
rect 193446 132450 193874 132510
rect 192707 132020 192773 132021
rect 192707 131956 192708 132020
rect 192772 131956 192773 132020
rect 192707 131955 192773 131956
rect 192710 131477 192770 131955
rect 193446 131477 193506 132450
rect 192707 131476 192773 131477
rect 192707 131412 192708 131476
rect 192772 131412 192773 131476
rect 192707 131411 192773 131412
rect 193443 131476 193509 131477
rect 193443 131412 193444 131476
rect 193508 131412 193509 131476
rect 193443 131411 193509 131412
rect 192339 123860 192405 123861
rect 192339 123796 192340 123860
rect 192404 123796 192405 123860
rect 192339 123795 192405 123796
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 188843 107812 188909 107813
rect 188843 107748 188844 107812
rect 188908 107748 188909 107812
rect 188843 107747 188909 107748
rect 189234 82894 189854 118338
rect 189947 96932 190013 96933
rect 189947 96868 189948 96932
rect 190012 96868 190013 96932
rect 189947 96867 190013 96868
rect 189950 86733 190010 96867
rect 192342 92581 192402 123795
rect 192339 92580 192405 92581
rect 192339 92516 192340 92580
rect 192404 92516 192405 92580
rect 192339 92515 192405 92516
rect 189947 86732 190013 86733
rect 189947 86668 189948 86732
rect 190012 86668 190013 86732
rect 189947 86667 190013 86668
rect 192710 86189 192770 131411
rect 193811 102236 193877 102237
rect 193811 102172 193812 102236
rect 193876 102172 193877 102236
rect 193811 102171 193877 102172
rect 192954 86614 193574 90782
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192707 86188 192773 86189
rect 192707 86124 192708 86188
rect 192772 86124 192773 86188
rect 192707 86123 192773 86124
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 186819 6220 186885 6221
rect 186819 6156 186820 6220
rect 186884 6156 186885 6220
rect 186819 6155 186885 6156
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 193814 85509 193874 102171
rect 193811 85508 193877 85509
rect 193811 85444 193812 85508
rect 193876 85444 193877 85508
rect 193811 85443 193877 85444
rect 194547 85508 194613 85509
rect 194547 85444 194548 85508
rect 194612 85444 194613 85508
rect 194547 85443 194613 85444
rect 194550 84829 194610 85443
rect 194547 84828 194613 84829
rect 194547 84764 194548 84828
rect 194612 84764 194613 84828
rect 194547 84763 194613 84764
rect 195102 82109 195162 140387
rect 195099 82108 195165 82109
rect 195099 82044 195100 82108
rect 195164 82044 195165 82108
rect 195099 82043 195165 82044
rect 196574 79389 196634 142291
rect 199388 111454 199708 111486
rect 199388 111218 199430 111454
rect 199666 111218 199708 111454
rect 199388 111134 199708 111218
rect 199388 110898 199430 111134
rect 199666 110898 199708 111134
rect 199388 110866 199708 110898
rect 200622 93397 200682 179963
rect 200619 93396 200685 93397
rect 200619 93332 200620 93396
rect 200684 93332 200685 93396
rect 200619 93331 200685 93332
rect 201542 92445 201602 239395
rect 203514 205174 204134 239592
rect 205587 215932 205653 215933
rect 205587 215868 205588 215932
rect 205652 215868 205653 215932
rect 205587 215867 205653 215868
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 143035 204134 168618
rect 205590 147690 205650 215867
rect 205406 147630 205650 147690
rect 207234 208894 207854 239592
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 203195 142220 203261 142221
rect 203195 142156 203196 142220
rect 203260 142156 203261 142220
rect 203195 142155 203261 142156
rect 201539 92444 201605 92445
rect 201539 92380 201540 92444
rect 201604 92380 201605 92444
rect 201539 92379 201605 92380
rect 196571 79388 196637 79389
rect 196571 79324 196572 79388
rect 196636 79324 196637 79388
rect 196571 79323 196637 79324
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 90782
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 203198 40629 203258 142155
rect 205406 138030 205466 147630
rect 207234 143035 207854 172338
rect 210954 212614 211574 239592
rect 211659 237964 211725 237965
rect 211659 237900 211660 237964
rect 211724 237900 211725 237964
rect 211659 237899 211725 237900
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 143035 211574 176058
rect 209819 140588 209885 140589
rect 209819 140524 209820 140588
rect 209884 140524 209885 140588
rect 209819 140523 209885 140524
rect 205406 137970 205650 138030
rect 204264 129454 204584 129486
rect 204264 129218 204306 129454
rect 204542 129218 204584 129454
rect 204264 129134 204584 129218
rect 204264 128898 204306 129134
rect 204542 128898 204584 129134
rect 204264 128866 204584 128898
rect 203514 61174 204134 90782
rect 205590 90269 205650 137970
rect 209140 111454 209460 111486
rect 209140 111218 209182 111454
rect 209418 111218 209460 111454
rect 209140 111134 209460 111218
rect 209140 110898 209182 111134
rect 209418 110898 209460 111134
rect 209140 110866 209460 110898
rect 209822 93397 209882 140523
rect 209819 93396 209885 93397
rect 209819 93332 209820 93396
rect 209884 93332 209885 93396
rect 209819 93331 209885 93332
rect 211662 92445 211722 237899
rect 217794 219454 218414 239592
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 215339 216748 215405 216749
rect 215339 216684 215340 216748
rect 215404 216684 215405 216748
rect 215339 216683 215405 216684
rect 214016 129454 214336 129486
rect 214016 129218 214058 129454
rect 214294 129218 214336 129454
rect 214016 129134 214336 129218
rect 214016 128898 214058 129134
rect 214294 128898 214336 129134
rect 214016 128866 214336 128898
rect 211659 92444 211725 92445
rect 211659 92380 211660 92444
rect 211724 92380 211725 92444
rect 211659 92379 211725 92380
rect 205587 90268 205653 90269
rect 205587 90204 205588 90268
rect 205652 90204 205653 90268
rect 205587 90203 205653 90204
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203195 40628 203261 40629
rect 203195 40564 203196 40628
rect 203260 40564 203261 40628
rect 203195 40563 203261 40564
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 90782
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 90782
rect 215342 90269 215402 216683
rect 217794 183454 218414 218898
rect 221514 223174 222134 239592
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 219571 208316 219637 208317
rect 219571 208252 219572 208316
rect 219636 208252 219637 208316
rect 219571 208251 219637 208252
rect 219574 207770 219634 208251
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 143035 218414 146898
rect 219206 207710 219634 207770
rect 219206 139090 219266 207710
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 143035 222134 150618
rect 225234 226894 225854 239592
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 224907 148476 224973 148477
rect 224907 148412 224908 148476
rect 224972 148412 224973 148476
rect 224907 148411 224973 148412
rect 223619 144804 223685 144805
rect 223619 144740 223620 144804
rect 223684 144740 223685 144804
rect 223619 144739 223685 144740
rect 219206 139030 219634 139090
rect 218892 111454 219212 111486
rect 218892 111218 218934 111454
rect 219170 111218 219212 111454
rect 218892 111134 219212 111218
rect 218892 110898 218934 111134
rect 219170 110898 219212 111134
rect 218892 110866 219212 110898
rect 219574 93870 219634 139030
rect 223622 132510 223682 144739
rect 224355 142492 224421 142493
rect 224355 142428 224356 142492
rect 224420 142428 224421 142492
rect 224355 142427 224421 142428
rect 224358 133517 224418 142427
rect 224355 133516 224421 133517
rect 224355 133452 224356 133516
rect 224420 133452 224421 133516
rect 224355 133451 224421 133452
rect 223622 132450 224418 132510
rect 224358 129029 224418 132450
rect 224355 129028 224421 129029
rect 224355 128964 224356 129028
rect 224420 128964 224421 129028
rect 224355 128963 224421 128964
rect 224910 121413 224970 148411
rect 225234 143035 225854 154338
rect 228954 230614 229574 239592
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 226379 140724 226445 140725
rect 226379 140660 226380 140724
rect 226444 140660 226445 140724
rect 226379 140659 226445 140660
rect 224907 121412 224973 121413
rect 224907 121348 224908 121412
rect 224972 121348 224973 121412
rect 224907 121347 224973 121348
rect 226382 119509 226442 140659
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 226379 119508 226445 119509
rect 226379 119444 226380 119508
rect 226444 119444 226445 119508
rect 226379 119443 226445 119444
rect 227667 108356 227733 108357
rect 227667 108292 227668 108356
rect 227732 108292 227733 108356
rect 227667 108291 227733 108292
rect 224355 99516 224421 99517
rect 224355 99452 224356 99516
rect 224420 99452 224421 99516
rect 224355 99451 224421 99452
rect 219206 93810 219634 93870
rect 219206 91085 219266 93810
rect 224358 92309 224418 99451
rect 226379 97204 226445 97205
rect 226379 97140 226380 97204
rect 226444 97140 226445 97204
rect 226379 97139 226445 97140
rect 224355 92308 224421 92309
rect 224355 92244 224356 92308
rect 224420 92244 224421 92308
rect 224355 92243 224421 92244
rect 219203 91084 219269 91085
rect 219203 91020 219204 91084
rect 219268 91020 219269 91084
rect 219203 91019 219269 91020
rect 215339 90268 215405 90269
rect 215339 90204 215340 90268
rect 215404 90204 215405 90268
rect 215339 90203 215405 90204
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 90782
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 90782
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 90782
rect 226382 86733 226442 97139
rect 227670 87957 227730 108291
rect 227667 87956 227733 87957
rect 227667 87892 227668 87956
rect 227732 87892 227733 87956
rect 227667 87891 227733 87892
rect 226379 86732 226445 86733
rect 226379 86668 226380 86732
rect 226444 86668 226445 86732
rect 226379 86667 226445 86668
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 237454 236414 239592
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 205174 240134 239592
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 242942 200701 243002 241979
rect 243234 208894 243854 239592
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 242939 200700 243005 200701
rect 242939 200636 242940 200700
rect 243004 200636 243005 200700
rect 242939 200635 243005 200636
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 212614 247574 239592
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 251774 92173 251834 300867
rect 255270 297397 255330 329019
rect 256739 311268 256805 311269
rect 256739 311204 256740 311268
rect 256804 311204 256805 311268
rect 256739 311203 256805 311204
rect 256742 298757 256802 311203
rect 256739 298756 256805 298757
rect 256739 298692 256740 298756
rect 256804 298692 256805 298756
rect 256739 298691 256805 298692
rect 255267 297396 255333 297397
rect 255267 297332 255268 297396
rect 255332 297332 255333 297396
rect 255267 297331 255333 297332
rect 257514 295174 258134 330618
rect 258398 316050 258458 333235
rect 259683 331804 259749 331805
rect 259683 331740 259684 331804
rect 259748 331740 259749 331804
rect 259683 331739 259749 331740
rect 259499 327180 259565 327181
rect 259499 327116 259500 327180
rect 259564 327116 259565 327180
rect 259499 327115 259565 327116
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 258214 315990 258458 316050
rect 258214 287070 258274 315990
rect 258763 300796 258829 300797
rect 258763 300732 258764 300796
rect 258828 300732 258829 300796
rect 258763 300731 258829 300732
rect 258766 298077 258826 300731
rect 258763 298076 258829 298077
rect 258763 298012 258764 298076
rect 258828 298012 258829 298076
rect 258763 298011 258829 298012
rect 258395 293996 258461 293997
rect 258395 293932 258396 293996
rect 258460 293932 258461 293996
rect 258395 293931 258461 293932
rect 258398 290869 258458 293931
rect 258395 290868 258461 290869
rect 258395 290804 258396 290868
rect 258460 290804 258461 290868
rect 258395 290803 258461 290804
rect 259502 288829 259562 327115
rect 259686 293589 259746 331739
rect 260971 307052 261037 307053
rect 260971 306988 260972 307052
rect 261036 306988 261037 307052
rect 260971 306987 261037 306988
rect 259683 293588 259749 293589
rect 259683 293524 259684 293588
rect 259748 293524 259749 293588
rect 259683 293523 259749 293524
rect 259683 289780 259749 289781
rect 259683 289716 259684 289780
rect 259748 289716 259749 289780
rect 259683 289715 259749 289716
rect 259499 288828 259565 288829
rect 259499 288764 259500 288828
rect 259564 288764 259565 288828
rect 259499 288763 259565 288764
rect 258214 287010 258458 287070
rect 258398 270877 258458 287010
rect 259686 277410 259746 289715
rect 260974 278221 261034 306987
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 260971 278220 261037 278221
rect 260971 278156 260972 278220
rect 261036 278156 261037 278220
rect 260971 278155 261037 278156
rect 259502 277350 259746 277410
rect 259315 272508 259381 272509
rect 259315 272444 259316 272508
rect 259380 272444 259381 272508
rect 259315 272443 259381 272444
rect 258395 270876 258461 270877
rect 258395 270812 258396 270876
rect 258460 270812 258461 270876
rect 258395 270811 258461 270812
rect 259131 270876 259197 270877
rect 259131 270812 259132 270876
rect 259196 270812 259197 270876
rect 259131 270811 259197 270812
rect 259134 265573 259194 270811
rect 259131 265572 259197 265573
rect 259131 265508 259132 265572
rect 259196 265508 259197 265572
rect 259131 265507 259197 265508
rect 259131 263668 259197 263669
rect 259131 263604 259132 263668
rect 259196 263604 259197 263668
rect 259131 263603 259197 263604
rect 258579 261084 258645 261085
rect 258579 261020 258580 261084
rect 258644 261020 258645 261084
rect 258579 261019 258645 261020
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257291 246396 257357 246397
rect 257291 246332 257292 246396
rect 257356 246332 257357 246396
rect 257291 246331 257357 246332
rect 252875 243268 252941 243269
rect 252875 243204 252876 243268
rect 252940 243204 252941 243268
rect 252875 243203 252941 243204
rect 252878 241093 252938 243203
rect 252875 241092 252941 241093
rect 252875 241028 252876 241092
rect 252940 241028 252941 241092
rect 252875 241027 252941 241028
rect 253794 219454 254414 239592
rect 257294 236061 257354 246331
rect 257291 236060 257357 236061
rect 257291 235996 257292 236060
rect 257356 235996 257357 236060
rect 257291 235995 257357 235996
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 251771 92172 251837 92173
rect 251771 92108 251772 92172
rect 251836 92108 251837 92172
rect 251771 92107 251837 92108
rect 251774 91765 251834 92107
rect 251771 91764 251837 91765
rect 251771 91700 251772 91764
rect 251836 91700 251837 91764
rect 251771 91699 251837 91700
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 223174 258134 258618
rect 258582 257141 258642 261019
rect 259134 260949 259194 263603
rect 259131 260948 259197 260949
rect 259131 260884 259132 260948
rect 259196 260884 259197 260948
rect 259131 260883 259197 260884
rect 258579 257140 258645 257141
rect 258579 257076 258580 257140
rect 258644 257076 258645 257140
rect 258579 257075 258645 257076
rect 258395 252788 258461 252789
rect 258395 252724 258396 252788
rect 258460 252724 258461 252788
rect 258395 252723 258461 252724
rect 258398 252650 258458 252723
rect 258214 252590 258458 252650
rect 258214 238770 258274 252590
rect 259318 250069 259378 272443
rect 258395 250068 258461 250069
rect 258395 250004 258396 250068
rect 258460 250004 258461 250068
rect 258395 250003 258461 250004
rect 259315 250068 259381 250069
rect 259315 250004 259316 250068
rect 259380 250004 259381 250068
rect 259315 250003 259381 250004
rect 258398 240957 258458 250003
rect 258395 240956 258461 240957
rect 258395 240892 258396 240956
rect 258460 240892 258461 240956
rect 258395 240891 258461 240892
rect 258214 238710 258458 238770
rect 258398 234565 258458 238710
rect 258395 234564 258461 234565
rect 258395 234500 258396 234564
rect 258460 234500 258461 234564
rect 258395 234499 258461 234500
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 259502 136645 259562 277350
rect 261234 262894 261854 298338
rect 262262 272781 262322 349827
rect 262446 348533 262506 478075
rect 262443 348532 262509 348533
rect 262443 348468 262444 348532
rect 262508 348468 262509 348532
rect 262443 348467 262509 348468
rect 263550 338741 263610 600475
rect 264954 590614 265574 626058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 270539 596324 270605 596325
rect 270539 596260 270540 596324
rect 270604 596260 270605 596324
rect 270539 596259 270605 596260
rect 269067 592652 269133 592653
rect 269067 592588 269068 592652
rect 269132 592588 269133 592652
rect 269067 592587 269133 592588
rect 267779 590748 267845 590749
rect 267779 590684 267780 590748
rect 267844 590684 267845 590748
rect 267779 590683 267845 590684
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 263731 563140 263797 563141
rect 263731 563076 263732 563140
rect 263796 563076 263797 563140
rect 263731 563075 263797 563076
rect 263734 362269 263794 563075
rect 264954 554614 265574 590058
rect 265755 587212 265821 587213
rect 265755 587148 265756 587212
rect 265820 587148 265821 587212
rect 265755 587147 265821 587148
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 265758 381581 265818 587147
rect 266307 586532 266373 586533
rect 266307 586468 266308 586532
rect 266372 586468 266373 586532
rect 266307 586467 266373 586468
rect 265939 382396 266005 382397
rect 265939 382332 265940 382396
rect 266004 382332 266005 382396
rect 265939 382331 266005 382332
rect 265755 381580 265821 381581
rect 265755 381516 265756 381580
rect 265820 381516 265821 381580
rect 265755 381515 265821 381516
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 263731 362268 263797 362269
rect 263731 362204 263732 362268
rect 263796 362204 263797 362268
rect 263731 362203 263797 362204
rect 263547 338740 263613 338741
rect 263547 338676 263548 338740
rect 263612 338676 263613 338740
rect 263547 338675 263613 338676
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 263547 334660 263613 334661
rect 263547 334596 263548 334660
rect 263612 334596 263613 334660
rect 263547 334595 263613 334596
rect 262443 305692 262509 305693
rect 262443 305628 262444 305692
rect 262508 305628 262509 305692
rect 262443 305627 262509 305628
rect 262446 277405 262506 305627
rect 263550 302250 263610 334595
rect 263731 303788 263797 303789
rect 263731 303724 263732 303788
rect 263796 303724 263797 303788
rect 263731 303723 263797 303724
rect 263366 302190 263610 302250
rect 263366 292590 263426 302190
rect 263366 292530 263610 292590
rect 262443 277404 262509 277405
rect 262443 277340 262444 277404
rect 262508 277340 262509 277404
rect 262443 277339 262509 277340
rect 262259 272780 262325 272781
rect 262259 272716 262260 272780
rect 262324 272716 262325 272780
rect 262259 272715 262325 272716
rect 262262 272370 262322 272715
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 262078 272310 262322 272370
rect 262078 205733 262138 272310
rect 263363 267068 263429 267069
rect 263363 267004 263364 267068
rect 263428 267004 263429 267068
rect 263363 267003 263429 267004
rect 263366 253333 263426 267003
rect 263550 259181 263610 292530
rect 263547 259180 263613 259181
rect 263547 259116 263548 259180
rect 263612 259116 263613 259180
rect 263547 259115 263613 259116
rect 263547 254012 263613 254013
rect 263547 253948 263548 254012
rect 263612 253948 263613 254012
rect 263547 253947 263613 253948
rect 262259 253332 262325 253333
rect 262259 253268 262260 253332
rect 262324 253268 262325 253332
rect 262259 253267 262325 253268
rect 263363 253332 263429 253333
rect 263363 253268 263364 253332
rect 263428 253268 263429 253332
rect 263363 253267 263429 253268
rect 262075 205732 262141 205733
rect 262075 205668 262076 205732
rect 262140 205668 262141 205732
rect 262075 205667 262141 205668
rect 262262 193901 262322 253267
rect 262443 253196 262509 253197
rect 262443 253132 262444 253196
rect 262508 253132 262509 253196
rect 262443 253131 262509 253132
rect 262446 236605 262506 253131
rect 262443 236604 262509 236605
rect 262443 236540 262444 236604
rect 262508 236540 262509 236604
rect 262443 236539 262509 236540
rect 262259 193900 262325 193901
rect 262259 193836 262260 193900
rect 262324 193836 262325 193900
rect 262259 193835 262325 193836
rect 263550 192541 263610 253947
rect 263734 239461 263794 303723
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 263731 239460 263797 239461
rect 263731 239396 263732 239460
rect 263796 239396 263797 239460
rect 263731 239395 263797 239396
rect 264954 230614 265574 266058
rect 265942 263533 266002 382331
rect 266310 351117 266370 586467
rect 266859 361724 266925 361725
rect 266859 361660 266860 361724
rect 266924 361660 266925 361724
rect 266859 361659 266925 361660
rect 266307 351116 266373 351117
rect 266307 351052 266308 351116
rect 266372 351052 266373 351116
rect 266307 351051 266373 351052
rect 266307 330444 266373 330445
rect 266307 330380 266308 330444
rect 266372 330380 266373 330444
rect 266307 330379 266373 330380
rect 265939 263532 266005 263533
rect 265939 263468 265940 263532
rect 266004 263468 266005 263532
rect 265939 263467 266005 263468
rect 265942 263125 266002 263467
rect 265939 263124 266005 263125
rect 265939 263060 265940 263124
rect 266004 263060 266005 263124
rect 265939 263059 266005 263060
rect 266310 262989 266370 330379
rect 266862 277410 266922 361659
rect 267782 320109 267842 590683
rect 267963 376684 268029 376685
rect 267963 376620 267964 376684
rect 268028 376620 268029 376684
rect 267963 376619 268029 376620
rect 267779 320108 267845 320109
rect 267779 320044 267780 320108
rect 267844 320044 267845 320108
rect 267779 320043 267845 320044
rect 267779 319428 267845 319429
rect 267779 319364 267780 319428
rect 267844 319364 267845 319428
rect 267779 319363 267845 319364
rect 267782 278901 267842 319363
rect 267779 278900 267845 278901
rect 267779 278836 267780 278900
rect 267844 278836 267845 278900
rect 267779 278835 267845 278836
rect 266494 277350 266922 277410
rect 266494 270197 266554 277350
rect 266491 270196 266557 270197
rect 266491 270132 266492 270196
rect 266556 270132 266557 270196
rect 266491 270131 266557 270132
rect 266494 269245 266554 270131
rect 266491 269244 266557 269245
rect 266491 269180 266492 269244
rect 266556 269180 266557 269244
rect 266491 269179 266557 269180
rect 266307 262988 266373 262989
rect 266307 262924 266308 262988
rect 266372 262924 266373 262988
rect 266307 262923 266373 262924
rect 266491 259724 266557 259725
rect 266491 259660 266492 259724
rect 266556 259660 266557 259724
rect 266491 259659 266557 259660
rect 266307 255916 266373 255917
rect 266307 255852 266308 255916
rect 266372 255852 266373 255916
rect 266307 255851 266373 255852
rect 266310 251973 266370 255851
rect 266307 251972 266373 251973
rect 266307 251908 266308 251972
rect 266372 251908 266373 251972
rect 266307 251907 266373 251908
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263547 192540 263613 192541
rect 263547 192476 263548 192540
rect 263612 192476 263613 192540
rect 263547 192475 263613 192476
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 259499 136644 259565 136645
rect 259499 136580 259500 136644
rect 259564 136580 259565 136644
rect 259499 136579 259565 136580
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 158614 265574 194058
rect 266310 166973 266370 251907
rect 266494 231301 266554 259659
rect 267966 257141 268026 376619
rect 269070 356693 269130 592587
rect 270542 376005 270602 596259
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 276243 600404 276309 600405
rect 276243 600340 276244 600404
rect 276308 600340 276309 600404
rect 276243 600339 276309 600340
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 273299 452436 273365 452437
rect 273299 452372 273300 452436
rect 273364 452372 273365 452436
rect 273299 452371 273365 452372
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 270539 376004 270605 376005
rect 270539 375940 270540 376004
rect 270604 375940 270605 376004
rect 270539 375939 270605 375940
rect 271091 360228 271157 360229
rect 271091 360164 271092 360228
rect 271156 360164 271157 360228
rect 271091 360163 271157 360164
rect 269067 356692 269133 356693
rect 269067 356628 269068 356692
rect 269132 356628 269133 356692
rect 269067 356627 269133 356628
rect 270539 329220 270605 329221
rect 270539 329156 270540 329220
rect 270604 329156 270605 329220
rect 270539 329155 270605 329156
rect 269619 307732 269685 307733
rect 269619 307668 269620 307732
rect 269684 307668 269685 307732
rect 269619 307667 269685 307668
rect 269622 301477 269682 307667
rect 269619 301476 269685 301477
rect 269619 301412 269620 301476
rect 269684 301412 269685 301476
rect 269619 301411 269685 301412
rect 269622 268429 269682 301411
rect 269803 296852 269869 296853
rect 269803 296788 269804 296852
rect 269868 296788 269869 296852
rect 269803 296787 269869 296788
rect 269806 283525 269866 296787
rect 269803 283524 269869 283525
rect 269803 283460 269804 283524
rect 269868 283460 269869 283524
rect 269803 283459 269869 283460
rect 269619 268428 269685 268429
rect 269619 268364 269620 268428
rect 269684 268364 269685 268428
rect 269619 268363 269685 268364
rect 269067 261220 269133 261221
rect 269067 261156 269068 261220
rect 269132 261156 269133 261220
rect 269067 261155 269133 261156
rect 267963 257140 268029 257141
rect 267963 257076 267964 257140
rect 268028 257076 268029 257140
rect 267963 257075 268029 257076
rect 267963 257004 268029 257005
rect 267963 256940 267964 257004
rect 268028 256940 268029 257004
rect 267963 256939 268029 256940
rect 267779 240548 267845 240549
rect 267779 240484 267780 240548
rect 267844 240484 267845 240548
rect 267779 240483 267845 240484
rect 266491 231300 266557 231301
rect 266491 231236 266492 231300
rect 266556 231236 266557 231300
rect 266491 231235 266557 231236
rect 267782 210357 267842 240483
rect 267966 227629 268026 256939
rect 269070 230349 269130 261155
rect 270542 243677 270602 329155
rect 271094 269109 271154 360163
rect 271794 345454 272414 380898
rect 273302 359413 273362 452371
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 273483 360908 273549 360909
rect 273483 360844 273484 360908
rect 273548 360844 273549 360908
rect 273483 360843 273549 360844
rect 273299 359412 273365 359413
rect 273299 359348 273300 359412
rect 273364 359348 273365 359412
rect 273299 359347 273365 359348
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 273299 305828 273365 305829
rect 273299 305764 273300 305828
rect 273364 305764 273365 305828
rect 273299 305763 273365 305764
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271091 269108 271157 269109
rect 271091 269044 271092 269108
rect 271156 269044 271157 269108
rect 271091 269043 271157 269044
rect 270723 257956 270789 257957
rect 270723 257892 270724 257956
rect 270788 257892 270789 257956
rect 270723 257891 270789 257892
rect 270539 243676 270605 243677
rect 270539 243612 270540 243676
rect 270604 243612 270605 243676
rect 270539 243611 270605 243612
rect 269067 230348 269133 230349
rect 269067 230284 269068 230348
rect 269132 230284 269133 230348
rect 269067 230283 269133 230284
rect 267963 227628 268029 227629
rect 267963 227564 267964 227628
rect 268028 227564 268029 227628
rect 267963 227563 268029 227564
rect 270726 223549 270786 257891
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 270723 223548 270789 223549
rect 270723 223484 270724 223548
rect 270788 223484 270789 223548
rect 270723 223483 270789 223484
rect 270726 219450 270786 223483
rect 270542 219390 270786 219450
rect 267779 210356 267845 210357
rect 267779 210292 267780 210356
rect 267844 210292 267845 210356
rect 267779 210291 267845 210292
rect 266307 166972 266373 166973
rect 266307 166908 266308 166972
rect 266372 166908 266373 166972
rect 266307 166907 266373 166908
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 270542 108357 270602 219390
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 270539 108356 270605 108357
rect 270539 108292 270540 108356
rect 270604 108292 270605 108356
rect 270539 108291 270605 108292
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 93454 272414 128898
rect 273302 95845 273362 305763
rect 273486 240005 273546 360843
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 274587 325004 274653 325005
rect 274587 324940 274588 325004
rect 274652 324940 274653 325004
rect 274587 324939 274653 324940
rect 274590 247077 274650 324939
rect 275514 313174 276134 348618
rect 276246 327725 276306 600339
rect 279234 568894 279854 604338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 281579 589932 281645 589933
rect 281579 589868 281580 589932
rect 281644 589868 281645 589932
rect 281579 589867 281645 589868
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 277347 441692 277413 441693
rect 277347 441630 277348 441692
rect 277166 441628 277348 441630
rect 277412 441628 277413 441692
rect 277166 441627 277413 441628
rect 277166 441570 277410 441627
rect 276427 395316 276493 395317
rect 276427 395252 276428 395316
rect 276492 395252 276493 395316
rect 276427 395251 276493 395252
rect 276430 379405 276490 395251
rect 276427 379404 276493 379405
rect 276427 379340 276428 379404
rect 276492 379340 276493 379404
rect 276427 379339 276493 379340
rect 276243 327724 276309 327725
rect 276243 327660 276244 327724
rect 276308 327660 276309 327724
rect 276243 327659 276309 327660
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 274587 247076 274653 247077
rect 274587 247012 274588 247076
rect 274652 247012 274653 247076
rect 274587 247011 274653 247012
rect 275514 241174 276134 276618
rect 276430 258093 276490 379339
rect 277166 304197 277226 441570
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 280291 416804 280357 416805
rect 280291 416740 280292 416804
rect 280356 416740 280357 416804
rect 280291 416739 280357 416740
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 280294 369749 280354 416739
rect 280291 369748 280357 369749
rect 280291 369684 280292 369748
rect 280356 369684 280357 369748
rect 280291 369683 280357 369684
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 277531 349756 277597 349757
rect 277531 349692 277532 349756
rect 277596 349692 277597 349756
rect 277531 349691 277597 349692
rect 277163 304196 277229 304197
rect 277163 304132 277164 304196
rect 277228 304132 277229 304196
rect 277163 304131 277229 304132
rect 276427 258092 276493 258093
rect 276427 258028 276428 258092
rect 276492 258028 276493 258092
rect 276427 258027 276493 258028
rect 277534 243677 277594 349691
rect 279234 316894 279854 352338
rect 280291 325820 280357 325821
rect 280291 325756 280292 325820
rect 280356 325756 280357 325820
rect 280291 325755 280357 325756
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 277899 261356 277965 261357
rect 277899 261292 277900 261356
rect 277964 261292 277965 261356
rect 277899 261291 277965 261292
rect 277531 243676 277597 243677
rect 277531 243612 277532 243676
rect 277596 243612 277597 243676
rect 277531 243611 277597 243612
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 273483 240004 273549 240005
rect 273483 239940 273484 240004
rect 273548 239940 273549 240004
rect 273483 239939 273549 239940
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 277902 181389 277962 261291
rect 279234 244894 279854 280338
rect 280294 255917 280354 325755
rect 281582 308413 281642 589867
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 285627 481676 285693 481677
rect 285627 481612 285628 481676
rect 285692 481612 285693 481676
rect 285627 481611 285693 481612
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 284339 454068 284405 454069
rect 284339 454004 284340 454068
rect 284404 454004 284405 454068
rect 284339 454003 284405 454004
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 281579 308412 281645 308413
rect 281579 308348 281580 308412
rect 281644 308348 281645 308412
rect 281579 308347 281645 308348
rect 281582 262173 281642 308347
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 281579 262172 281645 262173
rect 281579 262108 281580 262172
rect 281644 262108 281645 262172
rect 281579 262107 281645 262108
rect 280291 255916 280357 255917
rect 280291 255852 280292 255916
rect 280356 255852 280357 255916
rect 280291 255851 280357 255852
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 277899 181388 277965 181389
rect 277899 181324 277900 181388
rect 277964 181324 277965 181388
rect 277899 181323 277965 181324
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 273299 95844 273365 95845
rect 273299 95780 273300 95844
rect 273364 95780 273365 95844
rect 273299 95779 273365 95780
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 248614 283574 284058
rect 284342 260133 284402 454003
rect 284339 260132 284405 260133
rect 284339 260068 284340 260132
rect 284404 260068 284405 260132
rect 284339 260067 284405 260068
rect 285630 256733 285690 481611
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 287099 418300 287165 418301
rect 287099 418236 287100 418300
rect 287164 418236 287165 418300
rect 287099 418235 287165 418236
rect 287102 378045 287162 418235
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 287099 378044 287165 378045
rect 287099 377980 287100 378044
rect 287164 377980 287165 378044
rect 287099 377979 287165 377980
rect 287102 267205 287162 377979
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 287099 267204 287165 267205
rect 287099 267140 287100 267204
rect 287164 267140 287165 267204
rect 287099 267139 287165 267140
rect 285627 256732 285693 256733
rect 285627 256668 285628 256732
rect 285692 256668 285693 256732
rect 285627 256667 285693 256668
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 73721 543218 73957 543454
rect 73721 542898 73957 543134
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77686 561218 77922 561454
rect 77686 560898 77922 561134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81651 543218 81887 543454
rect 81651 542898 81887 543134
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 85617 561218 85853 561454
rect 85617 560898 85853 561134
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 89582 543218 89818 543454
rect 89582 542898 89818 543134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 79019 273218 79255 273454
rect 79019 272898 79255 273134
rect 74387 255218 74623 255454
rect 74387 254898 74623 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 83651 255218 83887 255454
rect 83651 254898 83887 255134
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 88283 273218 88519 273454
rect 88283 272898 88519 273134
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 92915 255218 93151 255454
rect 92915 254898 93151 255134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 77686 129218 77922 129454
rect 77686 128898 77922 129134
rect 85617 129218 85853 129454
rect 85617 128898 85853 129134
rect 73721 111218 73957 111454
rect 73721 110898 73957 111134
rect 81651 111218 81887 111454
rect 81651 110898 81887 111134
rect 89582 111218 89818 111454
rect 89582 110898 89818 111134
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 197818 579218 198054 579454
rect 197818 578898 198054 579134
rect 197818 543218 198054 543454
rect 197818 542898 198054 543134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 213178 561218 213414 561454
rect 213178 560898 213414 561134
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228538 579218 228774 579454
rect 228538 578898 228774 579134
rect 228538 543218 228774 543454
rect 228538 542898 228774 543134
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 197818 435218 198054 435454
rect 197818 434898 198054 435134
rect 228538 435218 228774 435454
rect 228538 434898 228774 435134
rect 213178 417218 213414 417454
rect 213178 416898 213414 417134
rect 197818 399218 198054 399454
rect 197818 398898 198054 399134
rect 228538 399218 228774 399454
rect 228538 398898 228774 399134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243898 561218 244134 561454
rect 243898 560898 244134 561134
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243898 417218 244134 417454
rect 243898 416898 244134 417134
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 197818 291218 198054 291454
rect 197818 290898 198054 291134
rect 228538 291218 228774 291454
rect 228538 290898 228774 291134
rect 213178 273218 213414 273454
rect 213178 272898 213414 273134
rect 243898 273218 244134 273454
rect 243898 272898 244134 273134
rect 197818 255218 198054 255454
rect 197818 254898 198054 255134
rect 228538 255218 228774 255454
rect 228538 254898 228774 255134
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 199430 111218 199666 111454
rect 199430 110898 199666 111134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 204306 129218 204542 129454
rect 204306 128898 204542 129134
rect 209182 111218 209418 111454
rect 209182 110898 209418 111134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 214058 129218 214294 129454
rect 214058 128898 214294 129134
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 218934 111218 219170 111454
rect 218934 110898 219170 111134
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 197818 579454
rect 198054 579218 228538 579454
rect 228774 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 197818 579134
rect 198054 578898 228538 579134
rect 228774 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 77686 561454
rect 77922 561218 85617 561454
rect 85853 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 213178 561454
rect 213414 561218 243898 561454
rect 244134 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 77686 561134
rect 77922 560898 85617 561134
rect 85853 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 213178 561134
rect 213414 560898 243898 561134
rect 244134 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73721 543454
rect 73957 543218 81651 543454
rect 81887 543218 89582 543454
rect 89818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 197818 543454
rect 198054 543218 228538 543454
rect 228774 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73721 543134
rect 73957 542898 81651 543134
rect 81887 542898 89582 543134
rect 89818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 197818 543134
rect 198054 542898 228538 543134
rect 228774 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 197818 435454
rect 198054 435218 228538 435454
rect 228774 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 197818 435134
rect 198054 434898 228538 435134
rect 228774 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 213178 417454
rect 213414 417218 243898 417454
rect 244134 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 213178 417134
rect 213414 416898 243898 417134
rect 244134 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 197818 399454
rect 198054 399218 228538 399454
rect 228774 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 197818 399134
rect 198054 398898 228538 399134
rect 228774 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 197818 291454
rect 198054 291218 228538 291454
rect 228774 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 197818 291134
rect 198054 290898 228538 291134
rect 228774 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 79019 273454
rect 79255 273218 88283 273454
rect 88519 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 213178 273454
rect 213414 273218 243898 273454
rect 244134 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 79019 273134
rect 79255 272898 88283 273134
rect 88519 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 213178 273134
rect 213414 272898 243898 273134
rect 244134 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74387 255454
rect 74623 255218 83651 255454
rect 83887 255218 92915 255454
rect 93151 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 197818 255454
rect 198054 255218 228538 255454
rect 228774 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74387 255134
rect 74623 254898 83651 255134
rect 83887 254898 92915 255134
rect 93151 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 197818 255134
rect 198054 254898 228538 255134
rect 228774 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 77686 129454
rect 77922 129218 85617 129454
rect 85853 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 204306 129454
rect 204542 129218 214058 129454
rect 214294 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 77686 129134
rect 77922 128898 85617 129134
rect 85853 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 204306 129134
rect 204542 128898 214058 129134
rect 214294 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73721 111454
rect 73957 111218 81651 111454
rect 81887 111218 89582 111454
rect 89818 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 199430 111454
rect 199666 111218 209182 111454
rect 209418 111218 218934 111454
rect 219170 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73721 111134
rect 73957 110898 81651 111134
rect 81887 110898 89582 111134
rect 89818 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 199430 111134
rect 199666 110898 209182 111134
rect 209418 110898 218934 111134
rect 219170 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use zube_wrapped_project  zube_wrapped_project_5
timestamp 1636115455
transform 1 0 193568 0 1 241592
box 0 0 60000 60000
use wrapped_ws2812  wrapped_ws2812_4
timestamp 1636115455
transform 1 0 193568 0 1 92782
box 0 0 31475 48253
use wrapped_vga_clock  wrapped_vga_clock_2
timestamp 1636115455
transform 1 0 68770 0 1 390356
box 0 0 44000 44000
use wrapped_tpm2137  wrapped_tpm2137_3
timestamp 1636115455
transform 1 0 68770 0 1 539166
box 0 0 26000 42000
use wrapped_rgb_mixer  wrapped_rgb_mixer_0
timestamp 1636115455
transform 1 0 68770 0 1 92782
box 0 0 26000 42000
use wrapped_nco  wrapped_nco_7
timestamp 1636115455
transform 1 0 193568 0 1 539166
box 0 0 60000 60000
use wrapped_hack_soc  wrapped_hack_soc_6
timestamp 1636115455
transform 1 0 193568 0 1 390356
box 0 0 60000 60000
use wrapped_frequency_counter  wrapped_frequency_counter_1
timestamp 1636115455
transform 1 0 68770 0 1 241592
box 0 0 30000 42000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 136782 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 143035 218414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 303592 218414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 303592 254414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 436356 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 452356 218414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 452356 254414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 583166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 436356 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 601166 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 601166 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 136782 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 143035 222134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 303592 222134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 436356 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 452356 222134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 583166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 436356 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 601166 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 136782 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 143035 225854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 303592 225854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 436356 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 452356 225854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 583166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 601166 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 136782 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 143035 193574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 303592 193574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 303592 229574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 436356 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 452356 193574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 452356 229574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 583166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 601166 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 601166 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 90782 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 143035 207854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 303592 207854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 303592 243854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 452356 207854 537166 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 452356 243854 537166 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 436356 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 601166 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 601166 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 136782 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 143035 211574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 303592 211574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 303592 247574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 436356 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 452356 211574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 452356 247574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 583166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 436356 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 601166 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 601166 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 136782 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 143035 200414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 303592 200414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 303592 236414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 436356 92414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 452356 200414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 452356 236414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 583166 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 601166 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 601166 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 136782 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 143035 204134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 303592 204134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 303592 240134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 436356 96134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 452356 204134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 452356 240134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 583166 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 601166 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 601166 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
